/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */


assign int_rd_req_desc_0_size_txn_size = int_rd_req_desc_n_size_txn_size['h0];
assign int_rd_req_desc_0_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h0];
assign int_rd_req_desc_0_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h0];
assign int_rd_req_desc_0_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h0];
assign int_rd_req_desc_0_attr_axbar = int_rd_req_desc_n_attr_axbar['h0];
assign int_rd_req_desc_0_attr_axregion = int_rd_req_desc_n_attr_axregion['h0];
assign int_rd_req_desc_0_attr_axqos = int_rd_req_desc_n_attr_axqos['h0];
assign int_rd_req_desc_0_attr_axprot = int_rd_req_desc_n_attr_axprot['h0];
assign int_rd_req_desc_0_attr_axcache = int_rd_req_desc_n_attr_axcache['h0];
assign int_rd_req_desc_0_attr_axlock = int_rd_req_desc_n_attr_axlock['h0];
assign int_rd_req_desc_0_attr_axburst = int_rd_req_desc_n_attr_axburst['h0];
assign int_rd_req_desc_0_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h0];
assign int_rd_req_desc_0_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h0];
assign int_rd_req_desc_0_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h0];
assign int_rd_req_desc_0_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h0];
assign int_rd_req_desc_0_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h0];
assign int_rd_req_desc_0_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h0];
assign int_rd_req_desc_0_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h0];
assign int_rd_req_desc_0_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h0];
assign int_rd_req_desc_0_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h0];
assign int_rd_req_desc_0_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h0];
assign int_rd_req_desc_0_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h0];
assign int_rd_req_desc_0_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h0];
assign int_rd_req_desc_0_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h0];
assign int_rd_req_desc_0_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h0];
assign int_rd_req_desc_0_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h0];
assign int_rd_req_desc_0_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h0];
assign int_rd_req_desc_0_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h0];
assign int_rd_req_desc_0_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h0];
assign int_rd_req_desc_0_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h0];
assign int_rd_req_desc_0_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h0];
assign int_rd_req_desc_0_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h0];
assign int_rd_req_desc_0_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h0];
assign int_rd_req_desc_0_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h0];
assign int_rd_req_desc_0_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h0];
assign int_wr_req_desc_0_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h0];
assign int_wr_req_desc_0_size_txn_size = int_wr_req_desc_n_size_txn_size['h0];
assign int_wr_req_desc_0_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h0];
assign int_wr_req_desc_0_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h0];
assign int_wr_req_desc_0_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h0];
assign int_wr_req_desc_0_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h0];
assign int_wr_req_desc_0_attr_axbar = int_wr_req_desc_n_attr_axbar['h0];
assign int_wr_req_desc_0_attr_awunique = int_wr_req_desc_n_attr_awunique['h0];
assign int_wr_req_desc_0_attr_axregion = int_wr_req_desc_n_attr_axregion['h0];
assign int_wr_req_desc_0_attr_axqos = int_wr_req_desc_n_attr_axqos['h0];
assign int_wr_req_desc_0_attr_axprot = int_wr_req_desc_n_attr_axprot['h0];
assign int_wr_req_desc_0_attr_axcache = int_wr_req_desc_n_attr_axcache['h0];
assign int_wr_req_desc_0_attr_axlock = int_wr_req_desc_n_attr_axlock['h0];
assign int_wr_req_desc_0_attr_axburst = int_wr_req_desc_n_attr_axburst['h0];
assign int_wr_req_desc_0_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h0];
assign int_wr_req_desc_0_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h0];
assign int_wr_req_desc_0_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h0];
assign int_wr_req_desc_0_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h0];
assign int_wr_req_desc_0_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h0];
assign int_wr_req_desc_0_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h0];
assign int_wr_req_desc_0_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h0];
assign int_wr_req_desc_0_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h0];
assign int_wr_req_desc_0_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h0];
assign int_wr_req_desc_0_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h0];
assign int_wr_req_desc_0_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h0];
assign int_wr_req_desc_0_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h0];
assign int_wr_req_desc_0_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h0];
assign int_wr_req_desc_0_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h0];
assign int_wr_req_desc_0_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h0];
assign int_wr_req_desc_0_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h0];
assign int_wr_req_desc_0_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h0];
assign int_wr_req_desc_0_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h0];
assign int_wr_req_desc_0_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h0];
assign int_wr_req_desc_0_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h0];
assign int_wr_req_desc_0_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h0];
assign int_wr_req_desc_0_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h0];
assign int_wr_req_desc_0_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h0];
assign int_wr_req_desc_0_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h0];
assign int_wr_req_desc_0_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h0];
assign int_wr_req_desc_0_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h0];
assign int_wr_req_desc_0_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h0];
assign int_wr_req_desc_0_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h0];
assign int_wr_req_desc_0_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h0];
assign int_wr_req_desc_0_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h0];
assign int_wr_req_desc_0_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h0];
assign int_wr_req_desc_0_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h0];
assign int_wr_req_desc_0_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h0];
assign int_wr_req_desc_0_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h0];
assign int_wr_req_desc_0_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h0];
assign int_wr_req_desc_0_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h0];
assign int_wr_req_desc_0_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h0];
assign int_wr_req_desc_0_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h0];
assign int_wr_req_desc_0_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h0];
assign int_wr_req_desc_0_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h0];
assign int_sn_resp_desc_0_resp_resp = int_sn_resp_desc_n_resp_resp['h0];
assign int_rd_req_desc_1_size_txn_size = int_rd_req_desc_n_size_txn_size['h1];
assign int_rd_req_desc_1_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h1];
assign int_rd_req_desc_1_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h1];
assign int_rd_req_desc_1_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h1];
assign int_rd_req_desc_1_attr_axbar = int_rd_req_desc_n_attr_axbar['h1];
assign int_rd_req_desc_1_attr_axregion = int_rd_req_desc_n_attr_axregion['h1];
assign int_rd_req_desc_1_attr_axqos = int_rd_req_desc_n_attr_axqos['h1];
assign int_rd_req_desc_1_attr_axprot = int_rd_req_desc_n_attr_axprot['h1];
assign int_rd_req_desc_1_attr_axcache = int_rd_req_desc_n_attr_axcache['h1];
assign int_rd_req_desc_1_attr_axlock = int_rd_req_desc_n_attr_axlock['h1];
assign int_rd_req_desc_1_attr_axburst = int_rd_req_desc_n_attr_axburst['h1];
assign int_rd_req_desc_1_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h1];
assign int_rd_req_desc_1_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h1];
assign int_rd_req_desc_1_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h1];
assign int_rd_req_desc_1_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h1];
assign int_rd_req_desc_1_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h1];
assign int_rd_req_desc_1_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h1];
assign int_rd_req_desc_1_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h1];
assign int_rd_req_desc_1_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h1];
assign int_rd_req_desc_1_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h1];
assign int_rd_req_desc_1_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h1];
assign int_rd_req_desc_1_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h1];
assign int_rd_req_desc_1_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h1];
assign int_rd_req_desc_1_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h1];
assign int_rd_req_desc_1_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h1];
assign int_rd_req_desc_1_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h1];
assign int_rd_req_desc_1_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h1];
assign int_rd_req_desc_1_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h1];
assign int_rd_req_desc_1_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h1];
assign int_rd_req_desc_1_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h1];
assign int_rd_req_desc_1_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h1];
assign int_rd_req_desc_1_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h1];
assign int_rd_req_desc_1_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h1];
assign int_rd_req_desc_1_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h1];
assign int_rd_req_desc_1_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h1];
assign int_wr_req_desc_1_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h1];
assign int_wr_req_desc_1_size_txn_size = int_wr_req_desc_n_size_txn_size['h1];
assign int_wr_req_desc_1_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h1];
assign int_wr_req_desc_1_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h1];
assign int_wr_req_desc_1_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h1];
assign int_wr_req_desc_1_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h1];
assign int_wr_req_desc_1_attr_axbar = int_wr_req_desc_n_attr_axbar['h1];
assign int_wr_req_desc_1_attr_awunique = int_wr_req_desc_n_attr_awunique['h1];
assign int_wr_req_desc_1_attr_axregion = int_wr_req_desc_n_attr_axregion['h1];
assign int_wr_req_desc_1_attr_axqos = int_wr_req_desc_n_attr_axqos['h1];
assign int_wr_req_desc_1_attr_axprot = int_wr_req_desc_n_attr_axprot['h1];
assign int_wr_req_desc_1_attr_axcache = int_wr_req_desc_n_attr_axcache['h1];
assign int_wr_req_desc_1_attr_axlock = int_wr_req_desc_n_attr_axlock['h1];
assign int_wr_req_desc_1_attr_axburst = int_wr_req_desc_n_attr_axburst['h1];
assign int_wr_req_desc_1_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h1];
assign int_wr_req_desc_1_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h1];
assign int_wr_req_desc_1_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h1];
assign int_wr_req_desc_1_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h1];
assign int_wr_req_desc_1_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h1];
assign int_wr_req_desc_1_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h1];
assign int_wr_req_desc_1_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h1];
assign int_wr_req_desc_1_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h1];
assign int_wr_req_desc_1_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h1];
assign int_wr_req_desc_1_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h1];
assign int_wr_req_desc_1_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h1];
assign int_wr_req_desc_1_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h1];
assign int_wr_req_desc_1_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h1];
assign int_wr_req_desc_1_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h1];
assign int_wr_req_desc_1_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h1];
assign int_wr_req_desc_1_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h1];
assign int_wr_req_desc_1_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h1];
assign int_wr_req_desc_1_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h1];
assign int_wr_req_desc_1_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h1];
assign int_wr_req_desc_1_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h1];
assign int_wr_req_desc_1_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h1];
assign int_wr_req_desc_1_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h1];
assign int_wr_req_desc_1_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h1];
assign int_wr_req_desc_1_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h1];
assign int_wr_req_desc_1_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h1];
assign int_wr_req_desc_1_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h1];
assign int_wr_req_desc_1_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h1];
assign int_wr_req_desc_1_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h1];
assign int_wr_req_desc_1_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h1];
assign int_wr_req_desc_1_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h1];
assign int_wr_req_desc_1_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h1];
assign int_wr_req_desc_1_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h1];
assign int_wr_req_desc_1_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h1];
assign int_wr_req_desc_1_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h1];
assign int_wr_req_desc_1_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h1];
assign int_wr_req_desc_1_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h1];
assign int_wr_req_desc_1_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h1];
assign int_wr_req_desc_1_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h1];
assign int_wr_req_desc_1_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h1];
assign int_wr_req_desc_1_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h1];
assign int_sn_resp_desc_1_resp_resp = int_sn_resp_desc_n_resp_resp['h1];
assign int_rd_req_desc_2_size_txn_size = int_rd_req_desc_n_size_txn_size['h2];
assign int_rd_req_desc_2_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h2];
assign int_rd_req_desc_2_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h2];
assign int_rd_req_desc_2_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h2];
assign int_rd_req_desc_2_attr_axbar = int_rd_req_desc_n_attr_axbar['h2];
assign int_rd_req_desc_2_attr_axregion = int_rd_req_desc_n_attr_axregion['h2];
assign int_rd_req_desc_2_attr_axqos = int_rd_req_desc_n_attr_axqos['h2];
assign int_rd_req_desc_2_attr_axprot = int_rd_req_desc_n_attr_axprot['h2];
assign int_rd_req_desc_2_attr_axcache = int_rd_req_desc_n_attr_axcache['h2];
assign int_rd_req_desc_2_attr_axlock = int_rd_req_desc_n_attr_axlock['h2];
assign int_rd_req_desc_2_attr_axburst = int_rd_req_desc_n_attr_axburst['h2];
assign int_rd_req_desc_2_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h2];
assign int_rd_req_desc_2_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h2];
assign int_rd_req_desc_2_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h2];
assign int_rd_req_desc_2_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h2];
assign int_rd_req_desc_2_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h2];
assign int_rd_req_desc_2_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h2];
assign int_rd_req_desc_2_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h2];
assign int_rd_req_desc_2_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h2];
assign int_rd_req_desc_2_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h2];
assign int_rd_req_desc_2_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h2];
assign int_rd_req_desc_2_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h2];
assign int_rd_req_desc_2_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h2];
assign int_rd_req_desc_2_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h2];
assign int_rd_req_desc_2_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h2];
assign int_rd_req_desc_2_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h2];
assign int_rd_req_desc_2_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h2];
assign int_rd_req_desc_2_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h2];
assign int_rd_req_desc_2_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h2];
assign int_rd_req_desc_2_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h2];
assign int_rd_req_desc_2_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h2];
assign int_rd_req_desc_2_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h2];
assign int_rd_req_desc_2_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h2];
assign int_rd_req_desc_2_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h2];
assign int_rd_req_desc_2_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h2];
assign int_wr_req_desc_2_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h2];
assign int_wr_req_desc_2_size_txn_size = int_wr_req_desc_n_size_txn_size['h2];
assign int_wr_req_desc_2_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h2];
assign int_wr_req_desc_2_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h2];
assign int_wr_req_desc_2_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h2];
assign int_wr_req_desc_2_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h2];
assign int_wr_req_desc_2_attr_axbar = int_wr_req_desc_n_attr_axbar['h2];
assign int_wr_req_desc_2_attr_awunique = int_wr_req_desc_n_attr_awunique['h2];
assign int_wr_req_desc_2_attr_axregion = int_wr_req_desc_n_attr_axregion['h2];
assign int_wr_req_desc_2_attr_axqos = int_wr_req_desc_n_attr_axqos['h2];
assign int_wr_req_desc_2_attr_axprot = int_wr_req_desc_n_attr_axprot['h2];
assign int_wr_req_desc_2_attr_axcache = int_wr_req_desc_n_attr_axcache['h2];
assign int_wr_req_desc_2_attr_axlock = int_wr_req_desc_n_attr_axlock['h2];
assign int_wr_req_desc_2_attr_axburst = int_wr_req_desc_n_attr_axburst['h2];
assign int_wr_req_desc_2_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h2];
assign int_wr_req_desc_2_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h2];
assign int_wr_req_desc_2_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h2];
assign int_wr_req_desc_2_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h2];
assign int_wr_req_desc_2_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h2];
assign int_wr_req_desc_2_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h2];
assign int_wr_req_desc_2_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h2];
assign int_wr_req_desc_2_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h2];
assign int_wr_req_desc_2_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h2];
assign int_wr_req_desc_2_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h2];
assign int_wr_req_desc_2_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h2];
assign int_wr_req_desc_2_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h2];
assign int_wr_req_desc_2_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h2];
assign int_wr_req_desc_2_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h2];
assign int_wr_req_desc_2_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h2];
assign int_wr_req_desc_2_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h2];
assign int_wr_req_desc_2_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h2];
assign int_wr_req_desc_2_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h2];
assign int_wr_req_desc_2_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h2];
assign int_wr_req_desc_2_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h2];
assign int_wr_req_desc_2_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h2];
assign int_wr_req_desc_2_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h2];
assign int_wr_req_desc_2_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h2];
assign int_wr_req_desc_2_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h2];
assign int_wr_req_desc_2_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h2];
assign int_wr_req_desc_2_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h2];
assign int_wr_req_desc_2_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h2];
assign int_wr_req_desc_2_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h2];
assign int_wr_req_desc_2_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h2];
assign int_wr_req_desc_2_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h2];
assign int_wr_req_desc_2_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h2];
assign int_wr_req_desc_2_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h2];
assign int_wr_req_desc_2_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h2];
assign int_wr_req_desc_2_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h2];
assign int_wr_req_desc_2_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h2];
assign int_wr_req_desc_2_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h2];
assign int_wr_req_desc_2_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h2];
assign int_wr_req_desc_2_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h2];
assign int_wr_req_desc_2_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h2];
assign int_wr_req_desc_2_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h2];
assign int_sn_resp_desc_2_resp_resp = int_sn_resp_desc_n_resp_resp['h2];
assign int_rd_req_desc_3_size_txn_size = int_rd_req_desc_n_size_txn_size['h3];
assign int_rd_req_desc_3_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h3];
assign int_rd_req_desc_3_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h3];
assign int_rd_req_desc_3_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h3];
assign int_rd_req_desc_3_attr_axbar = int_rd_req_desc_n_attr_axbar['h3];
assign int_rd_req_desc_3_attr_axregion = int_rd_req_desc_n_attr_axregion['h3];
assign int_rd_req_desc_3_attr_axqos = int_rd_req_desc_n_attr_axqos['h3];
assign int_rd_req_desc_3_attr_axprot = int_rd_req_desc_n_attr_axprot['h3];
assign int_rd_req_desc_3_attr_axcache = int_rd_req_desc_n_attr_axcache['h3];
assign int_rd_req_desc_3_attr_axlock = int_rd_req_desc_n_attr_axlock['h3];
assign int_rd_req_desc_3_attr_axburst = int_rd_req_desc_n_attr_axburst['h3];
assign int_rd_req_desc_3_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h3];
assign int_rd_req_desc_3_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h3];
assign int_rd_req_desc_3_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h3];
assign int_rd_req_desc_3_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h3];
assign int_rd_req_desc_3_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h3];
assign int_rd_req_desc_3_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h3];
assign int_rd_req_desc_3_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h3];
assign int_rd_req_desc_3_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h3];
assign int_rd_req_desc_3_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h3];
assign int_rd_req_desc_3_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h3];
assign int_rd_req_desc_3_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h3];
assign int_rd_req_desc_3_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h3];
assign int_rd_req_desc_3_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h3];
assign int_rd_req_desc_3_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h3];
assign int_rd_req_desc_3_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h3];
assign int_rd_req_desc_3_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h3];
assign int_rd_req_desc_3_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h3];
assign int_rd_req_desc_3_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h3];
assign int_rd_req_desc_3_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h3];
assign int_rd_req_desc_3_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h3];
assign int_rd_req_desc_3_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h3];
assign int_rd_req_desc_3_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h3];
assign int_rd_req_desc_3_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h3];
assign int_rd_req_desc_3_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h3];
assign int_wr_req_desc_3_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h3];
assign int_wr_req_desc_3_size_txn_size = int_wr_req_desc_n_size_txn_size['h3];
assign int_wr_req_desc_3_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h3];
assign int_wr_req_desc_3_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h3];
assign int_wr_req_desc_3_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h3];
assign int_wr_req_desc_3_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h3];
assign int_wr_req_desc_3_attr_axbar = int_wr_req_desc_n_attr_axbar['h3];
assign int_wr_req_desc_3_attr_awunique = int_wr_req_desc_n_attr_awunique['h3];
assign int_wr_req_desc_3_attr_axregion = int_wr_req_desc_n_attr_axregion['h3];
assign int_wr_req_desc_3_attr_axqos = int_wr_req_desc_n_attr_axqos['h3];
assign int_wr_req_desc_3_attr_axprot = int_wr_req_desc_n_attr_axprot['h3];
assign int_wr_req_desc_3_attr_axcache = int_wr_req_desc_n_attr_axcache['h3];
assign int_wr_req_desc_3_attr_axlock = int_wr_req_desc_n_attr_axlock['h3];
assign int_wr_req_desc_3_attr_axburst = int_wr_req_desc_n_attr_axburst['h3];
assign int_wr_req_desc_3_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h3];
assign int_wr_req_desc_3_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h3];
assign int_wr_req_desc_3_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h3];
assign int_wr_req_desc_3_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h3];
assign int_wr_req_desc_3_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h3];
assign int_wr_req_desc_3_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h3];
assign int_wr_req_desc_3_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h3];
assign int_wr_req_desc_3_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h3];
assign int_wr_req_desc_3_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h3];
assign int_wr_req_desc_3_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h3];
assign int_wr_req_desc_3_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h3];
assign int_wr_req_desc_3_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h3];
assign int_wr_req_desc_3_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h3];
assign int_wr_req_desc_3_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h3];
assign int_wr_req_desc_3_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h3];
assign int_wr_req_desc_3_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h3];
assign int_wr_req_desc_3_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h3];
assign int_wr_req_desc_3_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h3];
assign int_wr_req_desc_3_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h3];
assign int_wr_req_desc_3_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h3];
assign int_wr_req_desc_3_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h3];
assign int_wr_req_desc_3_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h3];
assign int_wr_req_desc_3_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h3];
assign int_wr_req_desc_3_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h3];
assign int_wr_req_desc_3_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h3];
assign int_wr_req_desc_3_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h3];
assign int_wr_req_desc_3_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h3];
assign int_wr_req_desc_3_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h3];
assign int_wr_req_desc_3_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h3];
assign int_wr_req_desc_3_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h3];
assign int_wr_req_desc_3_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h3];
assign int_wr_req_desc_3_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h3];
assign int_wr_req_desc_3_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h3];
assign int_wr_req_desc_3_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h3];
assign int_wr_req_desc_3_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h3];
assign int_wr_req_desc_3_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h3];
assign int_wr_req_desc_3_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h3];
assign int_wr_req_desc_3_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h3];
assign int_wr_req_desc_3_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h3];
assign int_wr_req_desc_3_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h3];
assign int_sn_resp_desc_3_resp_resp = int_sn_resp_desc_n_resp_resp['h3];
assign int_rd_req_desc_4_size_txn_size = int_rd_req_desc_n_size_txn_size['h4];
assign int_rd_req_desc_4_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h4];
assign int_rd_req_desc_4_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h4];
assign int_rd_req_desc_4_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h4];
assign int_rd_req_desc_4_attr_axbar = int_rd_req_desc_n_attr_axbar['h4];
assign int_rd_req_desc_4_attr_axregion = int_rd_req_desc_n_attr_axregion['h4];
assign int_rd_req_desc_4_attr_axqos = int_rd_req_desc_n_attr_axqos['h4];
assign int_rd_req_desc_4_attr_axprot = int_rd_req_desc_n_attr_axprot['h4];
assign int_rd_req_desc_4_attr_axcache = int_rd_req_desc_n_attr_axcache['h4];
assign int_rd_req_desc_4_attr_axlock = int_rd_req_desc_n_attr_axlock['h4];
assign int_rd_req_desc_4_attr_axburst = int_rd_req_desc_n_attr_axburst['h4];
assign int_rd_req_desc_4_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h4];
assign int_rd_req_desc_4_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h4];
assign int_rd_req_desc_4_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h4];
assign int_rd_req_desc_4_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h4];
assign int_rd_req_desc_4_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h4];
assign int_rd_req_desc_4_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h4];
assign int_rd_req_desc_4_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h4];
assign int_rd_req_desc_4_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h4];
assign int_rd_req_desc_4_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h4];
assign int_rd_req_desc_4_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h4];
assign int_rd_req_desc_4_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h4];
assign int_rd_req_desc_4_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h4];
assign int_rd_req_desc_4_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h4];
assign int_rd_req_desc_4_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h4];
assign int_rd_req_desc_4_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h4];
assign int_rd_req_desc_4_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h4];
assign int_rd_req_desc_4_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h4];
assign int_rd_req_desc_4_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h4];
assign int_rd_req_desc_4_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h4];
assign int_rd_req_desc_4_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h4];
assign int_rd_req_desc_4_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h4];
assign int_rd_req_desc_4_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h4];
assign int_rd_req_desc_4_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h4];
assign int_rd_req_desc_4_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h4];
assign int_wr_req_desc_4_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h4];
assign int_wr_req_desc_4_size_txn_size = int_wr_req_desc_n_size_txn_size['h4];
assign int_wr_req_desc_4_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h4];
assign int_wr_req_desc_4_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h4];
assign int_wr_req_desc_4_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h4];
assign int_wr_req_desc_4_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h4];
assign int_wr_req_desc_4_attr_axbar = int_wr_req_desc_n_attr_axbar['h4];
assign int_wr_req_desc_4_attr_awunique = int_wr_req_desc_n_attr_awunique['h4];
assign int_wr_req_desc_4_attr_axregion = int_wr_req_desc_n_attr_axregion['h4];
assign int_wr_req_desc_4_attr_axqos = int_wr_req_desc_n_attr_axqos['h4];
assign int_wr_req_desc_4_attr_axprot = int_wr_req_desc_n_attr_axprot['h4];
assign int_wr_req_desc_4_attr_axcache = int_wr_req_desc_n_attr_axcache['h4];
assign int_wr_req_desc_4_attr_axlock = int_wr_req_desc_n_attr_axlock['h4];
assign int_wr_req_desc_4_attr_axburst = int_wr_req_desc_n_attr_axburst['h4];
assign int_wr_req_desc_4_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h4];
assign int_wr_req_desc_4_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h4];
assign int_wr_req_desc_4_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h4];
assign int_wr_req_desc_4_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h4];
assign int_wr_req_desc_4_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h4];
assign int_wr_req_desc_4_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h4];
assign int_wr_req_desc_4_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h4];
assign int_wr_req_desc_4_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h4];
assign int_wr_req_desc_4_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h4];
assign int_wr_req_desc_4_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h4];
assign int_wr_req_desc_4_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h4];
assign int_wr_req_desc_4_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h4];
assign int_wr_req_desc_4_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h4];
assign int_wr_req_desc_4_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h4];
assign int_wr_req_desc_4_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h4];
assign int_wr_req_desc_4_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h4];
assign int_wr_req_desc_4_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h4];
assign int_wr_req_desc_4_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h4];
assign int_wr_req_desc_4_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h4];
assign int_wr_req_desc_4_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h4];
assign int_wr_req_desc_4_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h4];
assign int_wr_req_desc_4_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h4];
assign int_wr_req_desc_4_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h4];
assign int_wr_req_desc_4_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h4];
assign int_wr_req_desc_4_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h4];
assign int_wr_req_desc_4_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h4];
assign int_wr_req_desc_4_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h4];
assign int_wr_req_desc_4_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h4];
assign int_wr_req_desc_4_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h4];
assign int_wr_req_desc_4_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h4];
assign int_wr_req_desc_4_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h4];
assign int_wr_req_desc_4_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h4];
assign int_wr_req_desc_4_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h4];
assign int_wr_req_desc_4_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h4];
assign int_wr_req_desc_4_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h4];
assign int_wr_req_desc_4_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h4];
assign int_wr_req_desc_4_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h4];
assign int_wr_req_desc_4_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h4];
assign int_wr_req_desc_4_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h4];
assign int_wr_req_desc_4_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h4];
assign int_sn_resp_desc_4_resp_resp = int_sn_resp_desc_n_resp_resp['h4];
assign int_rd_req_desc_5_size_txn_size = int_rd_req_desc_n_size_txn_size['h5];
assign int_rd_req_desc_5_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h5];
assign int_rd_req_desc_5_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h5];
assign int_rd_req_desc_5_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h5];
assign int_rd_req_desc_5_attr_axbar = int_rd_req_desc_n_attr_axbar['h5];
assign int_rd_req_desc_5_attr_axregion = int_rd_req_desc_n_attr_axregion['h5];
assign int_rd_req_desc_5_attr_axqos = int_rd_req_desc_n_attr_axqos['h5];
assign int_rd_req_desc_5_attr_axprot = int_rd_req_desc_n_attr_axprot['h5];
assign int_rd_req_desc_5_attr_axcache = int_rd_req_desc_n_attr_axcache['h5];
assign int_rd_req_desc_5_attr_axlock = int_rd_req_desc_n_attr_axlock['h5];
assign int_rd_req_desc_5_attr_axburst = int_rd_req_desc_n_attr_axburst['h5];
assign int_rd_req_desc_5_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h5];
assign int_rd_req_desc_5_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h5];
assign int_rd_req_desc_5_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h5];
assign int_rd_req_desc_5_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h5];
assign int_rd_req_desc_5_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h5];
assign int_rd_req_desc_5_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h5];
assign int_rd_req_desc_5_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h5];
assign int_rd_req_desc_5_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h5];
assign int_rd_req_desc_5_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h5];
assign int_rd_req_desc_5_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h5];
assign int_rd_req_desc_5_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h5];
assign int_rd_req_desc_5_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h5];
assign int_rd_req_desc_5_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h5];
assign int_rd_req_desc_5_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h5];
assign int_rd_req_desc_5_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h5];
assign int_rd_req_desc_5_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h5];
assign int_rd_req_desc_5_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h5];
assign int_rd_req_desc_5_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h5];
assign int_rd_req_desc_5_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h5];
assign int_rd_req_desc_5_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h5];
assign int_rd_req_desc_5_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h5];
assign int_rd_req_desc_5_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h5];
assign int_rd_req_desc_5_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h5];
assign int_rd_req_desc_5_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h5];
assign int_wr_req_desc_5_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h5];
assign int_wr_req_desc_5_size_txn_size = int_wr_req_desc_n_size_txn_size['h5];
assign int_wr_req_desc_5_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h5];
assign int_wr_req_desc_5_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h5];
assign int_wr_req_desc_5_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h5];
assign int_wr_req_desc_5_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h5];
assign int_wr_req_desc_5_attr_axbar = int_wr_req_desc_n_attr_axbar['h5];
assign int_wr_req_desc_5_attr_awunique = int_wr_req_desc_n_attr_awunique['h5];
assign int_wr_req_desc_5_attr_axregion = int_wr_req_desc_n_attr_axregion['h5];
assign int_wr_req_desc_5_attr_axqos = int_wr_req_desc_n_attr_axqos['h5];
assign int_wr_req_desc_5_attr_axprot = int_wr_req_desc_n_attr_axprot['h5];
assign int_wr_req_desc_5_attr_axcache = int_wr_req_desc_n_attr_axcache['h5];
assign int_wr_req_desc_5_attr_axlock = int_wr_req_desc_n_attr_axlock['h5];
assign int_wr_req_desc_5_attr_axburst = int_wr_req_desc_n_attr_axburst['h5];
assign int_wr_req_desc_5_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h5];
assign int_wr_req_desc_5_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h5];
assign int_wr_req_desc_5_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h5];
assign int_wr_req_desc_5_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h5];
assign int_wr_req_desc_5_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h5];
assign int_wr_req_desc_5_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h5];
assign int_wr_req_desc_5_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h5];
assign int_wr_req_desc_5_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h5];
assign int_wr_req_desc_5_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h5];
assign int_wr_req_desc_5_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h5];
assign int_wr_req_desc_5_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h5];
assign int_wr_req_desc_5_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h5];
assign int_wr_req_desc_5_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h5];
assign int_wr_req_desc_5_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h5];
assign int_wr_req_desc_5_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h5];
assign int_wr_req_desc_5_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h5];
assign int_wr_req_desc_5_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h5];
assign int_wr_req_desc_5_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h5];
assign int_wr_req_desc_5_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h5];
assign int_wr_req_desc_5_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h5];
assign int_wr_req_desc_5_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h5];
assign int_wr_req_desc_5_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h5];
assign int_wr_req_desc_5_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h5];
assign int_wr_req_desc_5_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h5];
assign int_wr_req_desc_5_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h5];
assign int_wr_req_desc_5_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h5];
assign int_wr_req_desc_5_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h5];
assign int_wr_req_desc_5_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h5];
assign int_wr_req_desc_5_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h5];
assign int_wr_req_desc_5_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h5];
assign int_wr_req_desc_5_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h5];
assign int_wr_req_desc_5_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h5];
assign int_wr_req_desc_5_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h5];
assign int_wr_req_desc_5_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h5];
assign int_wr_req_desc_5_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h5];
assign int_wr_req_desc_5_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h5];
assign int_wr_req_desc_5_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h5];
assign int_wr_req_desc_5_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h5];
assign int_wr_req_desc_5_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h5];
assign int_wr_req_desc_5_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h5];
assign int_sn_resp_desc_5_resp_resp = int_sn_resp_desc_n_resp_resp['h5];
assign int_rd_req_desc_6_size_txn_size = int_rd_req_desc_n_size_txn_size['h6];
assign int_rd_req_desc_6_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h6];
assign int_rd_req_desc_6_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h6];
assign int_rd_req_desc_6_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h6];
assign int_rd_req_desc_6_attr_axbar = int_rd_req_desc_n_attr_axbar['h6];
assign int_rd_req_desc_6_attr_axregion = int_rd_req_desc_n_attr_axregion['h6];
assign int_rd_req_desc_6_attr_axqos = int_rd_req_desc_n_attr_axqos['h6];
assign int_rd_req_desc_6_attr_axprot = int_rd_req_desc_n_attr_axprot['h6];
assign int_rd_req_desc_6_attr_axcache = int_rd_req_desc_n_attr_axcache['h6];
assign int_rd_req_desc_6_attr_axlock = int_rd_req_desc_n_attr_axlock['h6];
assign int_rd_req_desc_6_attr_axburst = int_rd_req_desc_n_attr_axburst['h6];
assign int_rd_req_desc_6_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h6];
assign int_rd_req_desc_6_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h6];
assign int_rd_req_desc_6_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h6];
assign int_rd_req_desc_6_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h6];
assign int_rd_req_desc_6_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h6];
assign int_rd_req_desc_6_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h6];
assign int_rd_req_desc_6_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h6];
assign int_rd_req_desc_6_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h6];
assign int_rd_req_desc_6_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h6];
assign int_rd_req_desc_6_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h6];
assign int_rd_req_desc_6_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h6];
assign int_rd_req_desc_6_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h6];
assign int_rd_req_desc_6_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h6];
assign int_rd_req_desc_6_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h6];
assign int_rd_req_desc_6_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h6];
assign int_rd_req_desc_6_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h6];
assign int_rd_req_desc_6_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h6];
assign int_rd_req_desc_6_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h6];
assign int_rd_req_desc_6_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h6];
assign int_rd_req_desc_6_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h6];
assign int_rd_req_desc_6_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h6];
assign int_rd_req_desc_6_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h6];
assign int_rd_req_desc_6_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h6];
assign int_rd_req_desc_6_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h6];
assign int_wr_req_desc_6_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h6];
assign int_wr_req_desc_6_size_txn_size = int_wr_req_desc_n_size_txn_size['h6];
assign int_wr_req_desc_6_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h6];
assign int_wr_req_desc_6_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h6];
assign int_wr_req_desc_6_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h6];
assign int_wr_req_desc_6_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h6];
assign int_wr_req_desc_6_attr_axbar = int_wr_req_desc_n_attr_axbar['h6];
assign int_wr_req_desc_6_attr_awunique = int_wr_req_desc_n_attr_awunique['h6];
assign int_wr_req_desc_6_attr_axregion = int_wr_req_desc_n_attr_axregion['h6];
assign int_wr_req_desc_6_attr_axqos = int_wr_req_desc_n_attr_axqos['h6];
assign int_wr_req_desc_6_attr_axprot = int_wr_req_desc_n_attr_axprot['h6];
assign int_wr_req_desc_6_attr_axcache = int_wr_req_desc_n_attr_axcache['h6];
assign int_wr_req_desc_6_attr_axlock = int_wr_req_desc_n_attr_axlock['h6];
assign int_wr_req_desc_6_attr_axburst = int_wr_req_desc_n_attr_axburst['h6];
assign int_wr_req_desc_6_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h6];
assign int_wr_req_desc_6_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h6];
assign int_wr_req_desc_6_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h6];
assign int_wr_req_desc_6_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h6];
assign int_wr_req_desc_6_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h6];
assign int_wr_req_desc_6_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h6];
assign int_wr_req_desc_6_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h6];
assign int_wr_req_desc_6_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h6];
assign int_wr_req_desc_6_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h6];
assign int_wr_req_desc_6_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h6];
assign int_wr_req_desc_6_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h6];
assign int_wr_req_desc_6_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h6];
assign int_wr_req_desc_6_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h6];
assign int_wr_req_desc_6_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h6];
assign int_wr_req_desc_6_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h6];
assign int_wr_req_desc_6_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h6];
assign int_wr_req_desc_6_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h6];
assign int_wr_req_desc_6_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h6];
assign int_wr_req_desc_6_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h6];
assign int_wr_req_desc_6_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h6];
assign int_wr_req_desc_6_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h6];
assign int_wr_req_desc_6_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h6];
assign int_wr_req_desc_6_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h6];
assign int_wr_req_desc_6_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h6];
assign int_wr_req_desc_6_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h6];
assign int_wr_req_desc_6_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h6];
assign int_wr_req_desc_6_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h6];
assign int_wr_req_desc_6_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h6];
assign int_wr_req_desc_6_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h6];
assign int_wr_req_desc_6_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h6];
assign int_wr_req_desc_6_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h6];
assign int_wr_req_desc_6_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h6];
assign int_wr_req_desc_6_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h6];
assign int_wr_req_desc_6_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h6];
assign int_wr_req_desc_6_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h6];
assign int_wr_req_desc_6_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h6];
assign int_wr_req_desc_6_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h6];
assign int_wr_req_desc_6_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h6];
assign int_wr_req_desc_6_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h6];
assign int_wr_req_desc_6_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h6];
assign int_sn_resp_desc_6_resp_resp = int_sn_resp_desc_n_resp_resp['h6];
assign int_rd_req_desc_7_size_txn_size = int_rd_req_desc_n_size_txn_size['h7];
assign int_rd_req_desc_7_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h7];
assign int_rd_req_desc_7_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h7];
assign int_rd_req_desc_7_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h7];
assign int_rd_req_desc_7_attr_axbar = int_rd_req_desc_n_attr_axbar['h7];
assign int_rd_req_desc_7_attr_axregion = int_rd_req_desc_n_attr_axregion['h7];
assign int_rd_req_desc_7_attr_axqos = int_rd_req_desc_n_attr_axqos['h7];
assign int_rd_req_desc_7_attr_axprot = int_rd_req_desc_n_attr_axprot['h7];
assign int_rd_req_desc_7_attr_axcache = int_rd_req_desc_n_attr_axcache['h7];
assign int_rd_req_desc_7_attr_axlock = int_rd_req_desc_n_attr_axlock['h7];
assign int_rd_req_desc_7_attr_axburst = int_rd_req_desc_n_attr_axburst['h7];
assign int_rd_req_desc_7_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h7];
assign int_rd_req_desc_7_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h7];
assign int_rd_req_desc_7_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h7];
assign int_rd_req_desc_7_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h7];
assign int_rd_req_desc_7_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h7];
assign int_rd_req_desc_7_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h7];
assign int_rd_req_desc_7_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h7];
assign int_rd_req_desc_7_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h7];
assign int_rd_req_desc_7_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h7];
assign int_rd_req_desc_7_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h7];
assign int_rd_req_desc_7_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h7];
assign int_rd_req_desc_7_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h7];
assign int_rd_req_desc_7_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h7];
assign int_rd_req_desc_7_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h7];
assign int_rd_req_desc_7_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h7];
assign int_rd_req_desc_7_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h7];
assign int_rd_req_desc_7_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h7];
assign int_rd_req_desc_7_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h7];
assign int_rd_req_desc_7_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h7];
assign int_rd_req_desc_7_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h7];
assign int_rd_req_desc_7_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h7];
assign int_rd_req_desc_7_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h7];
assign int_rd_req_desc_7_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h7];
assign int_rd_req_desc_7_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h7];
assign int_wr_req_desc_7_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h7];
assign int_wr_req_desc_7_size_txn_size = int_wr_req_desc_n_size_txn_size['h7];
assign int_wr_req_desc_7_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h7];
assign int_wr_req_desc_7_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h7];
assign int_wr_req_desc_7_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h7];
assign int_wr_req_desc_7_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h7];
assign int_wr_req_desc_7_attr_axbar = int_wr_req_desc_n_attr_axbar['h7];
assign int_wr_req_desc_7_attr_awunique = int_wr_req_desc_n_attr_awunique['h7];
assign int_wr_req_desc_7_attr_axregion = int_wr_req_desc_n_attr_axregion['h7];
assign int_wr_req_desc_7_attr_axqos = int_wr_req_desc_n_attr_axqos['h7];
assign int_wr_req_desc_7_attr_axprot = int_wr_req_desc_n_attr_axprot['h7];
assign int_wr_req_desc_7_attr_axcache = int_wr_req_desc_n_attr_axcache['h7];
assign int_wr_req_desc_7_attr_axlock = int_wr_req_desc_n_attr_axlock['h7];
assign int_wr_req_desc_7_attr_axburst = int_wr_req_desc_n_attr_axburst['h7];
assign int_wr_req_desc_7_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h7];
assign int_wr_req_desc_7_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h7];
assign int_wr_req_desc_7_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h7];
assign int_wr_req_desc_7_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h7];
assign int_wr_req_desc_7_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h7];
assign int_wr_req_desc_7_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h7];
assign int_wr_req_desc_7_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h7];
assign int_wr_req_desc_7_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h7];
assign int_wr_req_desc_7_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h7];
assign int_wr_req_desc_7_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h7];
assign int_wr_req_desc_7_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h7];
assign int_wr_req_desc_7_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h7];
assign int_wr_req_desc_7_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h7];
assign int_wr_req_desc_7_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h7];
assign int_wr_req_desc_7_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h7];
assign int_wr_req_desc_7_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h7];
assign int_wr_req_desc_7_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h7];
assign int_wr_req_desc_7_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h7];
assign int_wr_req_desc_7_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h7];
assign int_wr_req_desc_7_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h7];
assign int_wr_req_desc_7_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h7];
assign int_wr_req_desc_7_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h7];
assign int_wr_req_desc_7_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h7];
assign int_wr_req_desc_7_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h7];
assign int_wr_req_desc_7_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h7];
assign int_wr_req_desc_7_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h7];
assign int_wr_req_desc_7_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h7];
assign int_wr_req_desc_7_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h7];
assign int_wr_req_desc_7_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h7];
assign int_wr_req_desc_7_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h7];
assign int_wr_req_desc_7_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h7];
assign int_wr_req_desc_7_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h7];
assign int_wr_req_desc_7_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h7];
assign int_wr_req_desc_7_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h7];
assign int_wr_req_desc_7_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h7];
assign int_wr_req_desc_7_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h7];
assign int_wr_req_desc_7_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h7];
assign int_wr_req_desc_7_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h7];
assign int_wr_req_desc_7_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h7];
assign int_wr_req_desc_7_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h7];
assign int_sn_resp_desc_7_resp_resp = int_sn_resp_desc_n_resp_resp['h7];
assign int_rd_req_desc_8_size_txn_size = int_rd_req_desc_n_size_txn_size['h8];
assign int_rd_req_desc_8_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h8];
assign int_rd_req_desc_8_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h8];
assign int_rd_req_desc_8_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h8];
assign int_rd_req_desc_8_attr_axbar = int_rd_req_desc_n_attr_axbar['h8];
assign int_rd_req_desc_8_attr_axregion = int_rd_req_desc_n_attr_axregion['h8];
assign int_rd_req_desc_8_attr_axqos = int_rd_req_desc_n_attr_axqos['h8];
assign int_rd_req_desc_8_attr_axprot = int_rd_req_desc_n_attr_axprot['h8];
assign int_rd_req_desc_8_attr_axcache = int_rd_req_desc_n_attr_axcache['h8];
assign int_rd_req_desc_8_attr_axlock = int_rd_req_desc_n_attr_axlock['h8];
assign int_rd_req_desc_8_attr_axburst = int_rd_req_desc_n_attr_axburst['h8];
assign int_rd_req_desc_8_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h8];
assign int_rd_req_desc_8_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h8];
assign int_rd_req_desc_8_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h8];
assign int_rd_req_desc_8_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h8];
assign int_rd_req_desc_8_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h8];
assign int_rd_req_desc_8_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h8];
assign int_rd_req_desc_8_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h8];
assign int_rd_req_desc_8_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h8];
assign int_rd_req_desc_8_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h8];
assign int_rd_req_desc_8_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h8];
assign int_rd_req_desc_8_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h8];
assign int_rd_req_desc_8_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h8];
assign int_rd_req_desc_8_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h8];
assign int_rd_req_desc_8_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h8];
assign int_rd_req_desc_8_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h8];
assign int_rd_req_desc_8_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h8];
assign int_rd_req_desc_8_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h8];
assign int_rd_req_desc_8_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h8];
assign int_rd_req_desc_8_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h8];
assign int_rd_req_desc_8_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h8];
assign int_rd_req_desc_8_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h8];
assign int_rd_req_desc_8_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h8];
assign int_rd_req_desc_8_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h8];
assign int_rd_req_desc_8_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h8];
assign int_wr_req_desc_8_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h8];
assign int_wr_req_desc_8_size_txn_size = int_wr_req_desc_n_size_txn_size['h8];
assign int_wr_req_desc_8_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h8];
assign int_wr_req_desc_8_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h8];
assign int_wr_req_desc_8_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h8];
assign int_wr_req_desc_8_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h8];
assign int_wr_req_desc_8_attr_axbar = int_wr_req_desc_n_attr_axbar['h8];
assign int_wr_req_desc_8_attr_awunique = int_wr_req_desc_n_attr_awunique['h8];
assign int_wr_req_desc_8_attr_axregion = int_wr_req_desc_n_attr_axregion['h8];
assign int_wr_req_desc_8_attr_axqos = int_wr_req_desc_n_attr_axqos['h8];
assign int_wr_req_desc_8_attr_axprot = int_wr_req_desc_n_attr_axprot['h8];
assign int_wr_req_desc_8_attr_axcache = int_wr_req_desc_n_attr_axcache['h8];
assign int_wr_req_desc_8_attr_axlock = int_wr_req_desc_n_attr_axlock['h8];
assign int_wr_req_desc_8_attr_axburst = int_wr_req_desc_n_attr_axburst['h8];
assign int_wr_req_desc_8_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h8];
assign int_wr_req_desc_8_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h8];
assign int_wr_req_desc_8_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h8];
assign int_wr_req_desc_8_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h8];
assign int_wr_req_desc_8_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h8];
assign int_wr_req_desc_8_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h8];
assign int_wr_req_desc_8_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h8];
assign int_wr_req_desc_8_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h8];
assign int_wr_req_desc_8_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h8];
assign int_wr_req_desc_8_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h8];
assign int_wr_req_desc_8_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h8];
assign int_wr_req_desc_8_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h8];
assign int_wr_req_desc_8_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h8];
assign int_wr_req_desc_8_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h8];
assign int_wr_req_desc_8_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h8];
assign int_wr_req_desc_8_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h8];
assign int_wr_req_desc_8_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h8];
assign int_wr_req_desc_8_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h8];
assign int_wr_req_desc_8_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h8];
assign int_wr_req_desc_8_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h8];
assign int_wr_req_desc_8_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h8];
assign int_wr_req_desc_8_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h8];
assign int_wr_req_desc_8_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h8];
assign int_wr_req_desc_8_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h8];
assign int_wr_req_desc_8_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h8];
assign int_wr_req_desc_8_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h8];
assign int_wr_req_desc_8_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h8];
assign int_wr_req_desc_8_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h8];
assign int_wr_req_desc_8_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h8];
assign int_wr_req_desc_8_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h8];
assign int_wr_req_desc_8_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h8];
assign int_wr_req_desc_8_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h8];
assign int_wr_req_desc_8_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h8];
assign int_wr_req_desc_8_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h8];
assign int_wr_req_desc_8_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h8];
assign int_wr_req_desc_8_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h8];
assign int_wr_req_desc_8_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h8];
assign int_wr_req_desc_8_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h8];
assign int_wr_req_desc_8_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h8];
assign int_wr_req_desc_8_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h8];
assign int_sn_resp_desc_8_resp_resp = int_sn_resp_desc_n_resp_resp['h8];
assign int_rd_req_desc_9_size_txn_size = int_rd_req_desc_n_size_txn_size['h9];
assign int_rd_req_desc_9_axsize_axsize = int_rd_req_desc_n_axsize_axsize['h9];
assign int_rd_req_desc_9_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['h9];
assign int_rd_req_desc_9_attr_axdomain = int_rd_req_desc_n_attr_axdomain['h9];
assign int_rd_req_desc_9_attr_axbar = int_rd_req_desc_n_attr_axbar['h9];
assign int_rd_req_desc_9_attr_axregion = int_rd_req_desc_n_attr_axregion['h9];
assign int_rd_req_desc_9_attr_axqos = int_rd_req_desc_n_attr_axqos['h9];
assign int_rd_req_desc_9_attr_axprot = int_rd_req_desc_n_attr_axprot['h9];
assign int_rd_req_desc_9_attr_axcache = int_rd_req_desc_n_attr_axcache['h9];
assign int_rd_req_desc_9_attr_axlock = int_rd_req_desc_n_attr_axlock['h9];
assign int_rd_req_desc_9_attr_axburst = int_rd_req_desc_n_attr_axburst['h9];
assign int_rd_req_desc_9_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['h9];
assign int_rd_req_desc_9_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['h9];
assign int_rd_req_desc_9_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['h9];
assign int_rd_req_desc_9_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['h9];
assign int_rd_req_desc_9_axid_0_axid = int_rd_req_desc_n_axid_0_axid['h9];
assign int_rd_req_desc_9_axid_1_axid = int_rd_req_desc_n_axid_1_axid['h9];
assign int_rd_req_desc_9_axid_2_axid = int_rd_req_desc_n_axid_2_axid['h9];
assign int_rd_req_desc_9_axid_3_axid = int_rd_req_desc_n_axid_3_axid['h9];
assign int_rd_req_desc_9_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['h9];
assign int_rd_req_desc_9_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['h9];
assign int_rd_req_desc_9_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['h9];
assign int_rd_req_desc_9_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['h9];
assign int_rd_req_desc_9_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['h9];
assign int_rd_req_desc_9_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['h9];
assign int_rd_req_desc_9_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['h9];
assign int_rd_req_desc_9_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['h9];
assign int_rd_req_desc_9_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['h9];
assign int_rd_req_desc_9_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['h9];
assign int_rd_req_desc_9_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['h9];
assign int_rd_req_desc_9_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['h9];
assign int_rd_req_desc_9_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['h9];
assign int_rd_req_desc_9_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['h9];
assign int_rd_req_desc_9_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['h9];
assign int_rd_req_desc_9_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['h9];
assign int_wr_req_desc_9_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['h9];
assign int_wr_req_desc_9_size_txn_size = int_wr_req_desc_n_size_txn_size['h9];
assign int_wr_req_desc_9_data_offset_addr = int_wr_req_desc_n_data_offset_addr['h9];
assign int_wr_req_desc_9_axsize_axsize = int_wr_req_desc_n_axsize_axsize['h9];
assign int_wr_req_desc_9_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['h9];
assign int_wr_req_desc_9_attr_axdomain = int_wr_req_desc_n_attr_axdomain['h9];
assign int_wr_req_desc_9_attr_axbar = int_wr_req_desc_n_attr_axbar['h9];
assign int_wr_req_desc_9_attr_awunique = int_wr_req_desc_n_attr_awunique['h9];
assign int_wr_req_desc_9_attr_axregion = int_wr_req_desc_n_attr_axregion['h9];
assign int_wr_req_desc_9_attr_axqos = int_wr_req_desc_n_attr_axqos['h9];
assign int_wr_req_desc_9_attr_axprot = int_wr_req_desc_n_attr_axprot['h9];
assign int_wr_req_desc_9_attr_axcache = int_wr_req_desc_n_attr_axcache['h9];
assign int_wr_req_desc_9_attr_axlock = int_wr_req_desc_n_attr_axlock['h9];
assign int_wr_req_desc_9_attr_axburst = int_wr_req_desc_n_attr_axburst['h9];
assign int_wr_req_desc_9_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['h9];
assign int_wr_req_desc_9_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['h9];
assign int_wr_req_desc_9_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['h9];
assign int_wr_req_desc_9_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['h9];
assign int_wr_req_desc_9_axid_0_axid = int_wr_req_desc_n_axid_0_axid['h9];
assign int_wr_req_desc_9_axid_1_axid = int_wr_req_desc_n_axid_1_axid['h9];
assign int_wr_req_desc_9_axid_2_axid = int_wr_req_desc_n_axid_2_axid['h9];
assign int_wr_req_desc_9_axid_3_axid = int_wr_req_desc_n_axid_3_axid['h9];
assign int_wr_req_desc_9_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['h9];
assign int_wr_req_desc_9_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['h9];
assign int_wr_req_desc_9_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['h9];
assign int_wr_req_desc_9_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['h9];
assign int_wr_req_desc_9_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['h9];
assign int_wr_req_desc_9_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['h9];
assign int_wr_req_desc_9_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['h9];
assign int_wr_req_desc_9_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['h9];
assign int_wr_req_desc_9_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['h9];
assign int_wr_req_desc_9_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['h9];
assign int_wr_req_desc_9_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['h9];
assign int_wr_req_desc_9_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['h9];
assign int_wr_req_desc_9_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['h9];
assign int_wr_req_desc_9_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['h9];
assign int_wr_req_desc_9_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['h9];
assign int_wr_req_desc_9_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['h9];
assign int_wr_req_desc_9_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['h9];
assign int_wr_req_desc_9_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['h9];
assign int_wr_req_desc_9_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['h9];
assign int_wr_req_desc_9_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['h9];
assign int_wr_req_desc_9_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['h9];
assign int_wr_req_desc_9_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['h9];
assign int_wr_req_desc_9_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['h9];
assign int_wr_req_desc_9_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['h9];
assign int_wr_req_desc_9_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['h9];
assign int_wr_req_desc_9_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['h9];
assign int_wr_req_desc_9_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['h9];
assign int_wr_req_desc_9_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['h9];
assign int_wr_req_desc_9_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['h9];
assign int_wr_req_desc_9_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['h9];
assign int_wr_req_desc_9_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['h9];
assign int_wr_req_desc_9_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['h9];
assign int_sn_resp_desc_9_resp_resp = int_sn_resp_desc_n_resp_resp['h9];
assign int_rd_req_desc_a_size_txn_size = int_rd_req_desc_n_size_txn_size['ha];
assign int_rd_req_desc_a_axsize_axsize = int_rd_req_desc_n_axsize_axsize['ha];
assign int_rd_req_desc_a_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['ha];
assign int_rd_req_desc_a_attr_axdomain = int_rd_req_desc_n_attr_axdomain['ha];
assign int_rd_req_desc_a_attr_axbar = int_rd_req_desc_n_attr_axbar['ha];
assign int_rd_req_desc_a_attr_axregion = int_rd_req_desc_n_attr_axregion['ha];
assign int_rd_req_desc_a_attr_axqos = int_rd_req_desc_n_attr_axqos['ha];
assign int_rd_req_desc_a_attr_axprot = int_rd_req_desc_n_attr_axprot['ha];
assign int_rd_req_desc_a_attr_axcache = int_rd_req_desc_n_attr_axcache['ha];
assign int_rd_req_desc_a_attr_axlock = int_rd_req_desc_n_attr_axlock['ha];
assign int_rd_req_desc_a_attr_axburst = int_rd_req_desc_n_attr_axburst['ha];
assign int_rd_req_desc_a_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['ha];
assign int_rd_req_desc_a_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['ha];
assign int_rd_req_desc_a_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['ha];
assign int_rd_req_desc_a_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['ha];
assign int_rd_req_desc_a_axid_0_axid = int_rd_req_desc_n_axid_0_axid['ha];
assign int_rd_req_desc_a_axid_1_axid = int_rd_req_desc_n_axid_1_axid['ha];
assign int_rd_req_desc_a_axid_2_axid = int_rd_req_desc_n_axid_2_axid['ha];
assign int_rd_req_desc_a_axid_3_axid = int_rd_req_desc_n_axid_3_axid['ha];
assign int_rd_req_desc_a_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['ha];
assign int_rd_req_desc_a_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['ha];
assign int_rd_req_desc_a_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['ha];
assign int_rd_req_desc_a_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['ha];
assign int_rd_req_desc_a_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['ha];
assign int_rd_req_desc_a_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['ha];
assign int_rd_req_desc_a_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['ha];
assign int_rd_req_desc_a_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['ha];
assign int_rd_req_desc_a_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['ha];
assign int_rd_req_desc_a_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['ha];
assign int_rd_req_desc_a_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['ha];
assign int_rd_req_desc_a_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['ha];
assign int_rd_req_desc_a_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['ha];
assign int_rd_req_desc_a_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['ha];
assign int_rd_req_desc_a_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['ha];
assign int_rd_req_desc_a_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['ha];
assign int_wr_req_desc_a_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['ha];
assign int_wr_req_desc_a_size_txn_size = int_wr_req_desc_n_size_txn_size['ha];
assign int_wr_req_desc_a_data_offset_addr = int_wr_req_desc_n_data_offset_addr['ha];
assign int_wr_req_desc_a_axsize_axsize = int_wr_req_desc_n_axsize_axsize['ha];
assign int_wr_req_desc_a_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['ha];
assign int_wr_req_desc_a_attr_axdomain = int_wr_req_desc_n_attr_axdomain['ha];
assign int_wr_req_desc_a_attr_axbar = int_wr_req_desc_n_attr_axbar['ha];
assign int_wr_req_desc_a_attr_awunique = int_wr_req_desc_n_attr_awunique['ha];
assign int_wr_req_desc_a_attr_axregion = int_wr_req_desc_n_attr_axregion['ha];
assign int_wr_req_desc_a_attr_axqos = int_wr_req_desc_n_attr_axqos['ha];
assign int_wr_req_desc_a_attr_axprot = int_wr_req_desc_n_attr_axprot['ha];
assign int_wr_req_desc_a_attr_axcache = int_wr_req_desc_n_attr_axcache['ha];
assign int_wr_req_desc_a_attr_axlock = int_wr_req_desc_n_attr_axlock['ha];
assign int_wr_req_desc_a_attr_axburst = int_wr_req_desc_n_attr_axburst['ha];
assign int_wr_req_desc_a_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['ha];
assign int_wr_req_desc_a_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['ha];
assign int_wr_req_desc_a_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['ha];
assign int_wr_req_desc_a_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['ha];
assign int_wr_req_desc_a_axid_0_axid = int_wr_req_desc_n_axid_0_axid['ha];
assign int_wr_req_desc_a_axid_1_axid = int_wr_req_desc_n_axid_1_axid['ha];
assign int_wr_req_desc_a_axid_2_axid = int_wr_req_desc_n_axid_2_axid['ha];
assign int_wr_req_desc_a_axid_3_axid = int_wr_req_desc_n_axid_3_axid['ha];
assign int_wr_req_desc_a_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['ha];
assign int_wr_req_desc_a_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['ha];
assign int_wr_req_desc_a_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['ha];
assign int_wr_req_desc_a_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['ha];
assign int_wr_req_desc_a_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['ha];
assign int_wr_req_desc_a_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['ha];
assign int_wr_req_desc_a_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['ha];
assign int_wr_req_desc_a_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['ha];
assign int_wr_req_desc_a_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['ha];
assign int_wr_req_desc_a_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['ha];
assign int_wr_req_desc_a_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['ha];
assign int_wr_req_desc_a_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['ha];
assign int_wr_req_desc_a_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['ha];
assign int_wr_req_desc_a_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['ha];
assign int_wr_req_desc_a_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['ha];
assign int_wr_req_desc_a_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['ha];
assign int_wr_req_desc_a_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['ha];
assign int_wr_req_desc_a_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['ha];
assign int_wr_req_desc_a_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['ha];
assign int_wr_req_desc_a_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['ha];
assign int_wr_req_desc_a_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['ha];
assign int_wr_req_desc_a_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['ha];
assign int_wr_req_desc_a_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['ha];
assign int_wr_req_desc_a_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['ha];
assign int_wr_req_desc_a_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['ha];
assign int_wr_req_desc_a_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['ha];
assign int_wr_req_desc_a_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['ha];
assign int_wr_req_desc_a_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['ha];
assign int_wr_req_desc_a_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['ha];
assign int_wr_req_desc_a_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['ha];
assign int_wr_req_desc_a_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['ha];
assign int_wr_req_desc_a_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['ha];
assign int_sn_resp_desc_a_resp_resp = int_sn_resp_desc_n_resp_resp['ha];
assign int_rd_req_desc_b_size_txn_size = int_rd_req_desc_n_size_txn_size['hb];
assign int_rd_req_desc_b_axsize_axsize = int_rd_req_desc_n_axsize_axsize['hb];
assign int_rd_req_desc_b_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['hb];
assign int_rd_req_desc_b_attr_axdomain = int_rd_req_desc_n_attr_axdomain['hb];
assign int_rd_req_desc_b_attr_axbar = int_rd_req_desc_n_attr_axbar['hb];
assign int_rd_req_desc_b_attr_axregion = int_rd_req_desc_n_attr_axregion['hb];
assign int_rd_req_desc_b_attr_axqos = int_rd_req_desc_n_attr_axqos['hb];
assign int_rd_req_desc_b_attr_axprot = int_rd_req_desc_n_attr_axprot['hb];
assign int_rd_req_desc_b_attr_axcache = int_rd_req_desc_n_attr_axcache['hb];
assign int_rd_req_desc_b_attr_axlock = int_rd_req_desc_n_attr_axlock['hb];
assign int_rd_req_desc_b_attr_axburst = int_rd_req_desc_n_attr_axburst['hb];
assign int_rd_req_desc_b_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['hb];
assign int_rd_req_desc_b_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['hb];
assign int_rd_req_desc_b_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['hb];
assign int_rd_req_desc_b_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['hb];
assign int_rd_req_desc_b_axid_0_axid = int_rd_req_desc_n_axid_0_axid['hb];
assign int_rd_req_desc_b_axid_1_axid = int_rd_req_desc_n_axid_1_axid['hb];
assign int_rd_req_desc_b_axid_2_axid = int_rd_req_desc_n_axid_2_axid['hb];
assign int_rd_req_desc_b_axid_3_axid = int_rd_req_desc_n_axid_3_axid['hb];
assign int_rd_req_desc_b_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['hb];
assign int_rd_req_desc_b_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['hb];
assign int_rd_req_desc_b_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['hb];
assign int_rd_req_desc_b_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['hb];
assign int_rd_req_desc_b_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['hb];
assign int_rd_req_desc_b_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['hb];
assign int_rd_req_desc_b_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['hb];
assign int_rd_req_desc_b_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['hb];
assign int_rd_req_desc_b_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['hb];
assign int_rd_req_desc_b_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['hb];
assign int_rd_req_desc_b_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['hb];
assign int_rd_req_desc_b_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['hb];
assign int_rd_req_desc_b_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['hb];
assign int_rd_req_desc_b_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['hb];
assign int_rd_req_desc_b_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['hb];
assign int_rd_req_desc_b_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['hb];
assign int_wr_req_desc_b_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['hb];
assign int_wr_req_desc_b_size_txn_size = int_wr_req_desc_n_size_txn_size['hb];
assign int_wr_req_desc_b_data_offset_addr = int_wr_req_desc_n_data_offset_addr['hb];
assign int_wr_req_desc_b_axsize_axsize = int_wr_req_desc_n_axsize_axsize['hb];
assign int_wr_req_desc_b_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['hb];
assign int_wr_req_desc_b_attr_axdomain = int_wr_req_desc_n_attr_axdomain['hb];
assign int_wr_req_desc_b_attr_axbar = int_wr_req_desc_n_attr_axbar['hb];
assign int_wr_req_desc_b_attr_awunique = int_wr_req_desc_n_attr_awunique['hb];
assign int_wr_req_desc_b_attr_axregion = int_wr_req_desc_n_attr_axregion['hb];
assign int_wr_req_desc_b_attr_axqos = int_wr_req_desc_n_attr_axqos['hb];
assign int_wr_req_desc_b_attr_axprot = int_wr_req_desc_n_attr_axprot['hb];
assign int_wr_req_desc_b_attr_axcache = int_wr_req_desc_n_attr_axcache['hb];
assign int_wr_req_desc_b_attr_axlock = int_wr_req_desc_n_attr_axlock['hb];
assign int_wr_req_desc_b_attr_axburst = int_wr_req_desc_n_attr_axburst['hb];
assign int_wr_req_desc_b_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['hb];
assign int_wr_req_desc_b_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['hb];
assign int_wr_req_desc_b_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['hb];
assign int_wr_req_desc_b_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['hb];
assign int_wr_req_desc_b_axid_0_axid = int_wr_req_desc_n_axid_0_axid['hb];
assign int_wr_req_desc_b_axid_1_axid = int_wr_req_desc_n_axid_1_axid['hb];
assign int_wr_req_desc_b_axid_2_axid = int_wr_req_desc_n_axid_2_axid['hb];
assign int_wr_req_desc_b_axid_3_axid = int_wr_req_desc_n_axid_3_axid['hb];
assign int_wr_req_desc_b_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['hb];
assign int_wr_req_desc_b_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['hb];
assign int_wr_req_desc_b_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['hb];
assign int_wr_req_desc_b_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['hb];
assign int_wr_req_desc_b_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['hb];
assign int_wr_req_desc_b_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['hb];
assign int_wr_req_desc_b_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['hb];
assign int_wr_req_desc_b_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['hb];
assign int_wr_req_desc_b_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['hb];
assign int_wr_req_desc_b_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['hb];
assign int_wr_req_desc_b_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['hb];
assign int_wr_req_desc_b_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['hb];
assign int_wr_req_desc_b_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['hb];
assign int_wr_req_desc_b_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['hb];
assign int_wr_req_desc_b_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['hb];
assign int_wr_req_desc_b_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['hb];
assign int_wr_req_desc_b_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['hb];
assign int_wr_req_desc_b_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['hb];
assign int_wr_req_desc_b_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['hb];
assign int_wr_req_desc_b_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['hb];
assign int_wr_req_desc_b_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['hb];
assign int_wr_req_desc_b_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['hb];
assign int_wr_req_desc_b_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['hb];
assign int_wr_req_desc_b_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['hb];
assign int_wr_req_desc_b_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['hb];
assign int_wr_req_desc_b_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['hb];
assign int_wr_req_desc_b_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['hb];
assign int_wr_req_desc_b_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['hb];
assign int_wr_req_desc_b_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['hb];
assign int_wr_req_desc_b_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['hb];
assign int_wr_req_desc_b_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['hb];
assign int_wr_req_desc_b_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['hb];
assign int_sn_resp_desc_b_resp_resp = int_sn_resp_desc_n_resp_resp['hb];
assign int_rd_req_desc_c_size_txn_size = int_rd_req_desc_n_size_txn_size['hc];
assign int_rd_req_desc_c_axsize_axsize = int_rd_req_desc_n_axsize_axsize['hc];
assign int_rd_req_desc_c_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['hc];
assign int_rd_req_desc_c_attr_axdomain = int_rd_req_desc_n_attr_axdomain['hc];
assign int_rd_req_desc_c_attr_axbar = int_rd_req_desc_n_attr_axbar['hc];
assign int_rd_req_desc_c_attr_axregion = int_rd_req_desc_n_attr_axregion['hc];
assign int_rd_req_desc_c_attr_axqos = int_rd_req_desc_n_attr_axqos['hc];
assign int_rd_req_desc_c_attr_axprot = int_rd_req_desc_n_attr_axprot['hc];
assign int_rd_req_desc_c_attr_axcache = int_rd_req_desc_n_attr_axcache['hc];
assign int_rd_req_desc_c_attr_axlock = int_rd_req_desc_n_attr_axlock['hc];
assign int_rd_req_desc_c_attr_axburst = int_rd_req_desc_n_attr_axburst['hc];
assign int_rd_req_desc_c_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['hc];
assign int_rd_req_desc_c_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['hc];
assign int_rd_req_desc_c_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['hc];
assign int_rd_req_desc_c_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['hc];
assign int_rd_req_desc_c_axid_0_axid = int_rd_req_desc_n_axid_0_axid['hc];
assign int_rd_req_desc_c_axid_1_axid = int_rd_req_desc_n_axid_1_axid['hc];
assign int_rd_req_desc_c_axid_2_axid = int_rd_req_desc_n_axid_2_axid['hc];
assign int_rd_req_desc_c_axid_3_axid = int_rd_req_desc_n_axid_3_axid['hc];
assign int_rd_req_desc_c_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['hc];
assign int_rd_req_desc_c_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['hc];
assign int_rd_req_desc_c_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['hc];
assign int_rd_req_desc_c_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['hc];
assign int_rd_req_desc_c_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['hc];
assign int_rd_req_desc_c_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['hc];
assign int_rd_req_desc_c_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['hc];
assign int_rd_req_desc_c_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['hc];
assign int_rd_req_desc_c_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['hc];
assign int_rd_req_desc_c_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['hc];
assign int_rd_req_desc_c_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['hc];
assign int_rd_req_desc_c_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['hc];
assign int_rd_req_desc_c_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['hc];
assign int_rd_req_desc_c_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['hc];
assign int_rd_req_desc_c_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['hc];
assign int_rd_req_desc_c_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['hc];
assign int_wr_req_desc_c_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['hc];
assign int_wr_req_desc_c_size_txn_size = int_wr_req_desc_n_size_txn_size['hc];
assign int_wr_req_desc_c_data_offset_addr = int_wr_req_desc_n_data_offset_addr['hc];
assign int_wr_req_desc_c_axsize_axsize = int_wr_req_desc_n_axsize_axsize['hc];
assign int_wr_req_desc_c_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['hc];
assign int_wr_req_desc_c_attr_axdomain = int_wr_req_desc_n_attr_axdomain['hc];
assign int_wr_req_desc_c_attr_axbar = int_wr_req_desc_n_attr_axbar['hc];
assign int_wr_req_desc_c_attr_awunique = int_wr_req_desc_n_attr_awunique['hc];
assign int_wr_req_desc_c_attr_axregion = int_wr_req_desc_n_attr_axregion['hc];
assign int_wr_req_desc_c_attr_axqos = int_wr_req_desc_n_attr_axqos['hc];
assign int_wr_req_desc_c_attr_axprot = int_wr_req_desc_n_attr_axprot['hc];
assign int_wr_req_desc_c_attr_axcache = int_wr_req_desc_n_attr_axcache['hc];
assign int_wr_req_desc_c_attr_axlock = int_wr_req_desc_n_attr_axlock['hc];
assign int_wr_req_desc_c_attr_axburst = int_wr_req_desc_n_attr_axburst['hc];
assign int_wr_req_desc_c_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['hc];
assign int_wr_req_desc_c_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['hc];
assign int_wr_req_desc_c_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['hc];
assign int_wr_req_desc_c_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['hc];
assign int_wr_req_desc_c_axid_0_axid = int_wr_req_desc_n_axid_0_axid['hc];
assign int_wr_req_desc_c_axid_1_axid = int_wr_req_desc_n_axid_1_axid['hc];
assign int_wr_req_desc_c_axid_2_axid = int_wr_req_desc_n_axid_2_axid['hc];
assign int_wr_req_desc_c_axid_3_axid = int_wr_req_desc_n_axid_3_axid['hc];
assign int_wr_req_desc_c_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['hc];
assign int_wr_req_desc_c_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['hc];
assign int_wr_req_desc_c_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['hc];
assign int_wr_req_desc_c_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['hc];
assign int_wr_req_desc_c_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['hc];
assign int_wr_req_desc_c_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['hc];
assign int_wr_req_desc_c_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['hc];
assign int_wr_req_desc_c_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['hc];
assign int_wr_req_desc_c_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['hc];
assign int_wr_req_desc_c_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['hc];
assign int_wr_req_desc_c_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['hc];
assign int_wr_req_desc_c_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['hc];
assign int_wr_req_desc_c_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['hc];
assign int_wr_req_desc_c_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['hc];
assign int_wr_req_desc_c_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['hc];
assign int_wr_req_desc_c_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['hc];
assign int_wr_req_desc_c_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['hc];
assign int_wr_req_desc_c_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['hc];
assign int_wr_req_desc_c_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['hc];
assign int_wr_req_desc_c_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['hc];
assign int_wr_req_desc_c_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['hc];
assign int_wr_req_desc_c_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['hc];
assign int_wr_req_desc_c_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['hc];
assign int_wr_req_desc_c_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['hc];
assign int_wr_req_desc_c_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['hc];
assign int_wr_req_desc_c_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['hc];
assign int_wr_req_desc_c_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['hc];
assign int_wr_req_desc_c_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['hc];
assign int_wr_req_desc_c_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['hc];
assign int_wr_req_desc_c_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['hc];
assign int_wr_req_desc_c_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['hc];
assign int_wr_req_desc_c_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['hc];
assign int_sn_resp_desc_c_resp_resp = int_sn_resp_desc_n_resp_resp['hc];
assign int_rd_req_desc_d_size_txn_size = int_rd_req_desc_n_size_txn_size['hd];
assign int_rd_req_desc_d_axsize_axsize = int_rd_req_desc_n_axsize_axsize['hd];
assign int_rd_req_desc_d_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['hd];
assign int_rd_req_desc_d_attr_axdomain = int_rd_req_desc_n_attr_axdomain['hd];
assign int_rd_req_desc_d_attr_axbar = int_rd_req_desc_n_attr_axbar['hd];
assign int_rd_req_desc_d_attr_axregion = int_rd_req_desc_n_attr_axregion['hd];
assign int_rd_req_desc_d_attr_axqos = int_rd_req_desc_n_attr_axqos['hd];
assign int_rd_req_desc_d_attr_axprot = int_rd_req_desc_n_attr_axprot['hd];
assign int_rd_req_desc_d_attr_axcache = int_rd_req_desc_n_attr_axcache['hd];
assign int_rd_req_desc_d_attr_axlock = int_rd_req_desc_n_attr_axlock['hd];
assign int_rd_req_desc_d_attr_axburst = int_rd_req_desc_n_attr_axburst['hd];
assign int_rd_req_desc_d_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['hd];
assign int_rd_req_desc_d_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['hd];
assign int_rd_req_desc_d_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['hd];
assign int_rd_req_desc_d_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['hd];
assign int_rd_req_desc_d_axid_0_axid = int_rd_req_desc_n_axid_0_axid['hd];
assign int_rd_req_desc_d_axid_1_axid = int_rd_req_desc_n_axid_1_axid['hd];
assign int_rd_req_desc_d_axid_2_axid = int_rd_req_desc_n_axid_2_axid['hd];
assign int_rd_req_desc_d_axid_3_axid = int_rd_req_desc_n_axid_3_axid['hd];
assign int_rd_req_desc_d_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['hd];
assign int_rd_req_desc_d_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['hd];
assign int_rd_req_desc_d_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['hd];
assign int_rd_req_desc_d_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['hd];
assign int_rd_req_desc_d_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['hd];
assign int_rd_req_desc_d_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['hd];
assign int_rd_req_desc_d_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['hd];
assign int_rd_req_desc_d_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['hd];
assign int_rd_req_desc_d_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['hd];
assign int_rd_req_desc_d_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['hd];
assign int_rd_req_desc_d_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['hd];
assign int_rd_req_desc_d_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['hd];
assign int_rd_req_desc_d_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['hd];
assign int_rd_req_desc_d_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['hd];
assign int_rd_req_desc_d_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['hd];
assign int_rd_req_desc_d_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['hd];
assign int_wr_req_desc_d_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['hd];
assign int_wr_req_desc_d_size_txn_size = int_wr_req_desc_n_size_txn_size['hd];
assign int_wr_req_desc_d_data_offset_addr = int_wr_req_desc_n_data_offset_addr['hd];
assign int_wr_req_desc_d_axsize_axsize = int_wr_req_desc_n_axsize_axsize['hd];
assign int_wr_req_desc_d_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['hd];
assign int_wr_req_desc_d_attr_axdomain = int_wr_req_desc_n_attr_axdomain['hd];
assign int_wr_req_desc_d_attr_axbar = int_wr_req_desc_n_attr_axbar['hd];
assign int_wr_req_desc_d_attr_awunique = int_wr_req_desc_n_attr_awunique['hd];
assign int_wr_req_desc_d_attr_axregion = int_wr_req_desc_n_attr_axregion['hd];
assign int_wr_req_desc_d_attr_axqos = int_wr_req_desc_n_attr_axqos['hd];
assign int_wr_req_desc_d_attr_axprot = int_wr_req_desc_n_attr_axprot['hd];
assign int_wr_req_desc_d_attr_axcache = int_wr_req_desc_n_attr_axcache['hd];
assign int_wr_req_desc_d_attr_axlock = int_wr_req_desc_n_attr_axlock['hd];
assign int_wr_req_desc_d_attr_axburst = int_wr_req_desc_n_attr_axburst['hd];
assign int_wr_req_desc_d_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['hd];
assign int_wr_req_desc_d_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['hd];
assign int_wr_req_desc_d_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['hd];
assign int_wr_req_desc_d_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['hd];
assign int_wr_req_desc_d_axid_0_axid = int_wr_req_desc_n_axid_0_axid['hd];
assign int_wr_req_desc_d_axid_1_axid = int_wr_req_desc_n_axid_1_axid['hd];
assign int_wr_req_desc_d_axid_2_axid = int_wr_req_desc_n_axid_2_axid['hd];
assign int_wr_req_desc_d_axid_3_axid = int_wr_req_desc_n_axid_3_axid['hd];
assign int_wr_req_desc_d_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['hd];
assign int_wr_req_desc_d_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['hd];
assign int_wr_req_desc_d_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['hd];
assign int_wr_req_desc_d_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['hd];
assign int_wr_req_desc_d_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['hd];
assign int_wr_req_desc_d_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['hd];
assign int_wr_req_desc_d_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['hd];
assign int_wr_req_desc_d_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['hd];
assign int_wr_req_desc_d_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['hd];
assign int_wr_req_desc_d_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['hd];
assign int_wr_req_desc_d_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['hd];
assign int_wr_req_desc_d_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['hd];
assign int_wr_req_desc_d_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['hd];
assign int_wr_req_desc_d_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['hd];
assign int_wr_req_desc_d_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['hd];
assign int_wr_req_desc_d_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['hd];
assign int_wr_req_desc_d_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['hd];
assign int_wr_req_desc_d_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['hd];
assign int_wr_req_desc_d_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['hd];
assign int_wr_req_desc_d_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['hd];
assign int_wr_req_desc_d_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['hd];
assign int_wr_req_desc_d_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['hd];
assign int_wr_req_desc_d_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['hd];
assign int_wr_req_desc_d_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['hd];
assign int_wr_req_desc_d_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['hd];
assign int_wr_req_desc_d_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['hd];
assign int_wr_req_desc_d_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['hd];
assign int_wr_req_desc_d_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['hd];
assign int_wr_req_desc_d_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['hd];
assign int_wr_req_desc_d_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['hd];
assign int_wr_req_desc_d_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['hd];
assign int_wr_req_desc_d_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['hd];
assign int_sn_resp_desc_d_resp_resp = int_sn_resp_desc_n_resp_resp['hd];
assign int_rd_req_desc_e_size_txn_size = int_rd_req_desc_n_size_txn_size['he];
assign int_rd_req_desc_e_axsize_axsize = int_rd_req_desc_n_axsize_axsize['he];
assign int_rd_req_desc_e_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['he];
assign int_rd_req_desc_e_attr_axdomain = int_rd_req_desc_n_attr_axdomain['he];
assign int_rd_req_desc_e_attr_axbar = int_rd_req_desc_n_attr_axbar['he];
assign int_rd_req_desc_e_attr_axregion = int_rd_req_desc_n_attr_axregion['he];
assign int_rd_req_desc_e_attr_axqos = int_rd_req_desc_n_attr_axqos['he];
assign int_rd_req_desc_e_attr_axprot = int_rd_req_desc_n_attr_axprot['he];
assign int_rd_req_desc_e_attr_axcache = int_rd_req_desc_n_attr_axcache['he];
assign int_rd_req_desc_e_attr_axlock = int_rd_req_desc_n_attr_axlock['he];
assign int_rd_req_desc_e_attr_axburst = int_rd_req_desc_n_attr_axburst['he];
assign int_rd_req_desc_e_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['he];
assign int_rd_req_desc_e_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['he];
assign int_rd_req_desc_e_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['he];
assign int_rd_req_desc_e_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['he];
assign int_rd_req_desc_e_axid_0_axid = int_rd_req_desc_n_axid_0_axid['he];
assign int_rd_req_desc_e_axid_1_axid = int_rd_req_desc_n_axid_1_axid['he];
assign int_rd_req_desc_e_axid_2_axid = int_rd_req_desc_n_axid_2_axid['he];
assign int_rd_req_desc_e_axid_3_axid = int_rd_req_desc_n_axid_3_axid['he];
assign int_rd_req_desc_e_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['he];
assign int_rd_req_desc_e_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['he];
assign int_rd_req_desc_e_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['he];
assign int_rd_req_desc_e_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['he];
assign int_rd_req_desc_e_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['he];
assign int_rd_req_desc_e_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['he];
assign int_rd_req_desc_e_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['he];
assign int_rd_req_desc_e_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['he];
assign int_rd_req_desc_e_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['he];
assign int_rd_req_desc_e_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['he];
assign int_rd_req_desc_e_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['he];
assign int_rd_req_desc_e_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['he];
assign int_rd_req_desc_e_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['he];
assign int_rd_req_desc_e_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['he];
assign int_rd_req_desc_e_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['he];
assign int_rd_req_desc_e_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['he];
assign int_wr_req_desc_e_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['he];
assign int_wr_req_desc_e_size_txn_size = int_wr_req_desc_n_size_txn_size['he];
assign int_wr_req_desc_e_data_offset_addr = int_wr_req_desc_n_data_offset_addr['he];
assign int_wr_req_desc_e_axsize_axsize = int_wr_req_desc_n_axsize_axsize['he];
assign int_wr_req_desc_e_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['he];
assign int_wr_req_desc_e_attr_axdomain = int_wr_req_desc_n_attr_axdomain['he];
assign int_wr_req_desc_e_attr_axbar = int_wr_req_desc_n_attr_axbar['he];
assign int_wr_req_desc_e_attr_awunique = int_wr_req_desc_n_attr_awunique['he];
assign int_wr_req_desc_e_attr_axregion = int_wr_req_desc_n_attr_axregion['he];
assign int_wr_req_desc_e_attr_axqos = int_wr_req_desc_n_attr_axqos['he];
assign int_wr_req_desc_e_attr_axprot = int_wr_req_desc_n_attr_axprot['he];
assign int_wr_req_desc_e_attr_axcache = int_wr_req_desc_n_attr_axcache['he];
assign int_wr_req_desc_e_attr_axlock = int_wr_req_desc_n_attr_axlock['he];
assign int_wr_req_desc_e_attr_axburst = int_wr_req_desc_n_attr_axburst['he];
assign int_wr_req_desc_e_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['he];
assign int_wr_req_desc_e_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['he];
assign int_wr_req_desc_e_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['he];
assign int_wr_req_desc_e_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['he];
assign int_wr_req_desc_e_axid_0_axid = int_wr_req_desc_n_axid_0_axid['he];
assign int_wr_req_desc_e_axid_1_axid = int_wr_req_desc_n_axid_1_axid['he];
assign int_wr_req_desc_e_axid_2_axid = int_wr_req_desc_n_axid_2_axid['he];
assign int_wr_req_desc_e_axid_3_axid = int_wr_req_desc_n_axid_3_axid['he];
assign int_wr_req_desc_e_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['he];
assign int_wr_req_desc_e_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['he];
assign int_wr_req_desc_e_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['he];
assign int_wr_req_desc_e_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['he];
assign int_wr_req_desc_e_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['he];
assign int_wr_req_desc_e_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['he];
assign int_wr_req_desc_e_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['he];
assign int_wr_req_desc_e_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['he];
assign int_wr_req_desc_e_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['he];
assign int_wr_req_desc_e_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['he];
assign int_wr_req_desc_e_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['he];
assign int_wr_req_desc_e_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['he];
assign int_wr_req_desc_e_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['he];
assign int_wr_req_desc_e_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['he];
assign int_wr_req_desc_e_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['he];
assign int_wr_req_desc_e_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['he];
assign int_wr_req_desc_e_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['he];
assign int_wr_req_desc_e_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['he];
assign int_wr_req_desc_e_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['he];
assign int_wr_req_desc_e_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['he];
assign int_wr_req_desc_e_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['he];
assign int_wr_req_desc_e_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['he];
assign int_wr_req_desc_e_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['he];
assign int_wr_req_desc_e_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['he];
assign int_wr_req_desc_e_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['he];
assign int_wr_req_desc_e_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['he];
assign int_wr_req_desc_e_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['he];
assign int_wr_req_desc_e_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['he];
assign int_wr_req_desc_e_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['he];
assign int_wr_req_desc_e_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['he];
assign int_wr_req_desc_e_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['he];
assign int_wr_req_desc_e_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['he];
assign int_sn_resp_desc_e_resp_resp = int_sn_resp_desc_n_resp_resp['he];
assign int_rd_req_desc_f_size_txn_size = int_rd_req_desc_n_size_txn_size['hf];
assign int_rd_req_desc_f_axsize_axsize = int_rd_req_desc_n_axsize_axsize['hf];
assign int_rd_req_desc_f_attr_axsnoop = int_rd_req_desc_n_attr_axsnoop['hf];
assign int_rd_req_desc_f_attr_axdomain = int_rd_req_desc_n_attr_axdomain['hf];
assign int_rd_req_desc_f_attr_axbar = int_rd_req_desc_n_attr_axbar['hf];
assign int_rd_req_desc_f_attr_axregion = int_rd_req_desc_n_attr_axregion['hf];
assign int_rd_req_desc_f_attr_axqos = int_rd_req_desc_n_attr_axqos['hf];
assign int_rd_req_desc_f_attr_axprot = int_rd_req_desc_n_attr_axprot['hf];
assign int_rd_req_desc_f_attr_axcache = int_rd_req_desc_n_attr_axcache['hf];
assign int_rd_req_desc_f_attr_axlock = int_rd_req_desc_n_attr_axlock['hf];
assign int_rd_req_desc_f_attr_axburst = int_rd_req_desc_n_attr_axburst['hf];
assign int_rd_req_desc_f_axaddr_0_addr = int_rd_req_desc_n_axaddr_0_addr['hf];
assign int_rd_req_desc_f_axaddr_1_addr = int_rd_req_desc_n_axaddr_1_addr['hf];
assign int_rd_req_desc_f_axaddr_2_addr = int_rd_req_desc_n_axaddr_2_addr['hf];
assign int_rd_req_desc_f_axaddr_3_addr = int_rd_req_desc_n_axaddr_3_addr['hf];
assign int_rd_req_desc_f_axid_0_axid = int_rd_req_desc_n_axid_0_axid['hf];
assign int_rd_req_desc_f_axid_1_axid = int_rd_req_desc_n_axid_1_axid['hf];
assign int_rd_req_desc_f_axid_2_axid = int_rd_req_desc_n_axid_2_axid['hf];
assign int_rd_req_desc_f_axid_3_axid = int_rd_req_desc_n_axid_3_axid['hf];
assign int_rd_req_desc_f_axuser_0_axuser = int_rd_req_desc_n_axuser_0_axuser['hf];
assign int_rd_req_desc_f_axuser_1_axuser = int_rd_req_desc_n_axuser_1_axuser['hf];
assign int_rd_req_desc_f_axuser_2_axuser = int_rd_req_desc_n_axuser_2_axuser['hf];
assign int_rd_req_desc_f_axuser_3_axuser = int_rd_req_desc_n_axuser_3_axuser['hf];
assign int_rd_req_desc_f_axuser_4_axuser = int_rd_req_desc_n_axuser_4_axuser['hf];
assign int_rd_req_desc_f_axuser_5_axuser = int_rd_req_desc_n_axuser_5_axuser['hf];
assign int_rd_req_desc_f_axuser_6_axuser = int_rd_req_desc_n_axuser_6_axuser['hf];
assign int_rd_req_desc_f_axuser_7_axuser = int_rd_req_desc_n_axuser_7_axuser['hf];
assign int_rd_req_desc_f_axuser_8_axuser = int_rd_req_desc_n_axuser_8_axuser['hf];
assign int_rd_req_desc_f_axuser_9_axuser = int_rd_req_desc_n_axuser_9_axuser['hf];
assign int_rd_req_desc_f_axuser_10_axuser = int_rd_req_desc_n_axuser_10_axuser['hf];
assign int_rd_req_desc_f_axuser_11_axuser = int_rd_req_desc_n_axuser_11_axuser['hf];
assign int_rd_req_desc_f_axuser_12_axuser = int_rd_req_desc_n_axuser_12_axuser['hf];
assign int_rd_req_desc_f_axuser_13_axuser = int_rd_req_desc_n_axuser_13_axuser['hf];
assign int_rd_req_desc_f_axuser_14_axuser = int_rd_req_desc_n_axuser_14_axuser['hf];
assign int_rd_req_desc_f_axuser_15_axuser = int_rd_req_desc_n_axuser_15_axuser['hf];
assign int_wr_req_desc_f_txn_type_wr_strb = int_wr_req_desc_n_txn_type_wr_strb['hf];
assign int_wr_req_desc_f_size_txn_size = int_wr_req_desc_n_size_txn_size['hf];
assign int_wr_req_desc_f_data_offset_addr = int_wr_req_desc_n_data_offset_addr['hf];
assign int_wr_req_desc_f_axsize_axsize = int_wr_req_desc_n_axsize_axsize['hf];
assign int_wr_req_desc_f_attr_axsnoop = int_wr_req_desc_n_attr_axsnoop['hf];
assign int_wr_req_desc_f_attr_axdomain = int_wr_req_desc_n_attr_axdomain['hf];
assign int_wr_req_desc_f_attr_axbar = int_wr_req_desc_n_attr_axbar['hf];
assign int_wr_req_desc_f_attr_awunique = int_wr_req_desc_n_attr_awunique['hf];
assign int_wr_req_desc_f_attr_axregion = int_wr_req_desc_n_attr_axregion['hf];
assign int_wr_req_desc_f_attr_axqos = int_wr_req_desc_n_attr_axqos['hf];
assign int_wr_req_desc_f_attr_axprot = int_wr_req_desc_n_attr_axprot['hf];
assign int_wr_req_desc_f_attr_axcache = int_wr_req_desc_n_attr_axcache['hf];
assign int_wr_req_desc_f_attr_axlock = int_wr_req_desc_n_attr_axlock['hf];
assign int_wr_req_desc_f_attr_axburst = int_wr_req_desc_n_attr_axburst['hf];
assign int_wr_req_desc_f_axaddr_0_addr = int_wr_req_desc_n_axaddr_0_addr['hf];
assign int_wr_req_desc_f_axaddr_1_addr = int_wr_req_desc_n_axaddr_1_addr['hf];
assign int_wr_req_desc_f_axaddr_2_addr = int_wr_req_desc_n_axaddr_2_addr['hf];
assign int_wr_req_desc_f_axaddr_3_addr = int_wr_req_desc_n_axaddr_3_addr['hf];
assign int_wr_req_desc_f_axid_0_axid = int_wr_req_desc_n_axid_0_axid['hf];
assign int_wr_req_desc_f_axid_1_axid = int_wr_req_desc_n_axid_1_axid['hf];
assign int_wr_req_desc_f_axid_2_axid = int_wr_req_desc_n_axid_2_axid['hf];
assign int_wr_req_desc_f_axid_3_axid = int_wr_req_desc_n_axid_3_axid['hf];
assign int_wr_req_desc_f_axuser_0_axuser = int_wr_req_desc_n_axuser_0_axuser['hf];
assign int_wr_req_desc_f_axuser_1_axuser = int_wr_req_desc_n_axuser_1_axuser['hf];
assign int_wr_req_desc_f_axuser_2_axuser = int_wr_req_desc_n_axuser_2_axuser['hf];
assign int_wr_req_desc_f_axuser_3_axuser = int_wr_req_desc_n_axuser_3_axuser['hf];
assign int_wr_req_desc_f_axuser_4_axuser = int_wr_req_desc_n_axuser_4_axuser['hf];
assign int_wr_req_desc_f_axuser_5_axuser = int_wr_req_desc_n_axuser_5_axuser['hf];
assign int_wr_req_desc_f_axuser_6_axuser = int_wr_req_desc_n_axuser_6_axuser['hf];
assign int_wr_req_desc_f_axuser_7_axuser = int_wr_req_desc_n_axuser_7_axuser['hf];
assign int_wr_req_desc_f_axuser_8_axuser = int_wr_req_desc_n_axuser_8_axuser['hf];
assign int_wr_req_desc_f_axuser_9_axuser = int_wr_req_desc_n_axuser_9_axuser['hf];
assign int_wr_req_desc_f_axuser_10_axuser = int_wr_req_desc_n_axuser_10_axuser['hf];
assign int_wr_req_desc_f_axuser_11_axuser = int_wr_req_desc_n_axuser_11_axuser['hf];
assign int_wr_req_desc_f_axuser_12_axuser = int_wr_req_desc_n_axuser_12_axuser['hf];
assign int_wr_req_desc_f_axuser_13_axuser = int_wr_req_desc_n_axuser_13_axuser['hf];
assign int_wr_req_desc_f_axuser_14_axuser = int_wr_req_desc_n_axuser_14_axuser['hf];
assign int_wr_req_desc_f_axuser_15_axuser = int_wr_req_desc_n_axuser_15_axuser['hf];
assign int_wr_req_desc_f_wuser_0_wuser = int_wr_req_desc_n_wuser_0_wuser['hf];
assign int_wr_req_desc_f_wuser_1_wuser = int_wr_req_desc_n_wuser_1_wuser['hf];
assign int_wr_req_desc_f_wuser_2_wuser = int_wr_req_desc_n_wuser_2_wuser['hf];
assign int_wr_req_desc_f_wuser_3_wuser = int_wr_req_desc_n_wuser_3_wuser['hf];
assign int_wr_req_desc_f_wuser_4_wuser = int_wr_req_desc_n_wuser_4_wuser['hf];
assign int_wr_req_desc_f_wuser_5_wuser = int_wr_req_desc_n_wuser_5_wuser['hf];
assign int_wr_req_desc_f_wuser_6_wuser = int_wr_req_desc_n_wuser_6_wuser['hf];
assign int_wr_req_desc_f_wuser_7_wuser = int_wr_req_desc_n_wuser_7_wuser['hf];
assign int_wr_req_desc_f_wuser_8_wuser = int_wr_req_desc_n_wuser_8_wuser['hf];
assign int_wr_req_desc_f_wuser_9_wuser = int_wr_req_desc_n_wuser_9_wuser['hf];
assign int_wr_req_desc_f_wuser_10_wuser = int_wr_req_desc_n_wuser_10_wuser['hf];
assign int_wr_req_desc_f_wuser_11_wuser = int_wr_req_desc_n_wuser_11_wuser['hf];
assign int_wr_req_desc_f_wuser_12_wuser = int_wr_req_desc_n_wuser_12_wuser['hf];
assign int_wr_req_desc_f_wuser_13_wuser = int_wr_req_desc_n_wuser_13_wuser['hf];
assign int_wr_req_desc_f_wuser_14_wuser = int_wr_req_desc_n_wuser_14_wuser['hf];
assign int_wr_req_desc_f_wuser_15_wuser = int_wr_req_desc_n_wuser_15_wuser['hf];
assign int_sn_resp_desc_f_resp_resp = int_sn_resp_desc_n_resp_resp['hf];
assign int_rd_resp_desc_n_data_offset_addr['h0] = int_rd_resp_desc_0_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h0] = int_rd_resp_desc_0_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h0] = int_rd_resp_desc_0_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h0] = int_rd_resp_desc_0_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h0] = int_rd_resp_desc_0_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h0] = int_rd_resp_desc_0_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h0] = int_rd_resp_desc_0_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h0] = int_rd_resp_desc_0_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h0] = int_rd_resp_desc_0_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h0] = int_rd_resp_desc_0_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h0] = int_rd_resp_desc_0_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h0] = int_rd_resp_desc_0_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h0] = int_rd_resp_desc_0_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h0] = int_rd_resp_desc_0_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h0] = int_rd_resp_desc_0_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h0] = int_rd_resp_desc_0_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h0] = int_rd_resp_desc_0_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h0] = int_rd_resp_desc_0_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h0] = int_rd_resp_desc_0_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h0] = int_rd_resp_desc_0_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h0] = int_rd_resp_desc_0_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h0] = int_rd_resp_desc_0_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h0] = int_rd_resp_desc_0_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h0] = int_rd_resp_desc_0_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h0] = int_rd_resp_desc_0_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h0] = int_rd_resp_desc_0_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h0] = int_rd_resp_desc_0_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h0] = int_wr_req_desc_0_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h0] = int_wr_req_desc_0_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h0] = int_wr_req_desc_0_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h0] = int_wr_req_desc_0_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h0] = int_wr_req_desc_0_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h0] = int_wr_req_desc_0_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h0] = int_wr_req_desc_0_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h0] = int_wr_req_desc_0_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h0] = int_wr_resp_desc_0_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h0] = int_wr_resp_desc_0_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h0] = int_wr_resp_desc_0_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h0] = int_wr_resp_desc_0_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h0] = int_wr_resp_desc_0_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h0] = int_wr_resp_desc_0_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h0] = int_wr_resp_desc_0_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h0] = int_wr_resp_desc_0_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h0] = int_wr_resp_desc_0_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h0] = int_wr_resp_desc_0_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h0] = int_wr_resp_desc_0_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h0] = int_wr_resp_desc_0_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h0] = int_wr_resp_desc_0_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h0] = int_wr_resp_desc_0_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h0] = int_wr_resp_desc_0_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h0] = int_wr_resp_desc_0_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h0] = int_wr_resp_desc_0_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h0] = int_wr_resp_desc_0_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h0] = int_wr_resp_desc_0_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h0] = int_wr_resp_desc_0_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h0] = int_wr_resp_desc_0_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h0] = int_sn_req_desc_0_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h0] = int_sn_req_desc_0_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h0] = int_sn_req_desc_0_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h0] = int_sn_req_desc_0_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h0] = int_sn_req_desc_0_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h0] = int_sn_req_desc_0_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h1] = int_rd_resp_desc_1_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h1] = int_rd_resp_desc_1_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h1] = int_rd_resp_desc_1_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h1] = int_rd_resp_desc_1_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h1] = int_rd_resp_desc_1_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h1] = int_rd_resp_desc_1_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h1] = int_rd_resp_desc_1_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h1] = int_rd_resp_desc_1_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h1] = int_rd_resp_desc_1_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h1] = int_rd_resp_desc_1_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h1] = int_rd_resp_desc_1_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h1] = int_rd_resp_desc_1_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h1] = int_rd_resp_desc_1_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h1] = int_rd_resp_desc_1_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h1] = int_rd_resp_desc_1_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h1] = int_rd_resp_desc_1_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h1] = int_rd_resp_desc_1_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h1] = int_rd_resp_desc_1_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h1] = int_rd_resp_desc_1_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h1] = int_rd_resp_desc_1_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h1] = int_rd_resp_desc_1_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h1] = int_rd_resp_desc_1_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h1] = int_rd_resp_desc_1_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h1] = int_rd_resp_desc_1_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h1] = int_rd_resp_desc_1_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h1] = int_rd_resp_desc_1_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h1] = int_rd_resp_desc_1_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h1] = int_wr_req_desc_1_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h1] = int_wr_req_desc_1_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h1] = int_wr_req_desc_1_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h1] = int_wr_req_desc_1_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h1] = int_wr_req_desc_1_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h1] = int_wr_req_desc_1_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h1] = int_wr_req_desc_1_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h1] = int_wr_req_desc_1_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h1] = int_wr_resp_desc_1_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h1] = int_wr_resp_desc_1_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h1] = int_wr_resp_desc_1_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h1] = int_wr_resp_desc_1_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h1] = int_wr_resp_desc_1_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h1] = int_wr_resp_desc_1_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h1] = int_wr_resp_desc_1_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h1] = int_wr_resp_desc_1_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h1] = int_wr_resp_desc_1_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h1] = int_wr_resp_desc_1_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h1] = int_wr_resp_desc_1_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h1] = int_wr_resp_desc_1_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h1] = int_wr_resp_desc_1_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h1] = int_wr_resp_desc_1_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h1] = int_wr_resp_desc_1_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h1] = int_wr_resp_desc_1_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h1] = int_wr_resp_desc_1_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h1] = int_wr_resp_desc_1_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h1] = int_wr_resp_desc_1_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h1] = int_wr_resp_desc_1_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h1] = int_wr_resp_desc_1_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h1] = int_sn_req_desc_1_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h1] = int_sn_req_desc_1_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h1] = int_sn_req_desc_1_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h1] = int_sn_req_desc_1_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h1] = int_sn_req_desc_1_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h1] = int_sn_req_desc_1_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h2] = int_rd_resp_desc_2_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h2] = int_rd_resp_desc_2_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h2] = int_rd_resp_desc_2_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h2] = int_rd_resp_desc_2_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h2] = int_rd_resp_desc_2_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h2] = int_rd_resp_desc_2_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h2] = int_rd_resp_desc_2_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h2] = int_rd_resp_desc_2_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h2] = int_rd_resp_desc_2_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h2] = int_rd_resp_desc_2_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h2] = int_rd_resp_desc_2_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h2] = int_rd_resp_desc_2_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h2] = int_rd_resp_desc_2_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h2] = int_rd_resp_desc_2_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h2] = int_rd_resp_desc_2_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h2] = int_rd_resp_desc_2_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h2] = int_rd_resp_desc_2_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h2] = int_rd_resp_desc_2_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h2] = int_rd_resp_desc_2_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h2] = int_rd_resp_desc_2_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h2] = int_rd_resp_desc_2_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h2] = int_rd_resp_desc_2_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h2] = int_rd_resp_desc_2_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h2] = int_rd_resp_desc_2_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h2] = int_rd_resp_desc_2_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h2] = int_rd_resp_desc_2_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h2] = int_rd_resp_desc_2_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h2] = int_wr_req_desc_2_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h2] = int_wr_req_desc_2_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h2] = int_wr_req_desc_2_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h2] = int_wr_req_desc_2_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h2] = int_wr_req_desc_2_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h2] = int_wr_req_desc_2_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h2] = int_wr_req_desc_2_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h2] = int_wr_req_desc_2_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h2] = int_wr_resp_desc_2_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h2] = int_wr_resp_desc_2_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h2] = int_wr_resp_desc_2_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h2] = int_wr_resp_desc_2_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h2] = int_wr_resp_desc_2_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h2] = int_wr_resp_desc_2_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h2] = int_wr_resp_desc_2_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h2] = int_wr_resp_desc_2_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h2] = int_wr_resp_desc_2_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h2] = int_wr_resp_desc_2_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h2] = int_wr_resp_desc_2_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h2] = int_wr_resp_desc_2_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h2] = int_wr_resp_desc_2_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h2] = int_wr_resp_desc_2_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h2] = int_wr_resp_desc_2_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h2] = int_wr_resp_desc_2_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h2] = int_wr_resp_desc_2_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h2] = int_wr_resp_desc_2_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h2] = int_wr_resp_desc_2_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h2] = int_wr_resp_desc_2_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h2] = int_wr_resp_desc_2_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h2] = int_sn_req_desc_2_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h2] = int_sn_req_desc_2_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h2] = int_sn_req_desc_2_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h2] = int_sn_req_desc_2_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h2] = int_sn_req_desc_2_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h2] = int_sn_req_desc_2_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h3] = int_rd_resp_desc_3_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h3] = int_rd_resp_desc_3_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h3] = int_rd_resp_desc_3_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h3] = int_rd_resp_desc_3_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h3] = int_rd_resp_desc_3_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h3] = int_rd_resp_desc_3_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h3] = int_rd_resp_desc_3_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h3] = int_rd_resp_desc_3_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h3] = int_rd_resp_desc_3_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h3] = int_rd_resp_desc_3_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h3] = int_rd_resp_desc_3_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h3] = int_rd_resp_desc_3_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h3] = int_rd_resp_desc_3_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h3] = int_rd_resp_desc_3_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h3] = int_rd_resp_desc_3_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h3] = int_rd_resp_desc_3_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h3] = int_rd_resp_desc_3_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h3] = int_rd_resp_desc_3_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h3] = int_rd_resp_desc_3_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h3] = int_rd_resp_desc_3_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h3] = int_rd_resp_desc_3_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h3] = int_rd_resp_desc_3_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h3] = int_rd_resp_desc_3_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h3] = int_rd_resp_desc_3_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h3] = int_rd_resp_desc_3_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h3] = int_rd_resp_desc_3_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h3] = int_rd_resp_desc_3_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h3] = int_wr_req_desc_3_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h3] = int_wr_req_desc_3_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h3] = int_wr_req_desc_3_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h3] = int_wr_req_desc_3_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h3] = int_wr_req_desc_3_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h3] = int_wr_req_desc_3_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h3] = int_wr_req_desc_3_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h3] = int_wr_req_desc_3_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h3] = int_wr_resp_desc_3_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h3] = int_wr_resp_desc_3_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h3] = int_wr_resp_desc_3_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h3] = int_wr_resp_desc_3_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h3] = int_wr_resp_desc_3_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h3] = int_wr_resp_desc_3_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h3] = int_wr_resp_desc_3_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h3] = int_wr_resp_desc_3_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h3] = int_wr_resp_desc_3_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h3] = int_wr_resp_desc_3_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h3] = int_wr_resp_desc_3_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h3] = int_wr_resp_desc_3_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h3] = int_wr_resp_desc_3_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h3] = int_wr_resp_desc_3_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h3] = int_wr_resp_desc_3_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h3] = int_wr_resp_desc_3_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h3] = int_wr_resp_desc_3_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h3] = int_wr_resp_desc_3_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h3] = int_wr_resp_desc_3_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h3] = int_wr_resp_desc_3_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h3] = int_wr_resp_desc_3_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h3] = int_sn_req_desc_3_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h3] = int_sn_req_desc_3_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h3] = int_sn_req_desc_3_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h3] = int_sn_req_desc_3_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h3] = int_sn_req_desc_3_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h3] = int_sn_req_desc_3_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h4] = int_rd_resp_desc_4_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h4] = int_rd_resp_desc_4_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h4] = int_rd_resp_desc_4_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h4] = int_rd_resp_desc_4_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h4] = int_rd_resp_desc_4_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h4] = int_rd_resp_desc_4_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h4] = int_rd_resp_desc_4_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h4] = int_rd_resp_desc_4_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h4] = int_rd_resp_desc_4_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h4] = int_rd_resp_desc_4_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h4] = int_rd_resp_desc_4_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h4] = int_rd_resp_desc_4_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h4] = int_rd_resp_desc_4_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h4] = int_rd_resp_desc_4_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h4] = int_rd_resp_desc_4_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h4] = int_rd_resp_desc_4_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h4] = int_rd_resp_desc_4_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h4] = int_rd_resp_desc_4_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h4] = int_rd_resp_desc_4_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h4] = int_rd_resp_desc_4_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h4] = int_rd_resp_desc_4_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h4] = int_rd_resp_desc_4_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h4] = int_rd_resp_desc_4_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h4] = int_rd_resp_desc_4_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h4] = int_rd_resp_desc_4_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h4] = int_rd_resp_desc_4_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h4] = int_rd_resp_desc_4_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h4] = int_wr_req_desc_4_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h4] = int_wr_req_desc_4_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h4] = int_wr_req_desc_4_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h4] = int_wr_req_desc_4_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h4] = int_wr_req_desc_4_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h4] = int_wr_req_desc_4_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h4] = int_wr_req_desc_4_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h4] = int_wr_req_desc_4_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h4] = int_wr_resp_desc_4_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h4] = int_wr_resp_desc_4_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h4] = int_wr_resp_desc_4_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h4] = int_wr_resp_desc_4_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h4] = int_wr_resp_desc_4_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h4] = int_wr_resp_desc_4_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h4] = int_wr_resp_desc_4_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h4] = int_wr_resp_desc_4_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h4] = int_wr_resp_desc_4_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h4] = int_wr_resp_desc_4_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h4] = int_wr_resp_desc_4_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h4] = int_wr_resp_desc_4_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h4] = int_wr_resp_desc_4_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h4] = int_wr_resp_desc_4_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h4] = int_wr_resp_desc_4_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h4] = int_wr_resp_desc_4_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h4] = int_wr_resp_desc_4_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h4] = int_wr_resp_desc_4_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h4] = int_wr_resp_desc_4_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h4] = int_wr_resp_desc_4_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h4] = int_wr_resp_desc_4_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h4] = int_sn_req_desc_4_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h4] = int_sn_req_desc_4_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h4] = int_sn_req_desc_4_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h4] = int_sn_req_desc_4_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h4] = int_sn_req_desc_4_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h4] = int_sn_req_desc_4_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h5] = int_rd_resp_desc_5_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h5] = int_rd_resp_desc_5_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h5] = int_rd_resp_desc_5_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h5] = int_rd_resp_desc_5_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h5] = int_rd_resp_desc_5_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h5] = int_rd_resp_desc_5_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h5] = int_rd_resp_desc_5_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h5] = int_rd_resp_desc_5_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h5] = int_rd_resp_desc_5_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h5] = int_rd_resp_desc_5_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h5] = int_rd_resp_desc_5_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h5] = int_rd_resp_desc_5_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h5] = int_rd_resp_desc_5_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h5] = int_rd_resp_desc_5_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h5] = int_rd_resp_desc_5_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h5] = int_rd_resp_desc_5_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h5] = int_rd_resp_desc_5_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h5] = int_rd_resp_desc_5_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h5] = int_rd_resp_desc_5_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h5] = int_rd_resp_desc_5_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h5] = int_rd_resp_desc_5_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h5] = int_rd_resp_desc_5_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h5] = int_rd_resp_desc_5_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h5] = int_rd_resp_desc_5_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h5] = int_rd_resp_desc_5_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h5] = int_rd_resp_desc_5_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h5] = int_rd_resp_desc_5_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h5] = int_wr_req_desc_5_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h5] = int_wr_req_desc_5_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h5] = int_wr_req_desc_5_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h5] = int_wr_req_desc_5_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h5] = int_wr_req_desc_5_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h5] = int_wr_req_desc_5_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h5] = int_wr_req_desc_5_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h5] = int_wr_req_desc_5_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h5] = int_wr_resp_desc_5_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h5] = int_wr_resp_desc_5_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h5] = int_wr_resp_desc_5_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h5] = int_wr_resp_desc_5_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h5] = int_wr_resp_desc_5_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h5] = int_wr_resp_desc_5_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h5] = int_wr_resp_desc_5_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h5] = int_wr_resp_desc_5_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h5] = int_wr_resp_desc_5_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h5] = int_wr_resp_desc_5_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h5] = int_wr_resp_desc_5_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h5] = int_wr_resp_desc_5_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h5] = int_wr_resp_desc_5_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h5] = int_wr_resp_desc_5_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h5] = int_wr_resp_desc_5_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h5] = int_wr_resp_desc_5_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h5] = int_wr_resp_desc_5_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h5] = int_wr_resp_desc_5_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h5] = int_wr_resp_desc_5_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h5] = int_wr_resp_desc_5_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h5] = int_wr_resp_desc_5_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h5] = int_sn_req_desc_5_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h5] = int_sn_req_desc_5_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h5] = int_sn_req_desc_5_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h5] = int_sn_req_desc_5_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h5] = int_sn_req_desc_5_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h5] = int_sn_req_desc_5_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h6] = int_rd_resp_desc_6_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h6] = int_rd_resp_desc_6_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h6] = int_rd_resp_desc_6_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h6] = int_rd_resp_desc_6_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h6] = int_rd_resp_desc_6_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h6] = int_rd_resp_desc_6_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h6] = int_rd_resp_desc_6_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h6] = int_rd_resp_desc_6_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h6] = int_rd_resp_desc_6_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h6] = int_rd_resp_desc_6_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h6] = int_rd_resp_desc_6_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h6] = int_rd_resp_desc_6_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h6] = int_rd_resp_desc_6_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h6] = int_rd_resp_desc_6_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h6] = int_rd_resp_desc_6_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h6] = int_rd_resp_desc_6_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h6] = int_rd_resp_desc_6_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h6] = int_rd_resp_desc_6_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h6] = int_rd_resp_desc_6_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h6] = int_rd_resp_desc_6_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h6] = int_rd_resp_desc_6_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h6] = int_rd_resp_desc_6_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h6] = int_rd_resp_desc_6_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h6] = int_rd_resp_desc_6_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h6] = int_rd_resp_desc_6_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h6] = int_rd_resp_desc_6_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h6] = int_rd_resp_desc_6_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h6] = int_wr_req_desc_6_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h6] = int_wr_req_desc_6_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h6] = int_wr_req_desc_6_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h6] = int_wr_req_desc_6_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h6] = int_wr_req_desc_6_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h6] = int_wr_req_desc_6_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h6] = int_wr_req_desc_6_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h6] = int_wr_req_desc_6_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h6] = int_wr_resp_desc_6_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h6] = int_wr_resp_desc_6_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h6] = int_wr_resp_desc_6_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h6] = int_wr_resp_desc_6_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h6] = int_wr_resp_desc_6_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h6] = int_wr_resp_desc_6_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h6] = int_wr_resp_desc_6_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h6] = int_wr_resp_desc_6_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h6] = int_wr_resp_desc_6_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h6] = int_wr_resp_desc_6_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h6] = int_wr_resp_desc_6_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h6] = int_wr_resp_desc_6_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h6] = int_wr_resp_desc_6_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h6] = int_wr_resp_desc_6_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h6] = int_wr_resp_desc_6_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h6] = int_wr_resp_desc_6_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h6] = int_wr_resp_desc_6_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h6] = int_wr_resp_desc_6_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h6] = int_wr_resp_desc_6_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h6] = int_wr_resp_desc_6_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h6] = int_wr_resp_desc_6_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h6] = int_sn_req_desc_6_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h6] = int_sn_req_desc_6_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h6] = int_sn_req_desc_6_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h6] = int_sn_req_desc_6_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h6] = int_sn_req_desc_6_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h6] = int_sn_req_desc_6_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h7] = int_rd_resp_desc_7_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h7] = int_rd_resp_desc_7_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h7] = int_rd_resp_desc_7_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h7] = int_rd_resp_desc_7_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h7] = int_rd_resp_desc_7_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h7] = int_rd_resp_desc_7_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h7] = int_rd_resp_desc_7_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h7] = int_rd_resp_desc_7_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h7] = int_rd_resp_desc_7_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h7] = int_rd_resp_desc_7_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h7] = int_rd_resp_desc_7_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h7] = int_rd_resp_desc_7_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h7] = int_rd_resp_desc_7_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h7] = int_rd_resp_desc_7_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h7] = int_rd_resp_desc_7_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h7] = int_rd_resp_desc_7_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h7] = int_rd_resp_desc_7_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h7] = int_rd_resp_desc_7_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h7] = int_rd_resp_desc_7_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h7] = int_rd_resp_desc_7_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h7] = int_rd_resp_desc_7_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h7] = int_rd_resp_desc_7_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h7] = int_rd_resp_desc_7_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h7] = int_rd_resp_desc_7_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h7] = int_rd_resp_desc_7_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h7] = int_rd_resp_desc_7_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h7] = int_rd_resp_desc_7_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h7] = int_wr_req_desc_7_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h7] = int_wr_req_desc_7_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h7] = int_wr_req_desc_7_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h7] = int_wr_req_desc_7_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h7] = int_wr_req_desc_7_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h7] = int_wr_req_desc_7_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h7] = int_wr_req_desc_7_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h7] = int_wr_req_desc_7_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h7] = int_wr_resp_desc_7_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h7] = int_wr_resp_desc_7_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h7] = int_wr_resp_desc_7_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h7] = int_wr_resp_desc_7_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h7] = int_wr_resp_desc_7_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h7] = int_wr_resp_desc_7_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h7] = int_wr_resp_desc_7_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h7] = int_wr_resp_desc_7_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h7] = int_wr_resp_desc_7_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h7] = int_wr_resp_desc_7_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h7] = int_wr_resp_desc_7_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h7] = int_wr_resp_desc_7_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h7] = int_wr_resp_desc_7_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h7] = int_wr_resp_desc_7_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h7] = int_wr_resp_desc_7_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h7] = int_wr_resp_desc_7_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h7] = int_wr_resp_desc_7_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h7] = int_wr_resp_desc_7_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h7] = int_wr_resp_desc_7_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h7] = int_wr_resp_desc_7_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h7] = int_wr_resp_desc_7_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h7] = int_sn_req_desc_7_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h7] = int_sn_req_desc_7_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h7] = int_sn_req_desc_7_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h7] = int_sn_req_desc_7_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h7] = int_sn_req_desc_7_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h7] = int_sn_req_desc_7_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h8] = int_rd_resp_desc_8_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h8] = int_rd_resp_desc_8_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h8] = int_rd_resp_desc_8_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h8] = int_rd_resp_desc_8_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h8] = int_rd_resp_desc_8_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h8] = int_rd_resp_desc_8_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h8] = int_rd_resp_desc_8_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h8] = int_rd_resp_desc_8_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h8] = int_rd_resp_desc_8_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h8] = int_rd_resp_desc_8_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h8] = int_rd_resp_desc_8_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h8] = int_rd_resp_desc_8_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h8] = int_rd_resp_desc_8_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h8] = int_rd_resp_desc_8_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h8] = int_rd_resp_desc_8_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h8] = int_rd_resp_desc_8_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h8] = int_rd_resp_desc_8_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h8] = int_rd_resp_desc_8_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h8] = int_rd_resp_desc_8_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h8] = int_rd_resp_desc_8_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h8] = int_rd_resp_desc_8_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h8] = int_rd_resp_desc_8_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h8] = int_rd_resp_desc_8_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h8] = int_rd_resp_desc_8_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h8] = int_rd_resp_desc_8_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h8] = int_rd_resp_desc_8_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h8] = int_rd_resp_desc_8_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h8] = int_wr_req_desc_8_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h8] = int_wr_req_desc_8_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h8] = int_wr_req_desc_8_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h8] = int_wr_req_desc_8_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h8] = int_wr_req_desc_8_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h8] = int_wr_req_desc_8_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h8] = int_wr_req_desc_8_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h8] = int_wr_req_desc_8_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h8] = int_wr_resp_desc_8_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h8] = int_wr_resp_desc_8_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h8] = int_wr_resp_desc_8_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h8] = int_wr_resp_desc_8_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h8] = int_wr_resp_desc_8_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h8] = int_wr_resp_desc_8_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h8] = int_wr_resp_desc_8_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h8] = int_wr_resp_desc_8_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h8] = int_wr_resp_desc_8_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h8] = int_wr_resp_desc_8_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h8] = int_wr_resp_desc_8_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h8] = int_wr_resp_desc_8_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h8] = int_wr_resp_desc_8_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h8] = int_wr_resp_desc_8_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h8] = int_wr_resp_desc_8_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h8] = int_wr_resp_desc_8_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h8] = int_wr_resp_desc_8_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h8] = int_wr_resp_desc_8_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h8] = int_wr_resp_desc_8_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h8] = int_wr_resp_desc_8_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h8] = int_wr_resp_desc_8_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h8] = int_sn_req_desc_8_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h8] = int_sn_req_desc_8_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h8] = int_sn_req_desc_8_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h8] = int_sn_req_desc_8_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h8] = int_sn_req_desc_8_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h8] = int_sn_req_desc_8_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['h9] = int_rd_resp_desc_9_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['h9] = int_rd_resp_desc_9_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['h9] = int_rd_resp_desc_9_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['h9] = int_rd_resp_desc_9_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['h9] = int_rd_resp_desc_9_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['h9] = int_rd_resp_desc_9_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['h9] = int_rd_resp_desc_9_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['h9] = int_rd_resp_desc_9_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['h9] = int_rd_resp_desc_9_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['h9] = int_rd_resp_desc_9_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['h9] = int_rd_resp_desc_9_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['h9] = int_rd_resp_desc_9_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['h9] = int_rd_resp_desc_9_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['h9] = int_rd_resp_desc_9_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['h9] = int_rd_resp_desc_9_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['h9] = int_rd_resp_desc_9_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['h9] = int_rd_resp_desc_9_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['h9] = int_rd_resp_desc_9_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['h9] = int_rd_resp_desc_9_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['h9] = int_rd_resp_desc_9_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['h9] = int_rd_resp_desc_9_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['h9] = int_rd_resp_desc_9_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['h9] = int_rd_resp_desc_9_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['h9] = int_rd_resp_desc_9_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['h9] = int_rd_resp_desc_9_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['h9] = int_rd_resp_desc_9_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['h9] = int_rd_resp_desc_9_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['h9] = int_wr_req_desc_9_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['h9] = int_wr_req_desc_9_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['h9] = int_wr_req_desc_9_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['h9] = int_wr_req_desc_9_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['h9] = int_wr_req_desc_9_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['h9] = int_wr_req_desc_9_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['h9] = int_wr_req_desc_9_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['h9] = int_wr_req_desc_9_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['h9] = int_wr_resp_desc_9_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['h9] = int_wr_resp_desc_9_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['h9] = int_wr_resp_desc_9_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['h9] = int_wr_resp_desc_9_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['h9] = int_wr_resp_desc_9_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['h9] = int_wr_resp_desc_9_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['h9] = int_wr_resp_desc_9_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['h9] = int_wr_resp_desc_9_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['h9] = int_wr_resp_desc_9_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['h9] = int_wr_resp_desc_9_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['h9] = int_wr_resp_desc_9_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['h9] = int_wr_resp_desc_9_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['h9] = int_wr_resp_desc_9_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['h9] = int_wr_resp_desc_9_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['h9] = int_wr_resp_desc_9_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['h9] = int_wr_resp_desc_9_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['h9] = int_wr_resp_desc_9_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['h9] = int_wr_resp_desc_9_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['h9] = int_wr_resp_desc_9_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['h9] = int_wr_resp_desc_9_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['h9] = int_wr_resp_desc_9_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['h9] = int_sn_req_desc_9_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['h9] = int_sn_req_desc_9_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['h9] = int_sn_req_desc_9_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['h9] = int_sn_req_desc_9_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['h9] = int_sn_req_desc_9_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['h9] = int_sn_req_desc_9_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['ha] = int_rd_resp_desc_a_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['ha] = int_rd_resp_desc_a_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['ha] = int_rd_resp_desc_a_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['ha] = int_rd_resp_desc_a_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['ha] = int_rd_resp_desc_a_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['ha] = int_rd_resp_desc_a_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['ha] = int_rd_resp_desc_a_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['ha] = int_rd_resp_desc_a_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['ha] = int_rd_resp_desc_a_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['ha] = int_rd_resp_desc_a_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['ha] = int_rd_resp_desc_a_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['ha] = int_rd_resp_desc_a_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['ha] = int_rd_resp_desc_a_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['ha] = int_rd_resp_desc_a_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['ha] = int_rd_resp_desc_a_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['ha] = int_rd_resp_desc_a_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['ha] = int_rd_resp_desc_a_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['ha] = int_rd_resp_desc_a_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['ha] = int_rd_resp_desc_a_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['ha] = int_rd_resp_desc_a_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['ha] = int_rd_resp_desc_a_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['ha] = int_rd_resp_desc_a_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['ha] = int_rd_resp_desc_a_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['ha] = int_rd_resp_desc_a_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['ha] = int_rd_resp_desc_a_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['ha] = int_rd_resp_desc_a_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['ha] = int_rd_resp_desc_a_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['ha] = int_wr_req_desc_a_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['ha] = int_wr_req_desc_a_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['ha] = int_wr_req_desc_a_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['ha] = int_wr_req_desc_a_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['ha] = int_wr_req_desc_a_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['ha] = int_wr_req_desc_a_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['ha] = int_wr_req_desc_a_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['ha] = int_wr_req_desc_a_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['ha] = int_wr_resp_desc_a_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['ha] = int_wr_resp_desc_a_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['ha] = int_wr_resp_desc_a_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['ha] = int_wr_resp_desc_a_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['ha] = int_wr_resp_desc_a_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['ha] = int_wr_resp_desc_a_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['ha] = int_wr_resp_desc_a_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['ha] = int_wr_resp_desc_a_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['ha] = int_wr_resp_desc_a_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['ha] = int_wr_resp_desc_a_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['ha] = int_wr_resp_desc_a_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['ha] = int_wr_resp_desc_a_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['ha] = int_wr_resp_desc_a_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['ha] = int_wr_resp_desc_a_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['ha] = int_wr_resp_desc_a_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['ha] = int_wr_resp_desc_a_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['ha] = int_wr_resp_desc_a_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['ha] = int_wr_resp_desc_a_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['ha] = int_wr_resp_desc_a_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['ha] = int_wr_resp_desc_a_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['ha] = int_wr_resp_desc_a_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['ha] = int_sn_req_desc_a_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['ha] = int_sn_req_desc_a_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['ha] = int_sn_req_desc_a_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['ha] = int_sn_req_desc_a_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['ha] = int_sn_req_desc_a_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['ha] = int_sn_req_desc_a_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['hb] = int_rd_resp_desc_b_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['hb] = int_rd_resp_desc_b_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['hb] = int_rd_resp_desc_b_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['hb] = int_rd_resp_desc_b_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['hb] = int_rd_resp_desc_b_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['hb] = int_rd_resp_desc_b_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['hb] = int_rd_resp_desc_b_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['hb] = int_rd_resp_desc_b_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['hb] = int_rd_resp_desc_b_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['hb] = int_rd_resp_desc_b_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['hb] = int_rd_resp_desc_b_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['hb] = int_rd_resp_desc_b_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['hb] = int_rd_resp_desc_b_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['hb] = int_rd_resp_desc_b_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['hb] = int_rd_resp_desc_b_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['hb] = int_rd_resp_desc_b_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['hb] = int_rd_resp_desc_b_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['hb] = int_rd_resp_desc_b_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['hb] = int_rd_resp_desc_b_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['hb] = int_rd_resp_desc_b_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['hb] = int_rd_resp_desc_b_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['hb] = int_rd_resp_desc_b_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['hb] = int_rd_resp_desc_b_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['hb] = int_rd_resp_desc_b_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['hb] = int_rd_resp_desc_b_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['hb] = int_rd_resp_desc_b_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['hb] = int_rd_resp_desc_b_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['hb] = int_wr_req_desc_b_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['hb] = int_wr_req_desc_b_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['hb] = int_wr_req_desc_b_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['hb] = int_wr_req_desc_b_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['hb] = int_wr_req_desc_b_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['hb] = int_wr_req_desc_b_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['hb] = int_wr_req_desc_b_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['hb] = int_wr_req_desc_b_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['hb] = int_wr_resp_desc_b_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['hb] = int_wr_resp_desc_b_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['hb] = int_wr_resp_desc_b_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['hb] = int_wr_resp_desc_b_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['hb] = int_wr_resp_desc_b_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['hb] = int_wr_resp_desc_b_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['hb] = int_wr_resp_desc_b_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['hb] = int_wr_resp_desc_b_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['hb] = int_wr_resp_desc_b_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['hb] = int_wr_resp_desc_b_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['hb] = int_wr_resp_desc_b_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['hb] = int_wr_resp_desc_b_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['hb] = int_wr_resp_desc_b_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['hb] = int_wr_resp_desc_b_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['hb] = int_wr_resp_desc_b_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['hb] = int_wr_resp_desc_b_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['hb] = int_wr_resp_desc_b_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['hb] = int_wr_resp_desc_b_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['hb] = int_wr_resp_desc_b_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['hb] = int_wr_resp_desc_b_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['hb] = int_wr_resp_desc_b_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['hb] = int_sn_req_desc_b_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['hb] = int_sn_req_desc_b_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['hb] = int_sn_req_desc_b_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['hb] = int_sn_req_desc_b_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['hb] = int_sn_req_desc_b_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['hb] = int_sn_req_desc_b_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['hc] = int_rd_resp_desc_c_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['hc] = int_rd_resp_desc_c_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['hc] = int_rd_resp_desc_c_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['hc] = int_rd_resp_desc_c_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['hc] = int_rd_resp_desc_c_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['hc] = int_rd_resp_desc_c_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['hc] = int_rd_resp_desc_c_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['hc] = int_rd_resp_desc_c_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['hc] = int_rd_resp_desc_c_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['hc] = int_rd_resp_desc_c_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['hc] = int_rd_resp_desc_c_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['hc] = int_rd_resp_desc_c_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['hc] = int_rd_resp_desc_c_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['hc] = int_rd_resp_desc_c_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['hc] = int_rd_resp_desc_c_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['hc] = int_rd_resp_desc_c_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['hc] = int_rd_resp_desc_c_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['hc] = int_rd_resp_desc_c_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['hc] = int_rd_resp_desc_c_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['hc] = int_rd_resp_desc_c_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['hc] = int_rd_resp_desc_c_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['hc] = int_rd_resp_desc_c_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['hc] = int_rd_resp_desc_c_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['hc] = int_rd_resp_desc_c_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['hc] = int_rd_resp_desc_c_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['hc] = int_rd_resp_desc_c_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['hc] = int_rd_resp_desc_c_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['hc] = int_wr_req_desc_c_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['hc] = int_wr_req_desc_c_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['hc] = int_wr_req_desc_c_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['hc] = int_wr_req_desc_c_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['hc] = int_wr_req_desc_c_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['hc] = int_wr_req_desc_c_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['hc] = int_wr_req_desc_c_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['hc] = int_wr_req_desc_c_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['hc] = int_wr_resp_desc_c_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['hc] = int_wr_resp_desc_c_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['hc] = int_wr_resp_desc_c_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['hc] = int_wr_resp_desc_c_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['hc] = int_wr_resp_desc_c_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['hc] = int_wr_resp_desc_c_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['hc] = int_wr_resp_desc_c_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['hc] = int_wr_resp_desc_c_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['hc] = int_wr_resp_desc_c_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['hc] = int_wr_resp_desc_c_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['hc] = int_wr_resp_desc_c_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['hc] = int_wr_resp_desc_c_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['hc] = int_wr_resp_desc_c_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['hc] = int_wr_resp_desc_c_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['hc] = int_wr_resp_desc_c_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['hc] = int_wr_resp_desc_c_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['hc] = int_wr_resp_desc_c_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['hc] = int_wr_resp_desc_c_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['hc] = int_wr_resp_desc_c_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['hc] = int_wr_resp_desc_c_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['hc] = int_wr_resp_desc_c_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['hc] = int_sn_req_desc_c_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['hc] = int_sn_req_desc_c_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['hc] = int_sn_req_desc_c_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['hc] = int_sn_req_desc_c_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['hc] = int_sn_req_desc_c_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['hc] = int_sn_req_desc_c_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['hd] = int_rd_resp_desc_d_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['hd] = int_rd_resp_desc_d_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['hd] = int_rd_resp_desc_d_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['hd] = int_rd_resp_desc_d_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['hd] = int_rd_resp_desc_d_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['hd] = int_rd_resp_desc_d_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['hd] = int_rd_resp_desc_d_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['hd] = int_rd_resp_desc_d_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['hd] = int_rd_resp_desc_d_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['hd] = int_rd_resp_desc_d_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['hd] = int_rd_resp_desc_d_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['hd] = int_rd_resp_desc_d_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['hd] = int_rd_resp_desc_d_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['hd] = int_rd_resp_desc_d_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['hd] = int_rd_resp_desc_d_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['hd] = int_rd_resp_desc_d_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['hd] = int_rd_resp_desc_d_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['hd] = int_rd_resp_desc_d_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['hd] = int_rd_resp_desc_d_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['hd] = int_rd_resp_desc_d_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['hd] = int_rd_resp_desc_d_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['hd] = int_rd_resp_desc_d_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['hd] = int_rd_resp_desc_d_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['hd] = int_rd_resp_desc_d_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['hd] = int_rd_resp_desc_d_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['hd] = int_rd_resp_desc_d_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['hd] = int_rd_resp_desc_d_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['hd] = int_wr_req_desc_d_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['hd] = int_wr_req_desc_d_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['hd] = int_wr_req_desc_d_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['hd] = int_wr_req_desc_d_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['hd] = int_wr_req_desc_d_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['hd] = int_wr_req_desc_d_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['hd] = int_wr_req_desc_d_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['hd] = int_wr_req_desc_d_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['hd] = int_wr_resp_desc_d_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['hd] = int_wr_resp_desc_d_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['hd] = int_wr_resp_desc_d_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['hd] = int_wr_resp_desc_d_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['hd] = int_wr_resp_desc_d_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['hd] = int_wr_resp_desc_d_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['hd] = int_wr_resp_desc_d_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['hd] = int_wr_resp_desc_d_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['hd] = int_wr_resp_desc_d_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['hd] = int_wr_resp_desc_d_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['hd] = int_wr_resp_desc_d_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['hd] = int_wr_resp_desc_d_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['hd] = int_wr_resp_desc_d_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['hd] = int_wr_resp_desc_d_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['hd] = int_wr_resp_desc_d_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['hd] = int_wr_resp_desc_d_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['hd] = int_wr_resp_desc_d_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['hd] = int_wr_resp_desc_d_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['hd] = int_wr_resp_desc_d_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['hd] = int_wr_resp_desc_d_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['hd] = int_wr_resp_desc_d_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['hd] = int_sn_req_desc_d_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['hd] = int_sn_req_desc_d_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['hd] = int_sn_req_desc_d_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['hd] = int_sn_req_desc_d_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['hd] = int_sn_req_desc_d_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['hd] = int_sn_req_desc_d_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['he] = int_rd_resp_desc_e_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['he] = int_rd_resp_desc_e_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['he] = int_rd_resp_desc_e_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['he] = int_rd_resp_desc_e_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['he] = int_rd_resp_desc_e_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['he] = int_rd_resp_desc_e_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['he] = int_rd_resp_desc_e_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['he] = int_rd_resp_desc_e_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['he] = int_rd_resp_desc_e_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['he] = int_rd_resp_desc_e_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['he] = int_rd_resp_desc_e_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['he] = int_rd_resp_desc_e_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['he] = int_rd_resp_desc_e_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['he] = int_rd_resp_desc_e_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['he] = int_rd_resp_desc_e_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['he] = int_rd_resp_desc_e_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['he] = int_rd_resp_desc_e_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['he] = int_rd_resp_desc_e_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['he] = int_rd_resp_desc_e_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['he] = int_rd_resp_desc_e_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['he] = int_rd_resp_desc_e_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['he] = int_rd_resp_desc_e_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['he] = int_rd_resp_desc_e_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['he] = int_rd_resp_desc_e_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['he] = int_rd_resp_desc_e_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['he] = int_rd_resp_desc_e_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['he] = int_rd_resp_desc_e_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['he] = int_wr_req_desc_e_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['he] = int_wr_req_desc_e_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['he] = int_wr_req_desc_e_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['he] = int_wr_req_desc_e_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['he] = int_wr_req_desc_e_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['he] = int_wr_req_desc_e_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['he] = int_wr_req_desc_e_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['he] = int_wr_req_desc_e_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['he] = int_wr_resp_desc_e_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['he] = int_wr_resp_desc_e_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['he] = int_wr_resp_desc_e_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['he] = int_wr_resp_desc_e_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['he] = int_wr_resp_desc_e_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['he] = int_wr_resp_desc_e_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['he] = int_wr_resp_desc_e_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['he] = int_wr_resp_desc_e_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['he] = int_wr_resp_desc_e_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['he] = int_wr_resp_desc_e_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['he] = int_wr_resp_desc_e_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['he] = int_wr_resp_desc_e_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['he] = int_wr_resp_desc_e_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['he] = int_wr_resp_desc_e_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['he] = int_wr_resp_desc_e_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['he] = int_wr_resp_desc_e_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['he] = int_wr_resp_desc_e_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['he] = int_wr_resp_desc_e_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['he] = int_wr_resp_desc_e_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['he] = int_wr_resp_desc_e_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['he] = int_wr_resp_desc_e_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['he] = int_sn_req_desc_e_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['he] = int_sn_req_desc_e_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['he] = int_sn_req_desc_e_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['he] = int_sn_req_desc_e_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['he] = int_sn_req_desc_e_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['he] = int_sn_req_desc_e_acaddr_3_addr;
assign int_rd_resp_desc_n_data_offset_addr['hf] = int_rd_resp_desc_f_data_offset_addr;
assign int_rd_resp_desc_n_data_size_size['hf] = int_rd_resp_desc_f_data_size_size;
assign int_rd_resp_desc_n_data_host_addr_0_addr['hf] = int_rd_resp_desc_f_data_host_addr_0_addr;
assign int_rd_resp_desc_n_data_host_addr_1_addr['hf] = int_rd_resp_desc_f_data_host_addr_1_addr;
assign int_rd_resp_desc_n_data_host_addr_2_addr['hf] = int_rd_resp_desc_f_data_host_addr_2_addr;
assign int_rd_resp_desc_n_data_host_addr_3_addr['hf] = int_rd_resp_desc_f_data_host_addr_3_addr;
assign int_rd_resp_desc_n_resp_resp['hf] = int_rd_resp_desc_f_resp_resp;
assign int_rd_resp_desc_n_xid_0_xid['hf] = int_rd_resp_desc_f_xid_0_xid;
assign int_rd_resp_desc_n_xid_1_xid['hf] = int_rd_resp_desc_f_xid_1_xid;
assign int_rd_resp_desc_n_xid_2_xid['hf] = int_rd_resp_desc_f_xid_2_xid;
assign int_rd_resp_desc_n_xid_3_xid['hf] = int_rd_resp_desc_f_xid_3_xid;
assign int_rd_resp_desc_n_xuser_0_xuser['hf] = int_rd_resp_desc_f_xuser_0_xuser;
assign int_rd_resp_desc_n_xuser_1_xuser['hf] = int_rd_resp_desc_f_xuser_1_xuser;
assign int_rd_resp_desc_n_xuser_2_xuser['hf] = int_rd_resp_desc_f_xuser_2_xuser;
assign int_rd_resp_desc_n_xuser_3_xuser['hf] = int_rd_resp_desc_f_xuser_3_xuser;
assign int_rd_resp_desc_n_xuser_4_xuser['hf] = int_rd_resp_desc_f_xuser_4_xuser;
assign int_rd_resp_desc_n_xuser_5_xuser['hf] = int_rd_resp_desc_f_xuser_5_xuser;
assign int_rd_resp_desc_n_xuser_6_xuser['hf] = int_rd_resp_desc_f_xuser_6_xuser;
assign int_rd_resp_desc_n_xuser_7_xuser['hf] = int_rd_resp_desc_f_xuser_7_xuser;
assign int_rd_resp_desc_n_xuser_8_xuser['hf] = int_rd_resp_desc_f_xuser_8_xuser;
assign int_rd_resp_desc_n_xuser_9_xuser['hf] = int_rd_resp_desc_f_xuser_9_xuser;
assign int_rd_resp_desc_n_xuser_10_xuser['hf] = int_rd_resp_desc_f_xuser_10_xuser;
assign int_rd_resp_desc_n_xuser_11_xuser['hf] = int_rd_resp_desc_f_xuser_11_xuser;
assign int_rd_resp_desc_n_xuser_12_xuser['hf] = int_rd_resp_desc_f_xuser_12_xuser;
assign int_rd_resp_desc_n_xuser_13_xuser['hf] = int_rd_resp_desc_f_xuser_13_xuser;
assign int_rd_resp_desc_n_xuser_14_xuser['hf] = int_rd_resp_desc_f_xuser_14_xuser;
assign int_rd_resp_desc_n_xuser_15_xuser['hf] = int_rd_resp_desc_f_xuser_15_xuser;
assign int_wr_req_desc_n_data_host_addr_0_addr['hf] = int_wr_req_desc_f_data_host_addr_0_addr;
assign int_wr_req_desc_n_data_host_addr_1_addr['hf] = int_wr_req_desc_f_data_host_addr_1_addr;
assign int_wr_req_desc_n_data_host_addr_2_addr['hf] = int_wr_req_desc_f_data_host_addr_2_addr;
assign int_wr_req_desc_n_data_host_addr_3_addr['hf] = int_wr_req_desc_f_data_host_addr_3_addr;
assign int_wr_req_desc_n_wstrb_host_addr_0_addr['hf] = int_wr_req_desc_f_wstrb_host_addr_0_addr;
assign int_wr_req_desc_n_wstrb_host_addr_1_addr['hf] = int_wr_req_desc_f_wstrb_host_addr_1_addr;
assign int_wr_req_desc_n_wstrb_host_addr_2_addr['hf] = int_wr_req_desc_f_wstrb_host_addr_2_addr;
assign int_wr_req_desc_n_wstrb_host_addr_3_addr['hf] = int_wr_req_desc_f_wstrb_host_addr_3_addr;
assign int_wr_resp_desc_n_resp_resp['hf] = int_wr_resp_desc_f_resp_resp;
assign int_wr_resp_desc_n_xid_0_xid['hf] = int_wr_resp_desc_f_xid_0_xid;
assign int_wr_resp_desc_n_xid_1_xid['hf] = int_wr_resp_desc_f_xid_1_xid;
assign int_wr_resp_desc_n_xid_2_xid['hf] = int_wr_resp_desc_f_xid_2_xid;
assign int_wr_resp_desc_n_xid_3_xid['hf] = int_wr_resp_desc_f_xid_3_xid;
assign int_wr_resp_desc_n_xuser_0_xuser['hf] = int_wr_resp_desc_f_xuser_0_xuser;
assign int_wr_resp_desc_n_xuser_1_xuser['hf] = int_wr_resp_desc_f_xuser_1_xuser;
assign int_wr_resp_desc_n_xuser_2_xuser['hf] = int_wr_resp_desc_f_xuser_2_xuser;
assign int_wr_resp_desc_n_xuser_3_xuser['hf] = int_wr_resp_desc_f_xuser_3_xuser;
assign int_wr_resp_desc_n_xuser_4_xuser['hf] = int_wr_resp_desc_f_xuser_4_xuser;
assign int_wr_resp_desc_n_xuser_5_xuser['hf] = int_wr_resp_desc_f_xuser_5_xuser;
assign int_wr_resp_desc_n_xuser_6_xuser['hf] = int_wr_resp_desc_f_xuser_6_xuser;
assign int_wr_resp_desc_n_xuser_7_xuser['hf] = int_wr_resp_desc_f_xuser_7_xuser;
assign int_wr_resp_desc_n_xuser_8_xuser['hf] = int_wr_resp_desc_f_xuser_8_xuser;
assign int_wr_resp_desc_n_xuser_9_xuser['hf] = int_wr_resp_desc_f_xuser_9_xuser;
assign int_wr_resp_desc_n_xuser_10_xuser['hf] = int_wr_resp_desc_f_xuser_10_xuser;
assign int_wr_resp_desc_n_xuser_11_xuser['hf] = int_wr_resp_desc_f_xuser_11_xuser;
assign int_wr_resp_desc_n_xuser_12_xuser['hf] = int_wr_resp_desc_f_xuser_12_xuser;
assign int_wr_resp_desc_n_xuser_13_xuser['hf] = int_wr_resp_desc_f_xuser_13_xuser;
assign int_wr_resp_desc_n_xuser_14_xuser['hf] = int_wr_resp_desc_f_xuser_14_xuser;
assign int_wr_resp_desc_n_xuser_15_xuser['hf] = int_wr_resp_desc_f_xuser_15_xuser;
assign int_sn_req_desc_n_attr_acsnoop['hf] = int_sn_req_desc_f_attr_acsnoop;
assign int_sn_req_desc_n_attr_acprot['hf] = int_sn_req_desc_f_attr_acprot;
assign int_sn_req_desc_n_acaddr_0_addr['hf] = int_sn_req_desc_f_acaddr_0_addr;
assign int_sn_req_desc_n_acaddr_1_addr['hf] = int_sn_req_desc_f_acaddr_1_addr;
assign int_sn_req_desc_n_acaddr_2_addr['hf] = int_sn_req_desc_f_acaddr_2_addr;
assign int_sn_req_desc_n_acaddr_3_addr['hf] = int_sn_req_desc_f_acaddr_3_addr;

