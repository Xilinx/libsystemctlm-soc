/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */

        ,output [0:0]	int_desc_0_txn_type_wr_strb
        ,output [0:0]	int_desc_0_txn_type_wr_rd
        ,output [3:0]	int_desc_0_attr_axregion
        ,output [3:0]	int_desc_0_attr_axqos
        ,output [2:0]	int_desc_0_attr_axprot
        ,output [3:0]	int_desc_0_attr_axcache
        ,output [1:0]	int_desc_0_attr_axlock
        ,output [1:0]	int_desc_0_attr_axburst
        ,output [31:0]	int_desc_0_axid_0_axid
        ,output [31:0]	int_desc_0_axid_1_axid
        ,output [31:0]	int_desc_0_axid_2_axid
        ,output [31:0]	int_desc_0_axid_3_axid
        ,output [31:0]	int_desc_0_axuser_0_axuser
        ,output [31:0]	int_desc_0_axuser_1_axuser
        ,output [31:0]	int_desc_0_axuser_2_axuser
        ,output [31:0]	int_desc_0_axuser_3_axuser
        ,output [31:0]	int_desc_0_axuser_4_axuser
        ,output [31:0]	int_desc_0_axuser_5_axuser
        ,output [31:0]	int_desc_0_axuser_6_axuser
        ,output [31:0]	int_desc_0_axuser_7_axuser
        ,output [31:0]	int_desc_0_axuser_8_axuser
        ,output [31:0]	int_desc_0_axuser_9_axuser
        ,output [31:0]	int_desc_0_axuser_10_axuser
        ,output [31:0]	int_desc_0_axuser_11_axuser
        ,output [31:0]	int_desc_0_axuser_12_axuser
        ,output [31:0]	int_desc_0_axuser_13_axuser
        ,output [31:0]	int_desc_0_axuser_14_axuser
        ,output [31:0]	int_desc_0_axuser_15_axuser
        ,output [15:0]	int_desc_0_size_txn_size
        ,output [2:0]	int_desc_0_axsize_axsize
        ,output [31:0]	int_desc_0_axaddr_0_addr
        ,output [31:0]	int_desc_0_axaddr_1_addr
        ,output [31:0]	int_desc_0_axaddr_2_addr
        ,output [31:0]	int_desc_0_axaddr_3_addr
        ,output [31:0]	int_desc_0_data_offset_addr
        ,output [31:0]	int_desc_0_wuser_0_wuser
        ,output [31:0]	int_desc_0_wuser_1_wuser
        ,output [31:0]	int_desc_0_wuser_2_wuser
        ,output [31:0]	int_desc_0_wuser_3_wuser
        ,output [31:0]	int_desc_0_wuser_4_wuser
        ,output [31:0]	int_desc_0_wuser_5_wuser
        ,output [31:0]	int_desc_0_wuser_6_wuser
        ,output [31:0]	int_desc_0_wuser_7_wuser
        ,output [31:0]	int_desc_0_wuser_8_wuser
        ,output [31:0]	int_desc_0_wuser_9_wuser
        ,output [31:0]	int_desc_0_wuser_10_wuser
        ,output [31:0]	int_desc_0_wuser_11_wuser
        ,output [31:0]	int_desc_0_wuser_12_wuser
        ,output [31:0]	int_desc_0_wuser_13_wuser
        ,output [31:0]	int_desc_0_wuser_14_wuser
        ,output [31:0]	int_desc_0_wuser_15_wuser
        ,output [0:0]	int_desc_1_txn_type_wr_strb
        ,output [0:0]	int_desc_1_txn_type_wr_rd
        ,output [3:0]	int_desc_1_attr_axregion
        ,output [3:0]	int_desc_1_attr_axqos
        ,output [2:0]	int_desc_1_attr_axprot
        ,output [3:0]	int_desc_1_attr_axcache
        ,output [1:0]	int_desc_1_attr_axlock
        ,output [1:0]	int_desc_1_attr_axburst
        ,output [31:0]	int_desc_1_axid_0_axid
        ,output [31:0]	int_desc_1_axid_1_axid
        ,output [31:0]	int_desc_1_axid_2_axid
        ,output [31:0]	int_desc_1_axid_3_axid
        ,output [31:0]	int_desc_1_axuser_0_axuser
        ,output [31:0]	int_desc_1_axuser_1_axuser
        ,output [31:0]	int_desc_1_axuser_2_axuser
        ,output [31:0]	int_desc_1_axuser_3_axuser
        ,output [31:0]	int_desc_1_axuser_4_axuser
        ,output [31:0]	int_desc_1_axuser_5_axuser
        ,output [31:0]	int_desc_1_axuser_6_axuser
        ,output [31:0]	int_desc_1_axuser_7_axuser
        ,output [31:0]	int_desc_1_axuser_8_axuser
        ,output [31:0]	int_desc_1_axuser_9_axuser
        ,output [31:0]	int_desc_1_axuser_10_axuser
        ,output [31:0]	int_desc_1_axuser_11_axuser
        ,output [31:0]	int_desc_1_axuser_12_axuser
        ,output [31:0]	int_desc_1_axuser_13_axuser
        ,output [31:0]	int_desc_1_axuser_14_axuser
        ,output [31:0]	int_desc_1_axuser_15_axuser
        ,output [15:0]	int_desc_1_size_txn_size
        ,output [2:0]	int_desc_1_axsize_axsize
        ,output [31:0]	int_desc_1_axaddr_0_addr
        ,output [31:0]	int_desc_1_axaddr_1_addr
        ,output [31:0]	int_desc_1_axaddr_2_addr
        ,output [31:0]	int_desc_1_axaddr_3_addr
        ,output [31:0]	int_desc_1_data_offset_addr
        ,output [31:0]	int_desc_1_wuser_0_wuser
        ,output [31:0]	int_desc_1_wuser_1_wuser
        ,output [31:0]	int_desc_1_wuser_2_wuser
        ,output [31:0]	int_desc_1_wuser_3_wuser
        ,output [31:0]	int_desc_1_wuser_4_wuser
        ,output [31:0]	int_desc_1_wuser_5_wuser
        ,output [31:0]	int_desc_1_wuser_6_wuser
        ,output [31:0]	int_desc_1_wuser_7_wuser
        ,output [31:0]	int_desc_1_wuser_8_wuser
        ,output [31:0]	int_desc_1_wuser_9_wuser
        ,output [31:0]	int_desc_1_wuser_10_wuser
        ,output [31:0]	int_desc_1_wuser_11_wuser
        ,output [31:0]	int_desc_1_wuser_12_wuser
        ,output [31:0]	int_desc_1_wuser_13_wuser
        ,output [31:0]	int_desc_1_wuser_14_wuser
        ,output [31:0]	int_desc_1_wuser_15_wuser
        ,output [0:0]	int_desc_2_txn_type_wr_strb
        ,output [0:0]	int_desc_2_txn_type_wr_rd
        ,output [3:0]	int_desc_2_attr_axregion
        ,output [3:0]	int_desc_2_attr_axqos
        ,output [2:0]	int_desc_2_attr_axprot
        ,output [3:0]	int_desc_2_attr_axcache
        ,output [1:0]	int_desc_2_attr_axlock
        ,output [1:0]	int_desc_2_attr_axburst
        ,output [31:0]	int_desc_2_axid_0_axid
        ,output [31:0]	int_desc_2_axid_1_axid
        ,output [31:0]	int_desc_2_axid_2_axid
        ,output [31:0]	int_desc_2_axid_3_axid
        ,output [31:0]	int_desc_2_axuser_0_axuser
        ,output [31:0]	int_desc_2_axuser_1_axuser
        ,output [31:0]	int_desc_2_axuser_2_axuser
        ,output [31:0]	int_desc_2_axuser_3_axuser
        ,output [31:0]	int_desc_2_axuser_4_axuser
        ,output [31:0]	int_desc_2_axuser_5_axuser
        ,output [31:0]	int_desc_2_axuser_6_axuser
        ,output [31:0]	int_desc_2_axuser_7_axuser
        ,output [31:0]	int_desc_2_axuser_8_axuser
        ,output [31:0]	int_desc_2_axuser_9_axuser
        ,output [31:0]	int_desc_2_axuser_10_axuser
        ,output [31:0]	int_desc_2_axuser_11_axuser
        ,output [31:0]	int_desc_2_axuser_12_axuser
        ,output [31:0]	int_desc_2_axuser_13_axuser
        ,output [31:0]	int_desc_2_axuser_14_axuser
        ,output [31:0]	int_desc_2_axuser_15_axuser
        ,output [15:0]	int_desc_2_size_txn_size
        ,output [2:0]	int_desc_2_axsize_axsize
        ,output [31:0]	int_desc_2_axaddr_0_addr
        ,output [31:0]	int_desc_2_axaddr_1_addr
        ,output [31:0]	int_desc_2_axaddr_2_addr
        ,output [31:0]	int_desc_2_axaddr_3_addr
        ,output [31:0]	int_desc_2_data_offset_addr
        ,output [31:0]	int_desc_2_wuser_0_wuser
        ,output [31:0]	int_desc_2_wuser_1_wuser
        ,output [31:0]	int_desc_2_wuser_2_wuser
        ,output [31:0]	int_desc_2_wuser_3_wuser
        ,output [31:0]	int_desc_2_wuser_4_wuser
        ,output [31:0]	int_desc_2_wuser_5_wuser
        ,output [31:0]	int_desc_2_wuser_6_wuser
        ,output [31:0]	int_desc_2_wuser_7_wuser
        ,output [31:0]	int_desc_2_wuser_8_wuser
        ,output [31:0]	int_desc_2_wuser_9_wuser
        ,output [31:0]	int_desc_2_wuser_10_wuser
        ,output [31:0]	int_desc_2_wuser_11_wuser
        ,output [31:0]	int_desc_2_wuser_12_wuser
        ,output [31:0]	int_desc_2_wuser_13_wuser
        ,output [31:0]	int_desc_2_wuser_14_wuser
        ,output [31:0]	int_desc_2_wuser_15_wuser
        ,output [0:0]	int_desc_3_txn_type_wr_strb
        ,output [0:0]	int_desc_3_txn_type_wr_rd
        ,output [3:0]	int_desc_3_attr_axregion
        ,output [3:0]	int_desc_3_attr_axqos
        ,output [2:0]	int_desc_3_attr_axprot
        ,output [3:0]	int_desc_3_attr_axcache
        ,output [1:0]	int_desc_3_attr_axlock
        ,output [1:0]	int_desc_3_attr_axburst
        ,output [31:0]	int_desc_3_axid_0_axid
        ,output [31:0]	int_desc_3_axid_1_axid
        ,output [31:0]	int_desc_3_axid_2_axid
        ,output [31:0]	int_desc_3_axid_3_axid
        ,output [31:0]	int_desc_3_axuser_0_axuser
        ,output [31:0]	int_desc_3_axuser_1_axuser
        ,output [31:0]	int_desc_3_axuser_2_axuser
        ,output [31:0]	int_desc_3_axuser_3_axuser
        ,output [31:0]	int_desc_3_axuser_4_axuser
        ,output [31:0]	int_desc_3_axuser_5_axuser
        ,output [31:0]	int_desc_3_axuser_6_axuser
        ,output [31:0]	int_desc_3_axuser_7_axuser
        ,output [31:0]	int_desc_3_axuser_8_axuser
        ,output [31:0]	int_desc_3_axuser_9_axuser
        ,output [31:0]	int_desc_3_axuser_10_axuser
        ,output [31:0]	int_desc_3_axuser_11_axuser
        ,output [31:0]	int_desc_3_axuser_12_axuser
        ,output [31:0]	int_desc_3_axuser_13_axuser
        ,output [31:0]	int_desc_3_axuser_14_axuser
        ,output [31:0]	int_desc_3_axuser_15_axuser
        ,output [15:0]	int_desc_3_size_txn_size
        ,output [2:0]	int_desc_3_axsize_axsize
        ,output [31:0]	int_desc_3_axaddr_0_addr
        ,output [31:0]	int_desc_3_axaddr_1_addr
        ,output [31:0]	int_desc_3_axaddr_2_addr
        ,output [31:0]	int_desc_3_axaddr_3_addr
        ,output [31:0]	int_desc_3_data_offset_addr
        ,output [31:0]	int_desc_3_wuser_0_wuser
        ,output [31:0]	int_desc_3_wuser_1_wuser
        ,output [31:0]	int_desc_3_wuser_2_wuser
        ,output [31:0]	int_desc_3_wuser_3_wuser
        ,output [31:0]	int_desc_3_wuser_4_wuser
        ,output [31:0]	int_desc_3_wuser_5_wuser
        ,output [31:0]	int_desc_3_wuser_6_wuser
        ,output [31:0]	int_desc_3_wuser_7_wuser
        ,output [31:0]	int_desc_3_wuser_8_wuser
        ,output [31:0]	int_desc_3_wuser_9_wuser
        ,output [31:0]	int_desc_3_wuser_10_wuser
        ,output [31:0]	int_desc_3_wuser_11_wuser
        ,output [31:0]	int_desc_3_wuser_12_wuser
        ,output [31:0]	int_desc_3_wuser_13_wuser
        ,output [31:0]	int_desc_3_wuser_14_wuser
        ,output [31:0]	int_desc_3_wuser_15_wuser
        ,output [0:0]	int_desc_4_txn_type_wr_strb
        ,output [0:0]	int_desc_4_txn_type_wr_rd
        ,output [3:0]	int_desc_4_attr_axregion
        ,output [3:0]	int_desc_4_attr_axqos
        ,output [2:0]	int_desc_4_attr_axprot
        ,output [3:0]	int_desc_4_attr_axcache
        ,output [1:0]	int_desc_4_attr_axlock
        ,output [1:0]	int_desc_4_attr_axburst
        ,output [31:0]	int_desc_4_axid_0_axid
        ,output [31:0]	int_desc_4_axid_1_axid
        ,output [31:0]	int_desc_4_axid_2_axid
        ,output [31:0]	int_desc_4_axid_3_axid
        ,output [31:0]	int_desc_4_axuser_0_axuser
        ,output [31:0]	int_desc_4_axuser_1_axuser
        ,output [31:0]	int_desc_4_axuser_2_axuser
        ,output [31:0]	int_desc_4_axuser_3_axuser
        ,output [31:0]	int_desc_4_axuser_4_axuser
        ,output [31:0]	int_desc_4_axuser_5_axuser
        ,output [31:0]	int_desc_4_axuser_6_axuser
        ,output [31:0]	int_desc_4_axuser_7_axuser
        ,output [31:0]	int_desc_4_axuser_8_axuser
        ,output [31:0]	int_desc_4_axuser_9_axuser
        ,output [31:0]	int_desc_4_axuser_10_axuser
        ,output [31:0]	int_desc_4_axuser_11_axuser
        ,output [31:0]	int_desc_4_axuser_12_axuser
        ,output [31:0]	int_desc_4_axuser_13_axuser
        ,output [31:0]	int_desc_4_axuser_14_axuser
        ,output [31:0]	int_desc_4_axuser_15_axuser
        ,output [15:0]	int_desc_4_size_txn_size
        ,output [2:0]	int_desc_4_axsize_axsize
        ,output [31:0]	int_desc_4_axaddr_0_addr
        ,output [31:0]	int_desc_4_axaddr_1_addr
        ,output [31:0]	int_desc_4_axaddr_2_addr
        ,output [31:0]	int_desc_4_axaddr_3_addr
        ,output [31:0]	int_desc_4_data_offset_addr
        ,output [31:0]	int_desc_4_wuser_0_wuser
        ,output [31:0]	int_desc_4_wuser_1_wuser
        ,output [31:0]	int_desc_4_wuser_2_wuser
        ,output [31:0]	int_desc_4_wuser_3_wuser
        ,output [31:0]	int_desc_4_wuser_4_wuser
        ,output [31:0]	int_desc_4_wuser_5_wuser
        ,output [31:0]	int_desc_4_wuser_6_wuser
        ,output [31:0]	int_desc_4_wuser_7_wuser
        ,output [31:0]	int_desc_4_wuser_8_wuser
        ,output [31:0]	int_desc_4_wuser_9_wuser
        ,output [31:0]	int_desc_4_wuser_10_wuser
        ,output [31:0]	int_desc_4_wuser_11_wuser
        ,output [31:0]	int_desc_4_wuser_12_wuser
        ,output [31:0]	int_desc_4_wuser_13_wuser
        ,output [31:0]	int_desc_4_wuser_14_wuser
        ,output [31:0]	int_desc_4_wuser_15_wuser
        ,output [0:0]	int_desc_5_txn_type_wr_strb
        ,output [0:0]	int_desc_5_txn_type_wr_rd
        ,output [3:0]	int_desc_5_attr_axregion
        ,output [3:0]	int_desc_5_attr_axqos
        ,output [2:0]	int_desc_5_attr_axprot
        ,output [3:0]	int_desc_5_attr_axcache
        ,output [1:0]	int_desc_5_attr_axlock
        ,output [1:0]	int_desc_5_attr_axburst
        ,output [31:0]	int_desc_5_axid_0_axid
        ,output [31:0]	int_desc_5_axid_1_axid
        ,output [31:0]	int_desc_5_axid_2_axid
        ,output [31:0]	int_desc_5_axid_3_axid
        ,output [31:0]	int_desc_5_axuser_0_axuser
        ,output [31:0]	int_desc_5_axuser_1_axuser
        ,output [31:0]	int_desc_5_axuser_2_axuser
        ,output [31:0]	int_desc_5_axuser_3_axuser
        ,output [31:0]	int_desc_5_axuser_4_axuser
        ,output [31:0]	int_desc_5_axuser_5_axuser
        ,output [31:0]	int_desc_5_axuser_6_axuser
        ,output [31:0]	int_desc_5_axuser_7_axuser
        ,output [31:0]	int_desc_5_axuser_8_axuser
        ,output [31:0]	int_desc_5_axuser_9_axuser
        ,output [31:0]	int_desc_5_axuser_10_axuser
        ,output [31:0]	int_desc_5_axuser_11_axuser
        ,output [31:0]	int_desc_5_axuser_12_axuser
        ,output [31:0]	int_desc_5_axuser_13_axuser
        ,output [31:0]	int_desc_5_axuser_14_axuser
        ,output [31:0]	int_desc_5_axuser_15_axuser
        ,output [15:0]	int_desc_5_size_txn_size
        ,output [2:0]	int_desc_5_axsize_axsize
        ,output [31:0]	int_desc_5_axaddr_0_addr
        ,output [31:0]	int_desc_5_axaddr_1_addr
        ,output [31:0]	int_desc_5_axaddr_2_addr
        ,output [31:0]	int_desc_5_axaddr_3_addr
        ,output [31:0]	int_desc_5_data_offset_addr
        ,output [31:0]	int_desc_5_wuser_0_wuser
        ,output [31:0]	int_desc_5_wuser_1_wuser
        ,output [31:0]	int_desc_5_wuser_2_wuser
        ,output [31:0]	int_desc_5_wuser_3_wuser
        ,output [31:0]	int_desc_5_wuser_4_wuser
        ,output [31:0]	int_desc_5_wuser_5_wuser
        ,output [31:0]	int_desc_5_wuser_6_wuser
        ,output [31:0]	int_desc_5_wuser_7_wuser
        ,output [31:0]	int_desc_5_wuser_8_wuser
        ,output [31:0]	int_desc_5_wuser_9_wuser
        ,output [31:0]	int_desc_5_wuser_10_wuser
        ,output [31:0]	int_desc_5_wuser_11_wuser
        ,output [31:0]	int_desc_5_wuser_12_wuser
        ,output [31:0]	int_desc_5_wuser_13_wuser
        ,output [31:0]	int_desc_5_wuser_14_wuser
        ,output [31:0]	int_desc_5_wuser_15_wuser
        ,output [0:0]	int_desc_6_txn_type_wr_strb
        ,output [0:0]	int_desc_6_txn_type_wr_rd
        ,output [3:0]	int_desc_6_attr_axregion
        ,output [3:0]	int_desc_6_attr_axqos
        ,output [2:0]	int_desc_6_attr_axprot
        ,output [3:0]	int_desc_6_attr_axcache
        ,output [1:0]	int_desc_6_attr_axlock
        ,output [1:0]	int_desc_6_attr_axburst
        ,output [31:0]	int_desc_6_axid_0_axid
        ,output [31:0]	int_desc_6_axid_1_axid
        ,output [31:0]	int_desc_6_axid_2_axid
        ,output [31:0]	int_desc_6_axid_3_axid
        ,output [31:0]	int_desc_6_axuser_0_axuser
        ,output [31:0]	int_desc_6_axuser_1_axuser
        ,output [31:0]	int_desc_6_axuser_2_axuser
        ,output [31:0]	int_desc_6_axuser_3_axuser
        ,output [31:0]	int_desc_6_axuser_4_axuser
        ,output [31:0]	int_desc_6_axuser_5_axuser
        ,output [31:0]	int_desc_6_axuser_6_axuser
        ,output [31:0]	int_desc_6_axuser_7_axuser
        ,output [31:0]	int_desc_6_axuser_8_axuser
        ,output [31:0]	int_desc_6_axuser_9_axuser
        ,output [31:0]	int_desc_6_axuser_10_axuser
        ,output [31:0]	int_desc_6_axuser_11_axuser
        ,output [31:0]	int_desc_6_axuser_12_axuser
        ,output [31:0]	int_desc_6_axuser_13_axuser
        ,output [31:0]	int_desc_6_axuser_14_axuser
        ,output [31:0]	int_desc_6_axuser_15_axuser
        ,output [15:0]	int_desc_6_size_txn_size
        ,output [2:0]	int_desc_6_axsize_axsize
        ,output [31:0]	int_desc_6_axaddr_0_addr
        ,output [31:0]	int_desc_6_axaddr_1_addr
        ,output [31:0]	int_desc_6_axaddr_2_addr
        ,output [31:0]	int_desc_6_axaddr_3_addr
        ,output [31:0]	int_desc_6_data_offset_addr
        ,output [31:0]	int_desc_6_wuser_0_wuser
        ,output [31:0]	int_desc_6_wuser_1_wuser
        ,output [31:0]	int_desc_6_wuser_2_wuser
        ,output [31:0]	int_desc_6_wuser_3_wuser
        ,output [31:0]	int_desc_6_wuser_4_wuser
        ,output [31:0]	int_desc_6_wuser_5_wuser
        ,output [31:0]	int_desc_6_wuser_6_wuser
        ,output [31:0]	int_desc_6_wuser_7_wuser
        ,output [31:0]	int_desc_6_wuser_8_wuser
        ,output [31:0]	int_desc_6_wuser_9_wuser
        ,output [31:0]	int_desc_6_wuser_10_wuser
        ,output [31:0]	int_desc_6_wuser_11_wuser
        ,output [31:0]	int_desc_6_wuser_12_wuser
        ,output [31:0]	int_desc_6_wuser_13_wuser
        ,output [31:0]	int_desc_6_wuser_14_wuser
        ,output [31:0]	int_desc_6_wuser_15_wuser
        ,output [0:0]	int_desc_7_txn_type_wr_strb
        ,output [0:0]	int_desc_7_txn_type_wr_rd
        ,output [3:0]	int_desc_7_attr_axregion
        ,output [3:0]	int_desc_7_attr_axqos
        ,output [2:0]	int_desc_7_attr_axprot
        ,output [3:0]	int_desc_7_attr_axcache
        ,output [1:0]	int_desc_7_attr_axlock
        ,output [1:0]	int_desc_7_attr_axburst
        ,output [31:0]	int_desc_7_axid_0_axid
        ,output [31:0]	int_desc_7_axid_1_axid
        ,output [31:0]	int_desc_7_axid_2_axid
        ,output [31:0]	int_desc_7_axid_3_axid
        ,output [31:0]	int_desc_7_axuser_0_axuser
        ,output [31:0]	int_desc_7_axuser_1_axuser
        ,output [31:0]	int_desc_7_axuser_2_axuser
        ,output [31:0]	int_desc_7_axuser_3_axuser
        ,output [31:0]	int_desc_7_axuser_4_axuser
        ,output [31:0]	int_desc_7_axuser_5_axuser
        ,output [31:0]	int_desc_7_axuser_6_axuser
        ,output [31:0]	int_desc_7_axuser_7_axuser
        ,output [31:0]	int_desc_7_axuser_8_axuser
        ,output [31:0]	int_desc_7_axuser_9_axuser
        ,output [31:0]	int_desc_7_axuser_10_axuser
        ,output [31:0]	int_desc_7_axuser_11_axuser
        ,output [31:0]	int_desc_7_axuser_12_axuser
        ,output [31:0]	int_desc_7_axuser_13_axuser
        ,output [31:0]	int_desc_7_axuser_14_axuser
        ,output [31:0]	int_desc_7_axuser_15_axuser
        ,output [15:0]	int_desc_7_size_txn_size
        ,output [2:0]	int_desc_7_axsize_axsize
        ,output [31:0]	int_desc_7_axaddr_0_addr
        ,output [31:0]	int_desc_7_axaddr_1_addr
        ,output [31:0]	int_desc_7_axaddr_2_addr
        ,output [31:0]	int_desc_7_axaddr_3_addr
        ,output [31:0]	int_desc_7_data_offset_addr
        ,output [31:0]	int_desc_7_wuser_0_wuser
        ,output [31:0]	int_desc_7_wuser_1_wuser
        ,output [31:0]	int_desc_7_wuser_2_wuser
        ,output [31:0]	int_desc_7_wuser_3_wuser
        ,output [31:0]	int_desc_7_wuser_4_wuser
        ,output [31:0]	int_desc_7_wuser_5_wuser
        ,output [31:0]	int_desc_7_wuser_6_wuser
        ,output [31:0]	int_desc_7_wuser_7_wuser
        ,output [31:0]	int_desc_7_wuser_8_wuser
        ,output [31:0]	int_desc_7_wuser_9_wuser
        ,output [31:0]	int_desc_7_wuser_10_wuser
        ,output [31:0]	int_desc_7_wuser_11_wuser
        ,output [31:0]	int_desc_7_wuser_12_wuser
        ,output [31:0]	int_desc_7_wuser_13_wuser
        ,output [31:0]	int_desc_7_wuser_14_wuser
        ,output [31:0]	int_desc_7_wuser_15_wuser
        ,output [0:0]	int_desc_8_txn_type_wr_strb
        ,output [0:0]	int_desc_8_txn_type_wr_rd
        ,output [3:0]	int_desc_8_attr_axregion
        ,output [3:0]	int_desc_8_attr_axqos
        ,output [2:0]	int_desc_8_attr_axprot
        ,output [3:0]	int_desc_8_attr_axcache
        ,output [1:0]	int_desc_8_attr_axlock
        ,output [1:0]	int_desc_8_attr_axburst
        ,output [31:0]	int_desc_8_axid_0_axid
        ,output [31:0]	int_desc_8_axid_1_axid
        ,output [31:0]	int_desc_8_axid_2_axid
        ,output [31:0]	int_desc_8_axid_3_axid
        ,output [31:0]	int_desc_8_axuser_0_axuser
        ,output [31:0]	int_desc_8_axuser_1_axuser
        ,output [31:0]	int_desc_8_axuser_2_axuser
        ,output [31:0]	int_desc_8_axuser_3_axuser
        ,output [31:0]	int_desc_8_axuser_4_axuser
        ,output [31:0]	int_desc_8_axuser_5_axuser
        ,output [31:0]	int_desc_8_axuser_6_axuser
        ,output [31:0]	int_desc_8_axuser_7_axuser
        ,output [31:0]	int_desc_8_axuser_8_axuser
        ,output [31:0]	int_desc_8_axuser_9_axuser
        ,output [31:0]	int_desc_8_axuser_10_axuser
        ,output [31:0]	int_desc_8_axuser_11_axuser
        ,output [31:0]	int_desc_8_axuser_12_axuser
        ,output [31:0]	int_desc_8_axuser_13_axuser
        ,output [31:0]	int_desc_8_axuser_14_axuser
        ,output [31:0]	int_desc_8_axuser_15_axuser
        ,output [15:0]	int_desc_8_size_txn_size
        ,output [2:0]	int_desc_8_axsize_axsize
        ,output [31:0]	int_desc_8_axaddr_0_addr
        ,output [31:0]	int_desc_8_axaddr_1_addr
        ,output [31:0]	int_desc_8_axaddr_2_addr
        ,output [31:0]	int_desc_8_axaddr_3_addr
        ,output [31:0]	int_desc_8_data_offset_addr
        ,output [31:0]	int_desc_8_wuser_0_wuser
        ,output [31:0]	int_desc_8_wuser_1_wuser
        ,output [31:0]	int_desc_8_wuser_2_wuser
        ,output [31:0]	int_desc_8_wuser_3_wuser
        ,output [31:0]	int_desc_8_wuser_4_wuser
        ,output [31:0]	int_desc_8_wuser_5_wuser
        ,output [31:0]	int_desc_8_wuser_6_wuser
        ,output [31:0]	int_desc_8_wuser_7_wuser
        ,output [31:0]	int_desc_8_wuser_8_wuser
        ,output [31:0]	int_desc_8_wuser_9_wuser
        ,output [31:0]	int_desc_8_wuser_10_wuser
        ,output [31:0]	int_desc_8_wuser_11_wuser
        ,output [31:0]	int_desc_8_wuser_12_wuser
        ,output [31:0]	int_desc_8_wuser_13_wuser
        ,output [31:0]	int_desc_8_wuser_14_wuser
        ,output [31:0]	int_desc_8_wuser_15_wuser
        ,output [0:0]	int_desc_9_txn_type_wr_strb
        ,output [0:0]	int_desc_9_txn_type_wr_rd
        ,output [3:0]	int_desc_9_attr_axregion
        ,output [3:0]	int_desc_9_attr_axqos
        ,output [2:0]	int_desc_9_attr_axprot
        ,output [3:0]	int_desc_9_attr_axcache
        ,output [1:0]	int_desc_9_attr_axlock
        ,output [1:0]	int_desc_9_attr_axburst
        ,output [31:0]	int_desc_9_axid_0_axid
        ,output [31:0]	int_desc_9_axid_1_axid
        ,output [31:0]	int_desc_9_axid_2_axid
        ,output [31:0]	int_desc_9_axid_3_axid
        ,output [31:0]	int_desc_9_axuser_0_axuser
        ,output [31:0]	int_desc_9_axuser_1_axuser
        ,output [31:0]	int_desc_9_axuser_2_axuser
        ,output [31:0]	int_desc_9_axuser_3_axuser
        ,output [31:0]	int_desc_9_axuser_4_axuser
        ,output [31:0]	int_desc_9_axuser_5_axuser
        ,output [31:0]	int_desc_9_axuser_6_axuser
        ,output [31:0]	int_desc_9_axuser_7_axuser
        ,output [31:0]	int_desc_9_axuser_8_axuser
        ,output [31:0]	int_desc_9_axuser_9_axuser
        ,output [31:0]	int_desc_9_axuser_10_axuser
        ,output [31:0]	int_desc_9_axuser_11_axuser
        ,output [31:0]	int_desc_9_axuser_12_axuser
        ,output [31:0]	int_desc_9_axuser_13_axuser
        ,output [31:0]	int_desc_9_axuser_14_axuser
        ,output [31:0]	int_desc_9_axuser_15_axuser
        ,output [15:0]	int_desc_9_size_txn_size
        ,output [2:0]	int_desc_9_axsize_axsize
        ,output [31:0]	int_desc_9_axaddr_0_addr
        ,output [31:0]	int_desc_9_axaddr_1_addr
        ,output [31:0]	int_desc_9_axaddr_2_addr
        ,output [31:0]	int_desc_9_axaddr_3_addr
        ,output [31:0]	int_desc_9_data_offset_addr
        ,output [31:0]	int_desc_9_wuser_0_wuser
        ,output [31:0]	int_desc_9_wuser_1_wuser
        ,output [31:0]	int_desc_9_wuser_2_wuser
        ,output [31:0]	int_desc_9_wuser_3_wuser
        ,output [31:0]	int_desc_9_wuser_4_wuser
        ,output [31:0]	int_desc_9_wuser_5_wuser
        ,output [31:0]	int_desc_9_wuser_6_wuser
        ,output [31:0]	int_desc_9_wuser_7_wuser
        ,output [31:0]	int_desc_9_wuser_8_wuser
        ,output [31:0]	int_desc_9_wuser_9_wuser
        ,output [31:0]	int_desc_9_wuser_10_wuser
        ,output [31:0]	int_desc_9_wuser_11_wuser
        ,output [31:0]	int_desc_9_wuser_12_wuser
        ,output [31:0]	int_desc_9_wuser_13_wuser
        ,output [31:0]	int_desc_9_wuser_14_wuser
        ,output [31:0]	int_desc_9_wuser_15_wuser
        ,output [0:0]	int_desc_10_txn_type_wr_strb
        ,output [0:0]	int_desc_10_txn_type_wr_rd
        ,output [3:0]	int_desc_10_attr_axregion
        ,output [3:0]	int_desc_10_attr_axqos
        ,output [2:0]	int_desc_10_attr_axprot
        ,output [3:0]	int_desc_10_attr_axcache
        ,output [1:0]	int_desc_10_attr_axlock
        ,output [1:0]	int_desc_10_attr_axburst
        ,output [31:0]	int_desc_10_axid_0_axid
        ,output [31:0]	int_desc_10_axid_1_axid
        ,output [31:0]	int_desc_10_axid_2_axid
        ,output [31:0]	int_desc_10_axid_3_axid
        ,output [31:0]	int_desc_10_axuser_0_axuser
        ,output [31:0]	int_desc_10_axuser_1_axuser
        ,output [31:0]	int_desc_10_axuser_2_axuser
        ,output [31:0]	int_desc_10_axuser_3_axuser
        ,output [31:0]	int_desc_10_axuser_4_axuser
        ,output [31:0]	int_desc_10_axuser_5_axuser
        ,output [31:0]	int_desc_10_axuser_6_axuser
        ,output [31:0]	int_desc_10_axuser_7_axuser
        ,output [31:0]	int_desc_10_axuser_8_axuser
        ,output [31:0]	int_desc_10_axuser_9_axuser
        ,output [31:0]	int_desc_10_axuser_10_axuser
        ,output [31:0]	int_desc_10_axuser_11_axuser
        ,output [31:0]	int_desc_10_axuser_12_axuser
        ,output [31:0]	int_desc_10_axuser_13_axuser
        ,output [31:0]	int_desc_10_axuser_14_axuser
        ,output [31:0]	int_desc_10_axuser_15_axuser
        ,output [15:0]	int_desc_10_size_txn_size
        ,output [2:0]	int_desc_10_axsize_axsize
        ,output [31:0]	int_desc_10_axaddr_0_addr
        ,output [31:0]	int_desc_10_axaddr_1_addr
        ,output [31:0]	int_desc_10_axaddr_2_addr
        ,output [31:0]	int_desc_10_axaddr_3_addr
        ,output [31:0]	int_desc_10_data_offset_addr
        ,output [31:0]	int_desc_10_wuser_0_wuser
        ,output [31:0]	int_desc_10_wuser_1_wuser
        ,output [31:0]	int_desc_10_wuser_2_wuser
        ,output [31:0]	int_desc_10_wuser_3_wuser
        ,output [31:0]	int_desc_10_wuser_4_wuser
        ,output [31:0]	int_desc_10_wuser_5_wuser
        ,output [31:0]	int_desc_10_wuser_6_wuser
        ,output [31:0]	int_desc_10_wuser_7_wuser
        ,output [31:0]	int_desc_10_wuser_8_wuser
        ,output [31:0]	int_desc_10_wuser_9_wuser
        ,output [31:0]	int_desc_10_wuser_10_wuser
        ,output [31:0]	int_desc_10_wuser_11_wuser
        ,output [31:0]	int_desc_10_wuser_12_wuser
        ,output [31:0]	int_desc_10_wuser_13_wuser
        ,output [31:0]	int_desc_10_wuser_14_wuser
        ,output [31:0]	int_desc_10_wuser_15_wuser
        ,output [0:0]	int_desc_11_txn_type_wr_strb
        ,output [0:0]	int_desc_11_txn_type_wr_rd
        ,output [3:0]	int_desc_11_attr_axregion
        ,output [3:0]	int_desc_11_attr_axqos
        ,output [2:0]	int_desc_11_attr_axprot
        ,output [3:0]	int_desc_11_attr_axcache
        ,output [1:0]	int_desc_11_attr_axlock
        ,output [1:0]	int_desc_11_attr_axburst
        ,output [31:0]	int_desc_11_axid_0_axid
        ,output [31:0]	int_desc_11_axid_1_axid
        ,output [31:0]	int_desc_11_axid_2_axid
        ,output [31:0]	int_desc_11_axid_3_axid
        ,output [31:0]	int_desc_11_axuser_0_axuser
        ,output [31:0]	int_desc_11_axuser_1_axuser
        ,output [31:0]	int_desc_11_axuser_2_axuser
        ,output [31:0]	int_desc_11_axuser_3_axuser
        ,output [31:0]	int_desc_11_axuser_4_axuser
        ,output [31:0]	int_desc_11_axuser_5_axuser
        ,output [31:0]	int_desc_11_axuser_6_axuser
        ,output [31:0]	int_desc_11_axuser_7_axuser
        ,output [31:0]	int_desc_11_axuser_8_axuser
        ,output [31:0]	int_desc_11_axuser_9_axuser
        ,output [31:0]	int_desc_11_axuser_10_axuser
        ,output [31:0]	int_desc_11_axuser_11_axuser
        ,output [31:0]	int_desc_11_axuser_12_axuser
        ,output [31:0]	int_desc_11_axuser_13_axuser
        ,output [31:0]	int_desc_11_axuser_14_axuser
        ,output [31:0]	int_desc_11_axuser_15_axuser
        ,output [15:0]	int_desc_11_size_txn_size
        ,output [2:0]	int_desc_11_axsize_axsize
        ,output [31:0]	int_desc_11_axaddr_0_addr
        ,output [31:0]	int_desc_11_axaddr_1_addr
        ,output [31:0]	int_desc_11_axaddr_2_addr
        ,output [31:0]	int_desc_11_axaddr_3_addr
        ,output [31:0]	int_desc_11_data_offset_addr
        ,output [31:0]	int_desc_11_wuser_0_wuser
        ,output [31:0]	int_desc_11_wuser_1_wuser
        ,output [31:0]	int_desc_11_wuser_2_wuser
        ,output [31:0]	int_desc_11_wuser_3_wuser
        ,output [31:0]	int_desc_11_wuser_4_wuser
        ,output [31:0]	int_desc_11_wuser_5_wuser
        ,output [31:0]	int_desc_11_wuser_6_wuser
        ,output [31:0]	int_desc_11_wuser_7_wuser
        ,output [31:0]	int_desc_11_wuser_8_wuser
        ,output [31:0]	int_desc_11_wuser_9_wuser
        ,output [31:0]	int_desc_11_wuser_10_wuser
        ,output [31:0]	int_desc_11_wuser_11_wuser
        ,output [31:0]	int_desc_11_wuser_12_wuser
        ,output [31:0]	int_desc_11_wuser_13_wuser
        ,output [31:0]	int_desc_11_wuser_14_wuser
        ,output [31:0]	int_desc_11_wuser_15_wuser
        ,output [0:0]	int_desc_12_txn_type_wr_strb
        ,output [0:0]	int_desc_12_txn_type_wr_rd
        ,output [3:0]	int_desc_12_attr_axregion
        ,output [3:0]	int_desc_12_attr_axqos
        ,output [2:0]	int_desc_12_attr_axprot
        ,output [3:0]	int_desc_12_attr_axcache
        ,output [1:0]	int_desc_12_attr_axlock
        ,output [1:0]	int_desc_12_attr_axburst
        ,output [31:0]	int_desc_12_axid_0_axid
        ,output [31:0]	int_desc_12_axid_1_axid
        ,output [31:0]	int_desc_12_axid_2_axid
        ,output [31:0]	int_desc_12_axid_3_axid
        ,output [31:0]	int_desc_12_axuser_0_axuser
        ,output [31:0]	int_desc_12_axuser_1_axuser
        ,output [31:0]	int_desc_12_axuser_2_axuser
        ,output [31:0]	int_desc_12_axuser_3_axuser
        ,output [31:0]	int_desc_12_axuser_4_axuser
        ,output [31:0]	int_desc_12_axuser_5_axuser
        ,output [31:0]	int_desc_12_axuser_6_axuser
        ,output [31:0]	int_desc_12_axuser_7_axuser
        ,output [31:0]	int_desc_12_axuser_8_axuser
        ,output [31:0]	int_desc_12_axuser_9_axuser
        ,output [31:0]	int_desc_12_axuser_10_axuser
        ,output [31:0]	int_desc_12_axuser_11_axuser
        ,output [31:0]	int_desc_12_axuser_12_axuser
        ,output [31:0]	int_desc_12_axuser_13_axuser
        ,output [31:0]	int_desc_12_axuser_14_axuser
        ,output [31:0]	int_desc_12_axuser_15_axuser
        ,output [15:0]	int_desc_12_size_txn_size
        ,output [2:0]	int_desc_12_axsize_axsize
        ,output [31:0]	int_desc_12_axaddr_0_addr
        ,output [31:0]	int_desc_12_axaddr_1_addr
        ,output [31:0]	int_desc_12_axaddr_2_addr
        ,output [31:0]	int_desc_12_axaddr_3_addr
        ,output [31:0]	int_desc_12_data_offset_addr
        ,output [31:0]	int_desc_12_wuser_0_wuser
        ,output [31:0]	int_desc_12_wuser_1_wuser
        ,output [31:0]	int_desc_12_wuser_2_wuser
        ,output [31:0]	int_desc_12_wuser_3_wuser
        ,output [31:0]	int_desc_12_wuser_4_wuser
        ,output [31:0]	int_desc_12_wuser_5_wuser
        ,output [31:0]	int_desc_12_wuser_6_wuser
        ,output [31:0]	int_desc_12_wuser_7_wuser
        ,output [31:0]	int_desc_12_wuser_8_wuser
        ,output [31:0]	int_desc_12_wuser_9_wuser
        ,output [31:0]	int_desc_12_wuser_10_wuser
        ,output [31:0]	int_desc_12_wuser_11_wuser
        ,output [31:0]	int_desc_12_wuser_12_wuser
        ,output [31:0]	int_desc_12_wuser_13_wuser
        ,output [31:0]	int_desc_12_wuser_14_wuser
        ,output [31:0]	int_desc_12_wuser_15_wuser
        ,output [0:0]	int_desc_13_txn_type_wr_strb
        ,output [0:0]	int_desc_13_txn_type_wr_rd
        ,output [3:0]	int_desc_13_attr_axregion
        ,output [3:0]	int_desc_13_attr_axqos
        ,output [2:0]	int_desc_13_attr_axprot
        ,output [3:0]	int_desc_13_attr_axcache
        ,output [1:0]	int_desc_13_attr_axlock
        ,output [1:0]	int_desc_13_attr_axburst
        ,output [31:0]	int_desc_13_axid_0_axid
        ,output [31:0]	int_desc_13_axid_1_axid
        ,output [31:0]	int_desc_13_axid_2_axid
        ,output [31:0]	int_desc_13_axid_3_axid
        ,output [31:0]	int_desc_13_axuser_0_axuser
        ,output [31:0]	int_desc_13_axuser_1_axuser
        ,output [31:0]	int_desc_13_axuser_2_axuser
        ,output [31:0]	int_desc_13_axuser_3_axuser
        ,output [31:0]	int_desc_13_axuser_4_axuser
        ,output [31:0]	int_desc_13_axuser_5_axuser
        ,output [31:0]	int_desc_13_axuser_6_axuser
        ,output [31:0]	int_desc_13_axuser_7_axuser
        ,output [31:0]	int_desc_13_axuser_8_axuser
        ,output [31:0]	int_desc_13_axuser_9_axuser
        ,output [31:0]	int_desc_13_axuser_10_axuser
        ,output [31:0]	int_desc_13_axuser_11_axuser
        ,output [31:0]	int_desc_13_axuser_12_axuser
        ,output [31:0]	int_desc_13_axuser_13_axuser
        ,output [31:0]	int_desc_13_axuser_14_axuser
        ,output [31:0]	int_desc_13_axuser_15_axuser
        ,output [15:0]	int_desc_13_size_txn_size
        ,output [2:0]	int_desc_13_axsize_axsize
        ,output [31:0]	int_desc_13_axaddr_0_addr
        ,output [31:0]	int_desc_13_axaddr_1_addr
        ,output [31:0]	int_desc_13_axaddr_2_addr
        ,output [31:0]	int_desc_13_axaddr_3_addr
        ,output [31:0]	int_desc_13_data_offset_addr
        ,output [31:0]	int_desc_13_wuser_0_wuser
        ,output [31:0]	int_desc_13_wuser_1_wuser
        ,output [31:0]	int_desc_13_wuser_2_wuser
        ,output [31:0]	int_desc_13_wuser_3_wuser
        ,output [31:0]	int_desc_13_wuser_4_wuser
        ,output [31:0]	int_desc_13_wuser_5_wuser
        ,output [31:0]	int_desc_13_wuser_6_wuser
        ,output [31:0]	int_desc_13_wuser_7_wuser
        ,output [31:0]	int_desc_13_wuser_8_wuser
        ,output [31:0]	int_desc_13_wuser_9_wuser
        ,output [31:0]	int_desc_13_wuser_10_wuser
        ,output [31:0]	int_desc_13_wuser_11_wuser
        ,output [31:0]	int_desc_13_wuser_12_wuser
        ,output [31:0]	int_desc_13_wuser_13_wuser
        ,output [31:0]	int_desc_13_wuser_14_wuser
        ,output [31:0]	int_desc_13_wuser_15_wuser
        ,output [0:0]	int_desc_14_txn_type_wr_strb
        ,output [0:0]	int_desc_14_txn_type_wr_rd
        ,output [3:0]	int_desc_14_attr_axregion
        ,output [3:0]	int_desc_14_attr_axqos
        ,output [2:0]	int_desc_14_attr_axprot
        ,output [3:0]	int_desc_14_attr_axcache
        ,output [1:0]	int_desc_14_attr_axlock
        ,output [1:0]	int_desc_14_attr_axburst
        ,output [31:0]	int_desc_14_axid_0_axid
        ,output [31:0]	int_desc_14_axid_1_axid
        ,output [31:0]	int_desc_14_axid_2_axid
        ,output [31:0]	int_desc_14_axid_3_axid
        ,output [31:0]	int_desc_14_axuser_0_axuser
        ,output [31:0]	int_desc_14_axuser_1_axuser
        ,output [31:0]	int_desc_14_axuser_2_axuser
        ,output [31:0]	int_desc_14_axuser_3_axuser
        ,output [31:0]	int_desc_14_axuser_4_axuser
        ,output [31:0]	int_desc_14_axuser_5_axuser
        ,output [31:0]	int_desc_14_axuser_6_axuser
        ,output [31:0]	int_desc_14_axuser_7_axuser
        ,output [31:0]	int_desc_14_axuser_8_axuser
        ,output [31:0]	int_desc_14_axuser_9_axuser
        ,output [31:0]	int_desc_14_axuser_10_axuser
        ,output [31:0]	int_desc_14_axuser_11_axuser
        ,output [31:0]	int_desc_14_axuser_12_axuser
        ,output [31:0]	int_desc_14_axuser_13_axuser
        ,output [31:0]	int_desc_14_axuser_14_axuser
        ,output [31:0]	int_desc_14_axuser_15_axuser
        ,output [15:0]	int_desc_14_size_txn_size
        ,output [2:0]	int_desc_14_axsize_axsize
        ,output [31:0]	int_desc_14_axaddr_0_addr
        ,output [31:0]	int_desc_14_axaddr_1_addr
        ,output [31:0]	int_desc_14_axaddr_2_addr
        ,output [31:0]	int_desc_14_axaddr_3_addr
        ,output [31:0]	int_desc_14_data_offset_addr
        ,output [31:0]	int_desc_14_wuser_0_wuser
        ,output [31:0]	int_desc_14_wuser_1_wuser
        ,output [31:0]	int_desc_14_wuser_2_wuser
        ,output [31:0]	int_desc_14_wuser_3_wuser
        ,output [31:0]	int_desc_14_wuser_4_wuser
        ,output [31:0]	int_desc_14_wuser_5_wuser
        ,output [31:0]	int_desc_14_wuser_6_wuser
        ,output [31:0]	int_desc_14_wuser_7_wuser
        ,output [31:0]	int_desc_14_wuser_8_wuser
        ,output [31:0]	int_desc_14_wuser_9_wuser
        ,output [31:0]	int_desc_14_wuser_10_wuser
        ,output [31:0]	int_desc_14_wuser_11_wuser
        ,output [31:0]	int_desc_14_wuser_12_wuser
        ,output [31:0]	int_desc_14_wuser_13_wuser
        ,output [31:0]	int_desc_14_wuser_14_wuser
        ,output [31:0]	int_desc_14_wuser_15_wuser
        ,output [0:0]	int_desc_15_txn_type_wr_strb
        ,output [0:0]	int_desc_15_txn_type_wr_rd
        ,output [3:0]	int_desc_15_attr_axregion
        ,output [3:0]	int_desc_15_attr_axqos
        ,output [2:0]	int_desc_15_attr_axprot
        ,output [3:0]	int_desc_15_attr_axcache
        ,output [1:0]	int_desc_15_attr_axlock
        ,output [1:0]	int_desc_15_attr_axburst
        ,output [31:0]	int_desc_15_axid_0_axid
        ,output [31:0]	int_desc_15_axid_1_axid
        ,output [31:0]	int_desc_15_axid_2_axid
        ,output [31:0]	int_desc_15_axid_3_axid
        ,output [31:0]	int_desc_15_axuser_0_axuser
        ,output [31:0]	int_desc_15_axuser_1_axuser
        ,output [31:0]	int_desc_15_axuser_2_axuser
        ,output [31:0]	int_desc_15_axuser_3_axuser
        ,output [31:0]	int_desc_15_axuser_4_axuser
        ,output [31:0]	int_desc_15_axuser_5_axuser
        ,output [31:0]	int_desc_15_axuser_6_axuser
        ,output [31:0]	int_desc_15_axuser_7_axuser
        ,output [31:0]	int_desc_15_axuser_8_axuser
        ,output [31:0]	int_desc_15_axuser_9_axuser
        ,output [31:0]	int_desc_15_axuser_10_axuser
        ,output [31:0]	int_desc_15_axuser_11_axuser
        ,output [31:0]	int_desc_15_axuser_12_axuser
        ,output [31:0]	int_desc_15_axuser_13_axuser
        ,output [31:0]	int_desc_15_axuser_14_axuser
        ,output [31:0]	int_desc_15_axuser_15_axuser
        ,output [15:0]	int_desc_15_size_txn_size
        ,output [2:0]	int_desc_15_axsize_axsize
        ,output [31:0]	int_desc_15_axaddr_0_addr
        ,output [31:0]	int_desc_15_axaddr_1_addr
        ,output [31:0]	int_desc_15_axaddr_2_addr
        ,output [31:0]	int_desc_15_axaddr_3_addr
        ,output [31:0]	int_desc_15_data_offset_addr
        ,output [31:0]	int_desc_15_wuser_0_wuser
        ,output [31:0]	int_desc_15_wuser_1_wuser
        ,output [31:0]	int_desc_15_wuser_2_wuser
        ,output [31:0]	int_desc_15_wuser_3_wuser
        ,output [31:0]	int_desc_15_wuser_4_wuser
        ,output [31:0]	int_desc_15_wuser_5_wuser
        ,output [31:0]	int_desc_15_wuser_6_wuser
        ,output [31:0]	int_desc_15_wuser_7_wuser
        ,output [31:0]	int_desc_15_wuser_8_wuser
        ,output [31:0]	int_desc_15_wuser_9_wuser
        ,output [31:0]	int_desc_15_wuser_10_wuser
        ,output [31:0]	int_desc_15_wuser_11_wuser
        ,output [31:0]	int_desc_15_wuser_12_wuser
        ,output [31:0]	int_desc_15_wuser_13_wuser
        ,output [31:0]	int_desc_15_wuser_14_wuser
        ,output [31:0]	int_desc_15_wuser_15_wuser
