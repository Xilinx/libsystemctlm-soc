/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *   This module is replica of ace_usr_slv_control module but it converts
 *   all registers into the internal fields as int_<reg>_<field> . Only these fields 
 *   are used in further hierarchy rather than registers.
 *
 *
 */

`include "ace_defines_common.vh"

module ace_usr_slv_control_field #(

				    parameter ACE_PROTOCOL                   = "FULLACE" 
				    
				    ,parameter ADDR_WIDTH                     = 64 
				    ,parameter XX_DATA_WIDTH                  = 128       
				    ,parameter SN_DATA_WIDTH                  = 128       
				    ,parameter ID_WIDTH                       = 16 
				    ,parameter AWUSER_WIDTH                   = 32 
				    ,parameter WUSER_WIDTH                    = 32 
				    ,parameter BUSER_WIDTH                    = 32 
				    ,parameter ARUSER_WIDTH                   = 32 
				    ,parameter RUSER_WIDTH                    = 32 
				    
				    ,parameter CACHE_LINE_SIZE                = 64 
				    ,parameter XX_MAX_DESC                    = 16         
				    ,parameter SN_MAX_DESC                    = 16         
				    ,parameter XX_RAM_SIZE                    = 16384     
				    ,parameter SN_RAM_SIZE                    = 512       

				    )(

				      //Clock and reset
				      input clk 
				      ,input resetn
   
				      //S_ACE_USR
				      ,input [ID_WIDTH-1:0] s_ace_usr_awid 
				      ,input [ADDR_WIDTH-1:0] s_ace_usr_awaddr 
				      ,input [7:0] s_ace_usr_awlen
				      ,input [2:0] s_ace_usr_awsize 
				      ,input [1:0] s_ace_usr_awburst 
				      ,input s_ace_usr_awlock 
				      ,input [3:0] s_ace_usr_awcache 
				      ,input [2:0] s_ace_usr_awprot 
				      ,input [3:0] s_ace_usr_awqos 
				      ,input [3:0] s_ace_usr_awregion 
				      ,input [AWUSER_WIDTH-1:0] s_ace_usr_awuser 
				      ,input [2:0] s_ace_usr_awsnoop 
				      ,input [1:0] s_ace_usr_awdomain 
				      ,input [1:0] s_ace_usr_awbar 
				      ,input s_ace_usr_awunique 
				      ,input s_ace_usr_awvalid 
				      ,output s_ace_usr_awready 
				      ,input [XX_DATA_WIDTH-1:0] s_ace_usr_wdata 
				      ,input [(XX_DATA_WIDTH/8)-1:0] s_ace_usr_wstrb
				      ,input s_ace_usr_wlast 
				      ,input [WUSER_WIDTH-1:0] s_ace_usr_wuser 
				      ,input s_ace_usr_wvalid 
				      ,output s_ace_usr_wready 
				      ,output [ID_WIDTH-1:0] s_ace_usr_bid 
				      ,output [1:0] s_ace_usr_bresp 
				      ,output [BUSER_WIDTH-1:0] s_ace_usr_buser 
				      ,output s_ace_usr_bvalid 
				      ,input s_ace_usr_bready 
				      ,input s_ace_usr_wack 
				      ,input [ID_WIDTH-1:0] s_ace_usr_arid 
				      ,input [ADDR_WIDTH-1:0] s_ace_usr_araddr 
				      ,input [7:0] s_ace_usr_arlen 
				      ,input [2:0] s_ace_usr_arsize 
				      ,input [1:0] s_ace_usr_arburst 
				      ,input s_ace_usr_arlock 
				      ,input [3:0] s_ace_usr_arcache 
				      ,input [2:0] s_ace_usr_arprot 
				      ,input [3:0] s_ace_usr_arqos 
				      ,input [3:0] s_ace_usr_arregion 
				      ,input [ARUSER_WIDTH-1:0] s_ace_usr_aruser 
				      ,input [3:0] s_ace_usr_arsnoop 
				      ,input [1:0] s_ace_usr_ardomain 
				      ,input [1:0] s_ace_usr_arbar 
				      ,input s_ace_usr_arvalid 
				      ,output s_ace_usr_arready 
				      ,output [ID_WIDTH-1:0] s_ace_usr_rid 
				      ,output [XX_DATA_WIDTH-1:0] s_ace_usr_rdata 
				      ,output [3:0] s_ace_usr_rresp 
				      ,output s_ace_usr_rlast 
				      ,output [RUSER_WIDTH-1:0] s_ace_usr_ruser 
				      ,output s_ace_usr_rvalid 
				      ,input s_ace_usr_rready 
				      ,input s_ace_usr_rack 
				      ,output [ADDR_WIDTH-1:0] s_ace_usr_acaddr 
				      ,output [3:0] s_ace_usr_acsnoop 
				      ,output [2:0] s_ace_usr_acprot 
				      ,output s_ace_usr_acvalid 
				      ,input s_ace_usr_acready 
				      ,input [4:0] s_ace_usr_crresp 
				      ,input s_ace_usr_crvalid 
				      ,output s_ace_usr_crready 
				      ,input [SN_DATA_WIDTH-1:0] s_ace_usr_cddata 
				      ,input s_ace_usr_cdlast 
				      ,input s_ace_usr_cdvalid 
				      ,output s_ace_usr_cdready 
   
				      ,input [31:0] bridge_identification_reg
				      ,input [31:0] last_bridge_reg
				      ,input [31:0] version_reg
				      ,input [31:0] bridge_type_reg
				      ,input [31:0] mode_select_reg
				      ,input [31:0] reset_reg
				      ,input [31:0] h2c_intr_0_reg
				      ,input [31:0] h2c_intr_1_reg
				      ,input [31:0] h2c_intr_2_reg
				      ,input [31:0] h2c_intr_3_reg
				      ,input [31:0] c2h_intr_status_0_reg
				      ,input [31:0] intr_c2h_toggle_status_0_reg
				      ,input [31:0] intr_c2h_toggle_clear_0_reg
				      ,input [31:0] intr_c2h_toggle_enable_0_reg
				      ,input [31:0] c2h_intr_status_1_reg
				      ,input [31:0] intr_c2h_toggle_status_1_reg
				      ,input [31:0] intr_c2h_toggle_clear_1_reg
				      ,input [31:0] intr_c2h_toggle_enable_1_reg
				      ,input [31:0] c2h_gpio_0_reg
				      ,input [31:0] c2h_gpio_1_reg
				      ,input [31:0] c2h_gpio_2_reg
				      ,input [31:0] c2h_gpio_3_reg
				      ,input [31:0] c2h_gpio_4_reg
				      ,input [31:0] c2h_gpio_5_reg
				      ,input [31:0] c2h_gpio_6_reg
				      ,input [31:0] c2h_gpio_7_reg
				      ,input [31:0] c2h_gpio_8_reg
				      ,input [31:0] c2h_gpio_9_reg
				      ,input [31:0] c2h_gpio_10_reg
				      ,input [31:0] c2h_gpio_11_reg
				      ,input [31:0] c2h_gpio_12_reg
				      ,input [31:0] c2h_gpio_13_reg
				      ,input [31:0] c2h_gpio_14_reg
				      ,input [31:0] c2h_gpio_15_reg
				      ,input [31:0] h2c_gpio_0_reg
				      ,input [31:0] h2c_gpio_1_reg
				      ,input [31:0] h2c_gpio_2_reg
				      ,input [31:0] h2c_gpio_3_reg
				      ,input [31:0] h2c_gpio_4_reg
				      ,input [31:0] h2c_gpio_5_reg
				      ,input [31:0] h2c_gpio_6_reg
				      ,input [31:0] h2c_gpio_7_reg
				      ,input [31:0] h2c_gpio_8_reg
				      ,input [31:0] h2c_gpio_9_reg
				      ,input [31:0] h2c_gpio_10_reg
				      ,input [31:0] h2c_gpio_11_reg
				      ,input [31:0] h2c_gpio_12_reg
				      ,input [31:0] h2c_gpio_13_reg
				      ,input [31:0] h2c_gpio_14_reg
				      ,input [31:0] h2c_gpio_15_reg
				      ,input [31:0] bridge_config_reg
				      ,input [31:0] intr_status_reg
				      ,input [31:0] intr_error_status_reg
				      ,input [31:0] intr_error_clear_reg
				      ,input [31:0] intr_error_enable_reg
				      ,input [31:0] bridge_rd_user_config_reg
				      ,input [31:0] bridge_wr_user_config_reg
				      ,input [31:0] rd_max_desc_reg
				      ,input [31:0] wr_max_desc_reg
				      ,input [31:0] sn_max_desc_reg
				      ,input [31:0] rd_req_free_desc_reg
				      ,input [31:0] rd_req_fifo_pop_desc_reg
				      ,input [31:0] rd_req_fifo_fill_level_reg
				      ,input [31:0] rd_resp_fifo_push_desc_reg
				      ,input [31:0] rd_resp_fifo_free_level_reg
				      ,input [31:0] rd_resp_intr_comp_status_reg
				      ,input [31:0] rd_resp_intr_comp_clear_reg
				      ,input [31:0] rd_resp_intr_comp_enable_reg
				      ,input [31:0] wr_req_free_desc_reg
				      ,input [31:0] wr_req_fifo_pop_desc_reg
				      ,input [31:0] wr_req_fifo_fill_level_reg
				      ,input [31:0] wr_resp_fifo_push_desc_reg
				      ,input [31:0] wr_resp_fifo_free_level_reg
				      ,input [31:0] wr_resp_intr_comp_status_reg
				      ,input [31:0] wr_resp_intr_comp_clear_reg
				      ,input [31:0] wr_resp_intr_comp_enable_reg
				      ,input [31:0] sn_req_fifo_push_desc_reg
				      ,input [31:0] sn_req_fifo_free_level_reg
				      ,input [31:0] sn_req_intr_comp_status_reg
				      ,input [31:0] sn_req_intr_comp_clear_reg
				      ,input [31:0] sn_req_intr_comp_enable_reg
				      ,input [31:0] sn_resp_free_desc_reg
				      ,input [31:0] sn_resp_fifo_pop_desc_reg
				      ,input [31:0] sn_resp_fifo_fill_level_reg
				      ,input [31:0] sn_data_free_desc_reg
				      ,input [31:0] sn_data_fifo_pop_desc_reg
				      ,input [31:0] sn_data_fifo_fill_level_reg
				      ,input [31:0] intr_fifo_enable_reg
				      ,input [31:0] rd_req_desc_0_txn_type_reg
				      ,input [31:0] rd_req_desc_0_size_reg
				      ,input [31:0] rd_req_desc_0_axsize_reg
				      ,input [31:0] rd_req_desc_0_attr_reg
				      ,input [31:0] rd_req_desc_0_axaddr_0_reg
				      ,input [31:0] rd_req_desc_0_axaddr_1_reg
				      ,input [31:0] rd_req_desc_0_axaddr_2_reg
				      ,input [31:0] rd_req_desc_0_axaddr_3_reg
				      ,input [31:0] rd_req_desc_0_axid_0_reg
				      ,input [31:0] rd_req_desc_0_axid_1_reg
				      ,input [31:0] rd_req_desc_0_axid_2_reg
				      ,input [31:0] rd_req_desc_0_axid_3_reg
				      ,input [31:0] rd_req_desc_0_axuser_0_reg
				      ,input [31:0] rd_req_desc_0_axuser_1_reg
				      ,input [31:0] rd_req_desc_0_axuser_2_reg
				      ,input [31:0] rd_req_desc_0_axuser_3_reg
				      ,input [31:0] rd_req_desc_0_axuser_4_reg
				      ,input [31:0] rd_req_desc_0_axuser_5_reg
				      ,input [31:0] rd_req_desc_0_axuser_6_reg
				      ,input [31:0] rd_req_desc_0_axuser_7_reg
				      ,input [31:0] rd_req_desc_0_axuser_8_reg
				      ,input [31:0] rd_req_desc_0_axuser_9_reg
				      ,input [31:0] rd_req_desc_0_axuser_10_reg
				      ,input [31:0] rd_req_desc_0_axuser_11_reg
				      ,input [31:0] rd_req_desc_0_axuser_12_reg
				      ,input [31:0] rd_req_desc_0_axuser_13_reg
				      ,input [31:0] rd_req_desc_0_axuser_14_reg
				      ,input [31:0] rd_req_desc_0_axuser_15_reg
				      ,input [31:0] rd_resp_desc_0_data_offset_reg
				      ,input [31:0] rd_resp_desc_0_data_size_reg
				      ,input [31:0] rd_resp_desc_0_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_0_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_0_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_0_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_0_resp_reg
				      ,input [31:0] rd_resp_desc_0_xid_0_reg
				      ,input [31:0] rd_resp_desc_0_xid_1_reg
				      ,input [31:0] rd_resp_desc_0_xid_2_reg
				      ,input [31:0] rd_resp_desc_0_xid_3_reg
				      ,input [31:0] rd_resp_desc_0_xuser_0_reg
				      ,input [31:0] rd_resp_desc_0_xuser_1_reg
				      ,input [31:0] rd_resp_desc_0_xuser_2_reg
				      ,input [31:0] rd_resp_desc_0_xuser_3_reg
				      ,input [31:0] rd_resp_desc_0_xuser_4_reg
				      ,input [31:0] rd_resp_desc_0_xuser_5_reg
				      ,input [31:0] rd_resp_desc_0_xuser_6_reg
				      ,input [31:0] rd_resp_desc_0_xuser_7_reg
				      ,input [31:0] rd_resp_desc_0_xuser_8_reg
				      ,input [31:0] rd_resp_desc_0_xuser_9_reg
				      ,input [31:0] rd_resp_desc_0_xuser_10_reg
				      ,input [31:0] rd_resp_desc_0_xuser_11_reg
				      ,input [31:0] rd_resp_desc_0_xuser_12_reg
				      ,input [31:0] rd_resp_desc_0_xuser_13_reg
				      ,input [31:0] rd_resp_desc_0_xuser_14_reg
				      ,input [31:0] rd_resp_desc_0_xuser_15_reg
				      ,input [31:0] wr_req_desc_0_txn_type_reg
				      ,input [31:0] wr_req_desc_0_size_reg
				      ,input [31:0] wr_req_desc_0_data_offset_reg
				      ,input [31:0] wr_req_desc_0_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_0_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_0_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_0_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_0_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_0_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_0_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_0_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_0_axsize_reg
				      ,input [31:0] wr_req_desc_0_attr_reg
				      ,input [31:0] wr_req_desc_0_axaddr_0_reg
				      ,input [31:0] wr_req_desc_0_axaddr_1_reg
				      ,input [31:0] wr_req_desc_0_axaddr_2_reg
				      ,input [31:0] wr_req_desc_0_axaddr_3_reg
				      ,input [31:0] wr_req_desc_0_axid_0_reg
				      ,input [31:0] wr_req_desc_0_axid_1_reg
				      ,input [31:0] wr_req_desc_0_axid_2_reg
				      ,input [31:0] wr_req_desc_0_axid_3_reg
				      ,input [31:0] wr_req_desc_0_axuser_0_reg
				      ,input [31:0] wr_req_desc_0_axuser_1_reg
				      ,input [31:0] wr_req_desc_0_axuser_2_reg
				      ,input [31:0] wr_req_desc_0_axuser_3_reg
				      ,input [31:0] wr_req_desc_0_axuser_4_reg
				      ,input [31:0] wr_req_desc_0_axuser_5_reg
				      ,input [31:0] wr_req_desc_0_axuser_6_reg
				      ,input [31:0] wr_req_desc_0_axuser_7_reg
				      ,input [31:0] wr_req_desc_0_axuser_8_reg
				      ,input [31:0] wr_req_desc_0_axuser_9_reg
				      ,input [31:0] wr_req_desc_0_axuser_10_reg
				      ,input [31:0] wr_req_desc_0_axuser_11_reg
				      ,input [31:0] wr_req_desc_0_axuser_12_reg
				      ,input [31:0] wr_req_desc_0_axuser_13_reg
				      ,input [31:0] wr_req_desc_0_axuser_14_reg
				      ,input [31:0] wr_req_desc_0_axuser_15_reg
				      ,input [31:0] wr_req_desc_0_wuser_0_reg
				      ,input [31:0] wr_req_desc_0_wuser_1_reg
				      ,input [31:0] wr_req_desc_0_wuser_2_reg
				      ,input [31:0] wr_req_desc_0_wuser_3_reg
				      ,input [31:0] wr_req_desc_0_wuser_4_reg
				      ,input [31:0] wr_req_desc_0_wuser_5_reg
				      ,input [31:0] wr_req_desc_0_wuser_6_reg
				      ,input [31:0] wr_req_desc_0_wuser_7_reg
				      ,input [31:0] wr_req_desc_0_wuser_8_reg
				      ,input [31:0] wr_req_desc_0_wuser_9_reg
				      ,input [31:0] wr_req_desc_0_wuser_10_reg
				      ,input [31:0] wr_req_desc_0_wuser_11_reg
				      ,input [31:0] wr_req_desc_0_wuser_12_reg
				      ,input [31:0] wr_req_desc_0_wuser_13_reg
				      ,input [31:0] wr_req_desc_0_wuser_14_reg
				      ,input [31:0] wr_req_desc_0_wuser_15_reg
				      ,input [31:0] wr_resp_desc_0_resp_reg
				      ,input [31:0] wr_resp_desc_0_xid_0_reg
				      ,input [31:0] wr_resp_desc_0_xid_1_reg
				      ,input [31:0] wr_resp_desc_0_xid_2_reg
				      ,input [31:0] wr_resp_desc_0_xid_3_reg
				      ,input [31:0] wr_resp_desc_0_xuser_0_reg
				      ,input [31:0] wr_resp_desc_0_xuser_1_reg
				      ,input [31:0] wr_resp_desc_0_xuser_2_reg
				      ,input [31:0] wr_resp_desc_0_xuser_3_reg
				      ,input [31:0] wr_resp_desc_0_xuser_4_reg
				      ,input [31:0] wr_resp_desc_0_xuser_5_reg
				      ,input [31:0] wr_resp_desc_0_xuser_6_reg
				      ,input [31:0] wr_resp_desc_0_xuser_7_reg
				      ,input [31:0] wr_resp_desc_0_xuser_8_reg
				      ,input [31:0] wr_resp_desc_0_xuser_9_reg
				      ,input [31:0] wr_resp_desc_0_xuser_10_reg
				      ,input [31:0] wr_resp_desc_0_xuser_11_reg
				      ,input [31:0] wr_resp_desc_0_xuser_12_reg
				      ,input [31:0] wr_resp_desc_0_xuser_13_reg
				      ,input [31:0] wr_resp_desc_0_xuser_14_reg
				      ,input [31:0] wr_resp_desc_0_xuser_15_reg
				      ,input [31:0] sn_req_desc_0_attr_reg
				      ,input [31:0] sn_req_desc_0_acaddr_0_reg
				      ,input [31:0] sn_req_desc_0_acaddr_1_reg
				      ,input [31:0] sn_req_desc_0_acaddr_2_reg
				      ,input [31:0] sn_req_desc_0_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_0_resp_reg
				      ,input [31:0] rd_req_desc_1_txn_type_reg
				      ,input [31:0] rd_req_desc_1_size_reg
				      ,input [31:0] rd_req_desc_1_axsize_reg
				      ,input [31:0] rd_req_desc_1_attr_reg
				      ,input [31:0] rd_req_desc_1_axaddr_0_reg
				      ,input [31:0] rd_req_desc_1_axaddr_1_reg
				      ,input [31:0] rd_req_desc_1_axaddr_2_reg
				      ,input [31:0] rd_req_desc_1_axaddr_3_reg
				      ,input [31:0] rd_req_desc_1_axid_0_reg
				      ,input [31:0] rd_req_desc_1_axid_1_reg
				      ,input [31:0] rd_req_desc_1_axid_2_reg
				      ,input [31:0] rd_req_desc_1_axid_3_reg
				      ,input [31:0] rd_req_desc_1_axuser_0_reg
				      ,input [31:0] rd_req_desc_1_axuser_1_reg
				      ,input [31:0] rd_req_desc_1_axuser_2_reg
				      ,input [31:0] rd_req_desc_1_axuser_3_reg
				      ,input [31:0] rd_req_desc_1_axuser_4_reg
				      ,input [31:0] rd_req_desc_1_axuser_5_reg
				      ,input [31:0] rd_req_desc_1_axuser_6_reg
				      ,input [31:0] rd_req_desc_1_axuser_7_reg
				      ,input [31:0] rd_req_desc_1_axuser_8_reg
				      ,input [31:0] rd_req_desc_1_axuser_9_reg
				      ,input [31:0] rd_req_desc_1_axuser_10_reg
				      ,input [31:0] rd_req_desc_1_axuser_11_reg
				      ,input [31:0] rd_req_desc_1_axuser_12_reg
				      ,input [31:0] rd_req_desc_1_axuser_13_reg
				      ,input [31:0] rd_req_desc_1_axuser_14_reg
				      ,input [31:0] rd_req_desc_1_axuser_15_reg
				      ,input [31:0] rd_resp_desc_1_data_offset_reg
				      ,input [31:0] rd_resp_desc_1_data_size_reg
				      ,input [31:0] rd_resp_desc_1_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_1_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_1_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_1_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_1_resp_reg
				      ,input [31:0] rd_resp_desc_1_xid_0_reg
				      ,input [31:0] rd_resp_desc_1_xid_1_reg
				      ,input [31:0] rd_resp_desc_1_xid_2_reg
				      ,input [31:0] rd_resp_desc_1_xid_3_reg
				      ,input [31:0] rd_resp_desc_1_xuser_0_reg
				      ,input [31:0] rd_resp_desc_1_xuser_1_reg
				      ,input [31:0] rd_resp_desc_1_xuser_2_reg
				      ,input [31:0] rd_resp_desc_1_xuser_3_reg
				      ,input [31:0] rd_resp_desc_1_xuser_4_reg
				      ,input [31:0] rd_resp_desc_1_xuser_5_reg
				      ,input [31:0] rd_resp_desc_1_xuser_6_reg
				      ,input [31:0] rd_resp_desc_1_xuser_7_reg
				      ,input [31:0] rd_resp_desc_1_xuser_8_reg
				      ,input [31:0] rd_resp_desc_1_xuser_9_reg
				      ,input [31:0] rd_resp_desc_1_xuser_10_reg
				      ,input [31:0] rd_resp_desc_1_xuser_11_reg
				      ,input [31:0] rd_resp_desc_1_xuser_12_reg
				      ,input [31:0] rd_resp_desc_1_xuser_13_reg
				      ,input [31:0] rd_resp_desc_1_xuser_14_reg
				      ,input [31:0] rd_resp_desc_1_xuser_15_reg
				      ,input [31:0] wr_req_desc_1_txn_type_reg
				      ,input [31:0] wr_req_desc_1_size_reg
				      ,input [31:0] wr_req_desc_1_data_offset_reg
				      ,input [31:0] wr_req_desc_1_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_1_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_1_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_1_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_1_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_1_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_1_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_1_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_1_axsize_reg
				      ,input [31:0] wr_req_desc_1_attr_reg
				      ,input [31:0] wr_req_desc_1_axaddr_0_reg
				      ,input [31:0] wr_req_desc_1_axaddr_1_reg
				      ,input [31:0] wr_req_desc_1_axaddr_2_reg
				      ,input [31:0] wr_req_desc_1_axaddr_3_reg
				      ,input [31:0] wr_req_desc_1_axid_0_reg
				      ,input [31:0] wr_req_desc_1_axid_1_reg
				      ,input [31:0] wr_req_desc_1_axid_2_reg
				      ,input [31:0] wr_req_desc_1_axid_3_reg
				      ,input [31:0] wr_req_desc_1_axuser_0_reg
				      ,input [31:0] wr_req_desc_1_axuser_1_reg
				      ,input [31:0] wr_req_desc_1_axuser_2_reg
				      ,input [31:0] wr_req_desc_1_axuser_3_reg
				      ,input [31:0] wr_req_desc_1_axuser_4_reg
				      ,input [31:0] wr_req_desc_1_axuser_5_reg
				      ,input [31:0] wr_req_desc_1_axuser_6_reg
				      ,input [31:0] wr_req_desc_1_axuser_7_reg
				      ,input [31:0] wr_req_desc_1_axuser_8_reg
				      ,input [31:0] wr_req_desc_1_axuser_9_reg
				      ,input [31:0] wr_req_desc_1_axuser_10_reg
				      ,input [31:0] wr_req_desc_1_axuser_11_reg
				      ,input [31:0] wr_req_desc_1_axuser_12_reg
				      ,input [31:0] wr_req_desc_1_axuser_13_reg
				      ,input [31:0] wr_req_desc_1_axuser_14_reg
				      ,input [31:0] wr_req_desc_1_axuser_15_reg
				      ,input [31:0] wr_req_desc_1_wuser_0_reg
				      ,input [31:0] wr_req_desc_1_wuser_1_reg
				      ,input [31:0] wr_req_desc_1_wuser_2_reg
				      ,input [31:0] wr_req_desc_1_wuser_3_reg
				      ,input [31:0] wr_req_desc_1_wuser_4_reg
				      ,input [31:0] wr_req_desc_1_wuser_5_reg
				      ,input [31:0] wr_req_desc_1_wuser_6_reg
				      ,input [31:0] wr_req_desc_1_wuser_7_reg
				      ,input [31:0] wr_req_desc_1_wuser_8_reg
				      ,input [31:0] wr_req_desc_1_wuser_9_reg
				      ,input [31:0] wr_req_desc_1_wuser_10_reg
				      ,input [31:0] wr_req_desc_1_wuser_11_reg
				      ,input [31:0] wr_req_desc_1_wuser_12_reg
				      ,input [31:0] wr_req_desc_1_wuser_13_reg
				      ,input [31:0] wr_req_desc_1_wuser_14_reg
				      ,input [31:0] wr_req_desc_1_wuser_15_reg
				      ,input [31:0] wr_resp_desc_1_resp_reg
				      ,input [31:0] wr_resp_desc_1_xid_0_reg
				      ,input [31:0] wr_resp_desc_1_xid_1_reg
				      ,input [31:0] wr_resp_desc_1_xid_2_reg
				      ,input [31:0] wr_resp_desc_1_xid_3_reg
				      ,input [31:0] wr_resp_desc_1_xuser_0_reg
				      ,input [31:0] wr_resp_desc_1_xuser_1_reg
				      ,input [31:0] wr_resp_desc_1_xuser_2_reg
				      ,input [31:0] wr_resp_desc_1_xuser_3_reg
				      ,input [31:0] wr_resp_desc_1_xuser_4_reg
				      ,input [31:0] wr_resp_desc_1_xuser_5_reg
				      ,input [31:0] wr_resp_desc_1_xuser_6_reg
				      ,input [31:0] wr_resp_desc_1_xuser_7_reg
				      ,input [31:0] wr_resp_desc_1_xuser_8_reg
				      ,input [31:0] wr_resp_desc_1_xuser_9_reg
				      ,input [31:0] wr_resp_desc_1_xuser_10_reg
				      ,input [31:0] wr_resp_desc_1_xuser_11_reg
				      ,input [31:0] wr_resp_desc_1_xuser_12_reg
				      ,input [31:0] wr_resp_desc_1_xuser_13_reg
				      ,input [31:0] wr_resp_desc_1_xuser_14_reg
				      ,input [31:0] wr_resp_desc_1_xuser_15_reg
				      ,input [31:0] sn_req_desc_1_attr_reg
				      ,input [31:0] sn_req_desc_1_acaddr_0_reg
				      ,input [31:0] sn_req_desc_1_acaddr_1_reg
				      ,input [31:0] sn_req_desc_1_acaddr_2_reg
				      ,input [31:0] sn_req_desc_1_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_1_resp_reg
				      ,input [31:0] rd_req_desc_2_txn_type_reg
				      ,input [31:0] rd_req_desc_2_size_reg
				      ,input [31:0] rd_req_desc_2_axsize_reg
				      ,input [31:0] rd_req_desc_2_attr_reg
				      ,input [31:0] rd_req_desc_2_axaddr_0_reg
				      ,input [31:0] rd_req_desc_2_axaddr_1_reg
				      ,input [31:0] rd_req_desc_2_axaddr_2_reg
				      ,input [31:0] rd_req_desc_2_axaddr_3_reg
				      ,input [31:0] rd_req_desc_2_axid_0_reg
				      ,input [31:0] rd_req_desc_2_axid_1_reg
				      ,input [31:0] rd_req_desc_2_axid_2_reg
				      ,input [31:0] rd_req_desc_2_axid_3_reg
				      ,input [31:0] rd_req_desc_2_axuser_0_reg
				      ,input [31:0] rd_req_desc_2_axuser_1_reg
				      ,input [31:0] rd_req_desc_2_axuser_2_reg
				      ,input [31:0] rd_req_desc_2_axuser_3_reg
				      ,input [31:0] rd_req_desc_2_axuser_4_reg
				      ,input [31:0] rd_req_desc_2_axuser_5_reg
				      ,input [31:0] rd_req_desc_2_axuser_6_reg
				      ,input [31:0] rd_req_desc_2_axuser_7_reg
				      ,input [31:0] rd_req_desc_2_axuser_8_reg
				      ,input [31:0] rd_req_desc_2_axuser_9_reg
				      ,input [31:0] rd_req_desc_2_axuser_10_reg
				      ,input [31:0] rd_req_desc_2_axuser_11_reg
				      ,input [31:0] rd_req_desc_2_axuser_12_reg
				      ,input [31:0] rd_req_desc_2_axuser_13_reg
				      ,input [31:0] rd_req_desc_2_axuser_14_reg
				      ,input [31:0] rd_req_desc_2_axuser_15_reg
				      ,input [31:0] rd_resp_desc_2_data_offset_reg
				      ,input [31:0] rd_resp_desc_2_data_size_reg
				      ,input [31:0] rd_resp_desc_2_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_2_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_2_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_2_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_2_resp_reg
				      ,input [31:0] rd_resp_desc_2_xid_0_reg
				      ,input [31:0] rd_resp_desc_2_xid_1_reg
				      ,input [31:0] rd_resp_desc_2_xid_2_reg
				      ,input [31:0] rd_resp_desc_2_xid_3_reg
				      ,input [31:0] rd_resp_desc_2_xuser_0_reg
				      ,input [31:0] rd_resp_desc_2_xuser_1_reg
				      ,input [31:0] rd_resp_desc_2_xuser_2_reg
				      ,input [31:0] rd_resp_desc_2_xuser_3_reg
				      ,input [31:0] rd_resp_desc_2_xuser_4_reg
				      ,input [31:0] rd_resp_desc_2_xuser_5_reg
				      ,input [31:0] rd_resp_desc_2_xuser_6_reg
				      ,input [31:0] rd_resp_desc_2_xuser_7_reg
				      ,input [31:0] rd_resp_desc_2_xuser_8_reg
				      ,input [31:0] rd_resp_desc_2_xuser_9_reg
				      ,input [31:0] rd_resp_desc_2_xuser_10_reg
				      ,input [31:0] rd_resp_desc_2_xuser_11_reg
				      ,input [31:0] rd_resp_desc_2_xuser_12_reg
				      ,input [31:0] rd_resp_desc_2_xuser_13_reg
				      ,input [31:0] rd_resp_desc_2_xuser_14_reg
				      ,input [31:0] rd_resp_desc_2_xuser_15_reg
				      ,input [31:0] wr_req_desc_2_txn_type_reg
				      ,input [31:0] wr_req_desc_2_size_reg
				      ,input [31:0] wr_req_desc_2_data_offset_reg
				      ,input [31:0] wr_req_desc_2_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_2_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_2_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_2_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_2_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_2_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_2_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_2_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_2_axsize_reg
				      ,input [31:0] wr_req_desc_2_attr_reg
				      ,input [31:0] wr_req_desc_2_axaddr_0_reg
				      ,input [31:0] wr_req_desc_2_axaddr_1_reg
				      ,input [31:0] wr_req_desc_2_axaddr_2_reg
				      ,input [31:0] wr_req_desc_2_axaddr_3_reg
				      ,input [31:0] wr_req_desc_2_axid_0_reg
				      ,input [31:0] wr_req_desc_2_axid_1_reg
				      ,input [31:0] wr_req_desc_2_axid_2_reg
				      ,input [31:0] wr_req_desc_2_axid_3_reg
				      ,input [31:0] wr_req_desc_2_axuser_0_reg
				      ,input [31:0] wr_req_desc_2_axuser_1_reg
				      ,input [31:0] wr_req_desc_2_axuser_2_reg
				      ,input [31:0] wr_req_desc_2_axuser_3_reg
				      ,input [31:0] wr_req_desc_2_axuser_4_reg
				      ,input [31:0] wr_req_desc_2_axuser_5_reg
				      ,input [31:0] wr_req_desc_2_axuser_6_reg
				      ,input [31:0] wr_req_desc_2_axuser_7_reg
				      ,input [31:0] wr_req_desc_2_axuser_8_reg
				      ,input [31:0] wr_req_desc_2_axuser_9_reg
				      ,input [31:0] wr_req_desc_2_axuser_10_reg
				      ,input [31:0] wr_req_desc_2_axuser_11_reg
				      ,input [31:0] wr_req_desc_2_axuser_12_reg
				      ,input [31:0] wr_req_desc_2_axuser_13_reg
				      ,input [31:0] wr_req_desc_2_axuser_14_reg
				      ,input [31:0] wr_req_desc_2_axuser_15_reg
				      ,input [31:0] wr_req_desc_2_wuser_0_reg
				      ,input [31:0] wr_req_desc_2_wuser_1_reg
				      ,input [31:0] wr_req_desc_2_wuser_2_reg
				      ,input [31:0] wr_req_desc_2_wuser_3_reg
				      ,input [31:0] wr_req_desc_2_wuser_4_reg
				      ,input [31:0] wr_req_desc_2_wuser_5_reg
				      ,input [31:0] wr_req_desc_2_wuser_6_reg
				      ,input [31:0] wr_req_desc_2_wuser_7_reg
				      ,input [31:0] wr_req_desc_2_wuser_8_reg
				      ,input [31:0] wr_req_desc_2_wuser_9_reg
				      ,input [31:0] wr_req_desc_2_wuser_10_reg
				      ,input [31:0] wr_req_desc_2_wuser_11_reg
				      ,input [31:0] wr_req_desc_2_wuser_12_reg
				      ,input [31:0] wr_req_desc_2_wuser_13_reg
				      ,input [31:0] wr_req_desc_2_wuser_14_reg
				      ,input [31:0] wr_req_desc_2_wuser_15_reg
				      ,input [31:0] wr_resp_desc_2_resp_reg
				      ,input [31:0] wr_resp_desc_2_xid_0_reg
				      ,input [31:0] wr_resp_desc_2_xid_1_reg
				      ,input [31:0] wr_resp_desc_2_xid_2_reg
				      ,input [31:0] wr_resp_desc_2_xid_3_reg
				      ,input [31:0] wr_resp_desc_2_xuser_0_reg
				      ,input [31:0] wr_resp_desc_2_xuser_1_reg
				      ,input [31:0] wr_resp_desc_2_xuser_2_reg
				      ,input [31:0] wr_resp_desc_2_xuser_3_reg
				      ,input [31:0] wr_resp_desc_2_xuser_4_reg
				      ,input [31:0] wr_resp_desc_2_xuser_5_reg
				      ,input [31:0] wr_resp_desc_2_xuser_6_reg
				      ,input [31:0] wr_resp_desc_2_xuser_7_reg
				      ,input [31:0] wr_resp_desc_2_xuser_8_reg
				      ,input [31:0] wr_resp_desc_2_xuser_9_reg
				      ,input [31:0] wr_resp_desc_2_xuser_10_reg
				      ,input [31:0] wr_resp_desc_2_xuser_11_reg
				      ,input [31:0] wr_resp_desc_2_xuser_12_reg
				      ,input [31:0] wr_resp_desc_2_xuser_13_reg
				      ,input [31:0] wr_resp_desc_2_xuser_14_reg
				      ,input [31:0] wr_resp_desc_2_xuser_15_reg
				      ,input [31:0] sn_req_desc_2_attr_reg
				      ,input [31:0] sn_req_desc_2_acaddr_0_reg
				      ,input [31:0] sn_req_desc_2_acaddr_1_reg
				      ,input [31:0] sn_req_desc_2_acaddr_2_reg
				      ,input [31:0] sn_req_desc_2_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_2_resp_reg
				      ,input [31:0] rd_req_desc_3_txn_type_reg
				      ,input [31:0] rd_req_desc_3_size_reg
				      ,input [31:0] rd_req_desc_3_axsize_reg
				      ,input [31:0] rd_req_desc_3_attr_reg
				      ,input [31:0] rd_req_desc_3_axaddr_0_reg
				      ,input [31:0] rd_req_desc_3_axaddr_1_reg
				      ,input [31:0] rd_req_desc_3_axaddr_2_reg
				      ,input [31:0] rd_req_desc_3_axaddr_3_reg
				      ,input [31:0] rd_req_desc_3_axid_0_reg
				      ,input [31:0] rd_req_desc_3_axid_1_reg
				      ,input [31:0] rd_req_desc_3_axid_2_reg
				      ,input [31:0] rd_req_desc_3_axid_3_reg
				      ,input [31:0] rd_req_desc_3_axuser_0_reg
				      ,input [31:0] rd_req_desc_3_axuser_1_reg
				      ,input [31:0] rd_req_desc_3_axuser_2_reg
				      ,input [31:0] rd_req_desc_3_axuser_3_reg
				      ,input [31:0] rd_req_desc_3_axuser_4_reg
				      ,input [31:0] rd_req_desc_3_axuser_5_reg
				      ,input [31:0] rd_req_desc_3_axuser_6_reg
				      ,input [31:0] rd_req_desc_3_axuser_7_reg
				      ,input [31:0] rd_req_desc_3_axuser_8_reg
				      ,input [31:0] rd_req_desc_3_axuser_9_reg
				      ,input [31:0] rd_req_desc_3_axuser_10_reg
				      ,input [31:0] rd_req_desc_3_axuser_11_reg
				      ,input [31:0] rd_req_desc_3_axuser_12_reg
				      ,input [31:0] rd_req_desc_3_axuser_13_reg
				      ,input [31:0] rd_req_desc_3_axuser_14_reg
				      ,input [31:0] rd_req_desc_3_axuser_15_reg
				      ,input [31:0] rd_resp_desc_3_data_offset_reg
				      ,input [31:0] rd_resp_desc_3_data_size_reg
				      ,input [31:0] rd_resp_desc_3_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_3_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_3_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_3_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_3_resp_reg
				      ,input [31:0] rd_resp_desc_3_xid_0_reg
				      ,input [31:0] rd_resp_desc_3_xid_1_reg
				      ,input [31:0] rd_resp_desc_3_xid_2_reg
				      ,input [31:0] rd_resp_desc_3_xid_3_reg
				      ,input [31:0] rd_resp_desc_3_xuser_0_reg
				      ,input [31:0] rd_resp_desc_3_xuser_1_reg
				      ,input [31:0] rd_resp_desc_3_xuser_2_reg
				      ,input [31:0] rd_resp_desc_3_xuser_3_reg
				      ,input [31:0] rd_resp_desc_3_xuser_4_reg
				      ,input [31:0] rd_resp_desc_3_xuser_5_reg
				      ,input [31:0] rd_resp_desc_3_xuser_6_reg
				      ,input [31:0] rd_resp_desc_3_xuser_7_reg
				      ,input [31:0] rd_resp_desc_3_xuser_8_reg
				      ,input [31:0] rd_resp_desc_3_xuser_9_reg
				      ,input [31:0] rd_resp_desc_3_xuser_10_reg
				      ,input [31:0] rd_resp_desc_3_xuser_11_reg
				      ,input [31:0] rd_resp_desc_3_xuser_12_reg
				      ,input [31:0] rd_resp_desc_3_xuser_13_reg
				      ,input [31:0] rd_resp_desc_3_xuser_14_reg
				      ,input [31:0] rd_resp_desc_3_xuser_15_reg
				      ,input [31:0] wr_req_desc_3_txn_type_reg
				      ,input [31:0] wr_req_desc_3_size_reg
				      ,input [31:0] wr_req_desc_3_data_offset_reg
				      ,input [31:0] wr_req_desc_3_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_3_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_3_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_3_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_3_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_3_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_3_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_3_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_3_axsize_reg
				      ,input [31:0] wr_req_desc_3_attr_reg
				      ,input [31:0] wr_req_desc_3_axaddr_0_reg
				      ,input [31:0] wr_req_desc_3_axaddr_1_reg
				      ,input [31:0] wr_req_desc_3_axaddr_2_reg
				      ,input [31:0] wr_req_desc_3_axaddr_3_reg
				      ,input [31:0] wr_req_desc_3_axid_0_reg
				      ,input [31:0] wr_req_desc_3_axid_1_reg
				      ,input [31:0] wr_req_desc_3_axid_2_reg
				      ,input [31:0] wr_req_desc_3_axid_3_reg
				      ,input [31:0] wr_req_desc_3_axuser_0_reg
				      ,input [31:0] wr_req_desc_3_axuser_1_reg
				      ,input [31:0] wr_req_desc_3_axuser_2_reg
				      ,input [31:0] wr_req_desc_3_axuser_3_reg
				      ,input [31:0] wr_req_desc_3_axuser_4_reg
				      ,input [31:0] wr_req_desc_3_axuser_5_reg
				      ,input [31:0] wr_req_desc_3_axuser_6_reg
				      ,input [31:0] wr_req_desc_3_axuser_7_reg
				      ,input [31:0] wr_req_desc_3_axuser_8_reg
				      ,input [31:0] wr_req_desc_3_axuser_9_reg
				      ,input [31:0] wr_req_desc_3_axuser_10_reg
				      ,input [31:0] wr_req_desc_3_axuser_11_reg
				      ,input [31:0] wr_req_desc_3_axuser_12_reg
				      ,input [31:0] wr_req_desc_3_axuser_13_reg
				      ,input [31:0] wr_req_desc_3_axuser_14_reg
				      ,input [31:0] wr_req_desc_3_axuser_15_reg
				      ,input [31:0] wr_req_desc_3_wuser_0_reg
				      ,input [31:0] wr_req_desc_3_wuser_1_reg
				      ,input [31:0] wr_req_desc_3_wuser_2_reg
				      ,input [31:0] wr_req_desc_3_wuser_3_reg
				      ,input [31:0] wr_req_desc_3_wuser_4_reg
				      ,input [31:0] wr_req_desc_3_wuser_5_reg
				      ,input [31:0] wr_req_desc_3_wuser_6_reg
				      ,input [31:0] wr_req_desc_3_wuser_7_reg
				      ,input [31:0] wr_req_desc_3_wuser_8_reg
				      ,input [31:0] wr_req_desc_3_wuser_9_reg
				      ,input [31:0] wr_req_desc_3_wuser_10_reg
				      ,input [31:0] wr_req_desc_3_wuser_11_reg
				      ,input [31:0] wr_req_desc_3_wuser_12_reg
				      ,input [31:0] wr_req_desc_3_wuser_13_reg
				      ,input [31:0] wr_req_desc_3_wuser_14_reg
				      ,input [31:0] wr_req_desc_3_wuser_15_reg
				      ,input [31:0] wr_resp_desc_3_resp_reg
				      ,input [31:0] wr_resp_desc_3_xid_0_reg
				      ,input [31:0] wr_resp_desc_3_xid_1_reg
				      ,input [31:0] wr_resp_desc_3_xid_2_reg
				      ,input [31:0] wr_resp_desc_3_xid_3_reg
				      ,input [31:0] wr_resp_desc_3_xuser_0_reg
				      ,input [31:0] wr_resp_desc_3_xuser_1_reg
				      ,input [31:0] wr_resp_desc_3_xuser_2_reg
				      ,input [31:0] wr_resp_desc_3_xuser_3_reg
				      ,input [31:0] wr_resp_desc_3_xuser_4_reg
				      ,input [31:0] wr_resp_desc_3_xuser_5_reg
				      ,input [31:0] wr_resp_desc_3_xuser_6_reg
				      ,input [31:0] wr_resp_desc_3_xuser_7_reg
				      ,input [31:0] wr_resp_desc_3_xuser_8_reg
				      ,input [31:0] wr_resp_desc_3_xuser_9_reg
				      ,input [31:0] wr_resp_desc_3_xuser_10_reg
				      ,input [31:0] wr_resp_desc_3_xuser_11_reg
				      ,input [31:0] wr_resp_desc_3_xuser_12_reg
				      ,input [31:0] wr_resp_desc_3_xuser_13_reg
				      ,input [31:0] wr_resp_desc_3_xuser_14_reg
				      ,input [31:0] wr_resp_desc_3_xuser_15_reg
				      ,input [31:0] sn_req_desc_3_attr_reg
				      ,input [31:0] sn_req_desc_3_acaddr_0_reg
				      ,input [31:0] sn_req_desc_3_acaddr_1_reg
				      ,input [31:0] sn_req_desc_3_acaddr_2_reg
				      ,input [31:0] sn_req_desc_3_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_3_resp_reg
				      ,input [31:0] rd_req_desc_4_txn_type_reg
				      ,input [31:0] rd_req_desc_4_size_reg
				      ,input [31:0] rd_req_desc_4_axsize_reg
				      ,input [31:0] rd_req_desc_4_attr_reg
				      ,input [31:0] rd_req_desc_4_axaddr_0_reg
				      ,input [31:0] rd_req_desc_4_axaddr_1_reg
				      ,input [31:0] rd_req_desc_4_axaddr_2_reg
				      ,input [31:0] rd_req_desc_4_axaddr_3_reg
				      ,input [31:0] rd_req_desc_4_axid_0_reg
				      ,input [31:0] rd_req_desc_4_axid_1_reg
				      ,input [31:0] rd_req_desc_4_axid_2_reg
				      ,input [31:0] rd_req_desc_4_axid_3_reg
				      ,input [31:0] rd_req_desc_4_axuser_0_reg
				      ,input [31:0] rd_req_desc_4_axuser_1_reg
				      ,input [31:0] rd_req_desc_4_axuser_2_reg
				      ,input [31:0] rd_req_desc_4_axuser_3_reg
				      ,input [31:0] rd_req_desc_4_axuser_4_reg
				      ,input [31:0] rd_req_desc_4_axuser_5_reg
				      ,input [31:0] rd_req_desc_4_axuser_6_reg
				      ,input [31:0] rd_req_desc_4_axuser_7_reg
				      ,input [31:0] rd_req_desc_4_axuser_8_reg
				      ,input [31:0] rd_req_desc_4_axuser_9_reg
				      ,input [31:0] rd_req_desc_4_axuser_10_reg
				      ,input [31:0] rd_req_desc_4_axuser_11_reg
				      ,input [31:0] rd_req_desc_4_axuser_12_reg
				      ,input [31:0] rd_req_desc_4_axuser_13_reg
				      ,input [31:0] rd_req_desc_4_axuser_14_reg
				      ,input [31:0] rd_req_desc_4_axuser_15_reg
				      ,input [31:0] rd_resp_desc_4_data_offset_reg
				      ,input [31:0] rd_resp_desc_4_data_size_reg
				      ,input [31:0] rd_resp_desc_4_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_4_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_4_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_4_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_4_resp_reg
				      ,input [31:0] rd_resp_desc_4_xid_0_reg
				      ,input [31:0] rd_resp_desc_4_xid_1_reg
				      ,input [31:0] rd_resp_desc_4_xid_2_reg
				      ,input [31:0] rd_resp_desc_4_xid_3_reg
				      ,input [31:0] rd_resp_desc_4_xuser_0_reg
				      ,input [31:0] rd_resp_desc_4_xuser_1_reg
				      ,input [31:0] rd_resp_desc_4_xuser_2_reg
				      ,input [31:0] rd_resp_desc_4_xuser_3_reg
				      ,input [31:0] rd_resp_desc_4_xuser_4_reg
				      ,input [31:0] rd_resp_desc_4_xuser_5_reg
				      ,input [31:0] rd_resp_desc_4_xuser_6_reg
				      ,input [31:0] rd_resp_desc_4_xuser_7_reg
				      ,input [31:0] rd_resp_desc_4_xuser_8_reg
				      ,input [31:0] rd_resp_desc_4_xuser_9_reg
				      ,input [31:0] rd_resp_desc_4_xuser_10_reg
				      ,input [31:0] rd_resp_desc_4_xuser_11_reg
				      ,input [31:0] rd_resp_desc_4_xuser_12_reg
				      ,input [31:0] rd_resp_desc_4_xuser_13_reg
				      ,input [31:0] rd_resp_desc_4_xuser_14_reg
				      ,input [31:0] rd_resp_desc_4_xuser_15_reg
				      ,input [31:0] wr_req_desc_4_txn_type_reg
				      ,input [31:0] wr_req_desc_4_size_reg
				      ,input [31:0] wr_req_desc_4_data_offset_reg
				      ,input [31:0] wr_req_desc_4_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_4_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_4_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_4_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_4_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_4_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_4_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_4_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_4_axsize_reg
				      ,input [31:0] wr_req_desc_4_attr_reg
				      ,input [31:0] wr_req_desc_4_axaddr_0_reg
				      ,input [31:0] wr_req_desc_4_axaddr_1_reg
				      ,input [31:0] wr_req_desc_4_axaddr_2_reg
				      ,input [31:0] wr_req_desc_4_axaddr_3_reg
				      ,input [31:0] wr_req_desc_4_axid_0_reg
				      ,input [31:0] wr_req_desc_4_axid_1_reg
				      ,input [31:0] wr_req_desc_4_axid_2_reg
				      ,input [31:0] wr_req_desc_4_axid_3_reg
				      ,input [31:0] wr_req_desc_4_axuser_0_reg
				      ,input [31:0] wr_req_desc_4_axuser_1_reg
				      ,input [31:0] wr_req_desc_4_axuser_2_reg
				      ,input [31:0] wr_req_desc_4_axuser_3_reg
				      ,input [31:0] wr_req_desc_4_axuser_4_reg
				      ,input [31:0] wr_req_desc_4_axuser_5_reg
				      ,input [31:0] wr_req_desc_4_axuser_6_reg
				      ,input [31:0] wr_req_desc_4_axuser_7_reg
				      ,input [31:0] wr_req_desc_4_axuser_8_reg
				      ,input [31:0] wr_req_desc_4_axuser_9_reg
				      ,input [31:0] wr_req_desc_4_axuser_10_reg
				      ,input [31:0] wr_req_desc_4_axuser_11_reg
				      ,input [31:0] wr_req_desc_4_axuser_12_reg
				      ,input [31:0] wr_req_desc_4_axuser_13_reg
				      ,input [31:0] wr_req_desc_4_axuser_14_reg
				      ,input [31:0] wr_req_desc_4_axuser_15_reg
				      ,input [31:0] wr_req_desc_4_wuser_0_reg
				      ,input [31:0] wr_req_desc_4_wuser_1_reg
				      ,input [31:0] wr_req_desc_4_wuser_2_reg
				      ,input [31:0] wr_req_desc_4_wuser_3_reg
				      ,input [31:0] wr_req_desc_4_wuser_4_reg
				      ,input [31:0] wr_req_desc_4_wuser_5_reg
				      ,input [31:0] wr_req_desc_4_wuser_6_reg
				      ,input [31:0] wr_req_desc_4_wuser_7_reg
				      ,input [31:0] wr_req_desc_4_wuser_8_reg
				      ,input [31:0] wr_req_desc_4_wuser_9_reg
				      ,input [31:0] wr_req_desc_4_wuser_10_reg
				      ,input [31:0] wr_req_desc_4_wuser_11_reg
				      ,input [31:0] wr_req_desc_4_wuser_12_reg
				      ,input [31:0] wr_req_desc_4_wuser_13_reg
				      ,input [31:0] wr_req_desc_4_wuser_14_reg
				      ,input [31:0] wr_req_desc_4_wuser_15_reg
				      ,input [31:0] wr_resp_desc_4_resp_reg
				      ,input [31:0] wr_resp_desc_4_xid_0_reg
				      ,input [31:0] wr_resp_desc_4_xid_1_reg
				      ,input [31:0] wr_resp_desc_4_xid_2_reg
				      ,input [31:0] wr_resp_desc_4_xid_3_reg
				      ,input [31:0] wr_resp_desc_4_xuser_0_reg
				      ,input [31:0] wr_resp_desc_4_xuser_1_reg
				      ,input [31:0] wr_resp_desc_4_xuser_2_reg
				      ,input [31:0] wr_resp_desc_4_xuser_3_reg
				      ,input [31:0] wr_resp_desc_4_xuser_4_reg
				      ,input [31:0] wr_resp_desc_4_xuser_5_reg
				      ,input [31:0] wr_resp_desc_4_xuser_6_reg
				      ,input [31:0] wr_resp_desc_4_xuser_7_reg
				      ,input [31:0] wr_resp_desc_4_xuser_8_reg
				      ,input [31:0] wr_resp_desc_4_xuser_9_reg
				      ,input [31:0] wr_resp_desc_4_xuser_10_reg
				      ,input [31:0] wr_resp_desc_4_xuser_11_reg
				      ,input [31:0] wr_resp_desc_4_xuser_12_reg
				      ,input [31:0] wr_resp_desc_4_xuser_13_reg
				      ,input [31:0] wr_resp_desc_4_xuser_14_reg
				      ,input [31:0] wr_resp_desc_4_xuser_15_reg
				      ,input [31:0] sn_req_desc_4_attr_reg
				      ,input [31:0] sn_req_desc_4_acaddr_0_reg
				      ,input [31:0] sn_req_desc_4_acaddr_1_reg
				      ,input [31:0] sn_req_desc_4_acaddr_2_reg
				      ,input [31:0] sn_req_desc_4_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_4_resp_reg
				      ,input [31:0] rd_req_desc_5_txn_type_reg
				      ,input [31:0] rd_req_desc_5_size_reg
				      ,input [31:0] rd_req_desc_5_axsize_reg
				      ,input [31:0] rd_req_desc_5_attr_reg
				      ,input [31:0] rd_req_desc_5_axaddr_0_reg
				      ,input [31:0] rd_req_desc_5_axaddr_1_reg
				      ,input [31:0] rd_req_desc_5_axaddr_2_reg
				      ,input [31:0] rd_req_desc_5_axaddr_3_reg
				      ,input [31:0] rd_req_desc_5_axid_0_reg
				      ,input [31:0] rd_req_desc_5_axid_1_reg
				      ,input [31:0] rd_req_desc_5_axid_2_reg
				      ,input [31:0] rd_req_desc_5_axid_3_reg
				      ,input [31:0] rd_req_desc_5_axuser_0_reg
				      ,input [31:0] rd_req_desc_5_axuser_1_reg
				      ,input [31:0] rd_req_desc_5_axuser_2_reg
				      ,input [31:0] rd_req_desc_5_axuser_3_reg
				      ,input [31:0] rd_req_desc_5_axuser_4_reg
				      ,input [31:0] rd_req_desc_5_axuser_5_reg
				      ,input [31:0] rd_req_desc_5_axuser_6_reg
				      ,input [31:0] rd_req_desc_5_axuser_7_reg
				      ,input [31:0] rd_req_desc_5_axuser_8_reg
				      ,input [31:0] rd_req_desc_5_axuser_9_reg
				      ,input [31:0] rd_req_desc_5_axuser_10_reg
				      ,input [31:0] rd_req_desc_5_axuser_11_reg
				      ,input [31:0] rd_req_desc_5_axuser_12_reg
				      ,input [31:0] rd_req_desc_5_axuser_13_reg
				      ,input [31:0] rd_req_desc_5_axuser_14_reg
				      ,input [31:0] rd_req_desc_5_axuser_15_reg
				      ,input [31:0] rd_resp_desc_5_data_offset_reg
				      ,input [31:0] rd_resp_desc_5_data_size_reg
				      ,input [31:0] rd_resp_desc_5_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_5_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_5_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_5_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_5_resp_reg
				      ,input [31:0] rd_resp_desc_5_xid_0_reg
				      ,input [31:0] rd_resp_desc_5_xid_1_reg
				      ,input [31:0] rd_resp_desc_5_xid_2_reg
				      ,input [31:0] rd_resp_desc_5_xid_3_reg
				      ,input [31:0] rd_resp_desc_5_xuser_0_reg
				      ,input [31:0] rd_resp_desc_5_xuser_1_reg
				      ,input [31:0] rd_resp_desc_5_xuser_2_reg
				      ,input [31:0] rd_resp_desc_5_xuser_3_reg
				      ,input [31:0] rd_resp_desc_5_xuser_4_reg
				      ,input [31:0] rd_resp_desc_5_xuser_5_reg
				      ,input [31:0] rd_resp_desc_5_xuser_6_reg
				      ,input [31:0] rd_resp_desc_5_xuser_7_reg
				      ,input [31:0] rd_resp_desc_5_xuser_8_reg
				      ,input [31:0] rd_resp_desc_5_xuser_9_reg
				      ,input [31:0] rd_resp_desc_5_xuser_10_reg
				      ,input [31:0] rd_resp_desc_5_xuser_11_reg
				      ,input [31:0] rd_resp_desc_5_xuser_12_reg
				      ,input [31:0] rd_resp_desc_5_xuser_13_reg
				      ,input [31:0] rd_resp_desc_5_xuser_14_reg
				      ,input [31:0] rd_resp_desc_5_xuser_15_reg
				      ,input [31:0] wr_req_desc_5_txn_type_reg
				      ,input [31:0] wr_req_desc_5_size_reg
				      ,input [31:0] wr_req_desc_5_data_offset_reg
				      ,input [31:0] wr_req_desc_5_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_5_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_5_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_5_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_5_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_5_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_5_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_5_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_5_axsize_reg
				      ,input [31:0] wr_req_desc_5_attr_reg
				      ,input [31:0] wr_req_desc_5_axaddr_0_reg
				      ,input [31:0] wr_req_desc_5_axaddr_1_reg
				      ,input [31:0] wr_req_desc_5_axaddr_2_reg
				      ,input [31:0] wr_req_desc_5_axaddr_3_reg
				      ,input [31:0] wr_req_desc_5_axid_0_reg
				      ,input [31:0] wr_req_desc_5_axid_1_reg
				      ,input [31:0] wr_req_desc_5_axid_2_reg
				      ,input [31:0] wr_req_desc_5_axid_3_reg
				      ,input [31:0] wr_req_desc_5_axuser_0_reg
				      ,input [31:0] wr_req_desc_5_axuser_1_reg
				      ,input [31:0] wr_req_desc_5_axuser_2_reg
				      ,input [31:0] wr_req_desc_5_axuser_3_reg
				      ,input [31:0] wr_req_desc_5_axuser_4_reg
				      ,input [31:0] wr_req_desc_5_axuser_5_reg
				      ,input [31:0] wr_req_desc_5_axuser_6_reg
				      ,input [31:0] wr_req_desc_5_axuser_7_reg
				      ,input [31:0] wr_req_desc_5_axuser_8_reg
				      ,input [31:0] wr_req_desc_5_axuser_9_reg
				      ,input [31:0] wr_req_desc_5_axuser_10_reg
				      ,input [31:0] wr_req_desc_5_axuser_11_reg
				      ,input [31:0] wr_req_desc_5_axuser_12_reg
				      ,input [31:0] wr_req_desc_5_axuser_13_reg
				      ,input [31:0] wr_req_desc_5_axuser_14_reg
				      ,input [31:0] wr_req_desc_5_axuser_15_reg
				      ,input [31:0] wr_req_desc_5_wuser_0_reg
				      ,input [31:0] wr_req_desc_5_wuser_1_reg
				      ,input [31:0] wr_req_desc_5_wuser_2_reg
				      ,input [31:0] wr_req_desc_5_wuser_3_reg
				      ,input [31:0] wr_req_desc_5_wuser_4_reg
				      ,input [31:0] wr_req_desc_5_wuser_5_reg
				      ,input [31:0] wr_req_desc_5_wuser_6_reg
				      ,input [31:0] wr_req_desc_5_wuser_7_reg
				      ,input [31:0] wr_req_desc_5_wuser_8_reg
				      ,input [31:0] wr_req_desc_5_wuser_9_reg
				      ,input [31:0] wr_req_desc_5_wuser_10_reg
				      ,input [31:0] wr_req_desc_5_wuser_11_reg
				      ,input [31:0] wr_req_desc_5_wuser_12_reg
				      ,input [31:0] wr_req_desc_5_wuser_13_reg
				      ,input [31:0] wr_req_desc_5_wuser_14_reg
				      ,input [31:0] wr_req_desc_5_wuser_15_reg
				      ,input [31:0] wr_resp_desc_5_resp_reg
				      ,input [31:0] wr_resp_desc_5_xid_0_reg
				      ,input [31:0] wr_resp_desc_5_xid_1_reg
				      ,input [31:0] wr_resp_desc_5_xid_2_reg
				      ,input [31:0] wr_resp_desc_5_xid_3_reg
				      ,input [31:0] wr_resp_desc_5_xuser_0_reg
				      ,input [31:0] wr_resp_desc_5_xuser_1_reg
				      ,input [31:0] wr_resp_desc_5_xuser_2_reg
				      ,input [31:0] wr_resp_desc_5_xuser_3_reg
				      ,input [31:0] wr_resp_desc_5_xuser_4_reg
				      ,input [31:0] wr_resp_desc_5_xuser_5_reg
				      ,input [31:0] wr_resp_desc_5_xuser_6_reg
				      ,input [31:0] wr_resp_desc_5_xuser_7_reg
				      ,input [31:0] wr_resp_desc_5_xuser_8_reg
				      ,input [31:0] wr_resp_desc_5_xuser_9_reg
				      ,input [31:0] wr_resp_desc_5_xuser_10_reg
				      ,input [31:0] wr_resp_desc_5_xuser_11_reg
				      ,input [31:0] wr_resp_desc_5_xuser_12_reg
				      ,input [31:0] wr_resp_desc_5_xuser_13_reg
				      ,input [31:0] wr_resp_desc_5_xuser_14_reg
				      ,input [31:0] wr_resp_desc_5_xuser_15_reg
				      ,input [31:0] sn_req_desc_5_attr_reg
				      ,input [31:0] sn_req_desc_5_acaddr_0_reg
				      ,input [31:0] sn_req_desc_5_acaddr_1_reg
				      ,input [31:0] sn_req_desc_5_acaddr_2_reg
				      ,input [31:0] sn_req_desc_5_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_5_resp_reg
				      ,input [31:0] rd_req_desc_6_txn_type_reg
				      ,input [31:0] rd_req_desc_6_size_reg
				      ,input [31:0] rd_req_desc_6_axsize_reg
				      ,input [31:0] rd_req_desc_6_attr_reg
				      ,input [31:0] rd_req_desc_6_axaddr_0_reg
				      ,input [31:0] rd_req_desc_6_axaddr_1_reg
				      ,input [31:0] rd_req_desc_6_axaddr_2_reg
				      ,input [31:0] rd_req_desc_6_axaddr_3_reg
				      ,input [31:0] rd_req_desc_6_axid_0_reg
				      ,input [31:0] rd_req_desc_6_axid_1_reg
				      ,input [31:0] rd_req_desc_6_axid_2_reg
				      ,input [31:0] rd_req_desc_6_axid_3_reg
				      ,input [31:0] rd_req_desc_6_axuser_0_reg
				      ,input [31:0] rd_req_desc_6_axuser_1_reg
				      ,input [31:0] rd_req_desc_6_axuser_2_reg
				      ,input [31:0] rd_req_desc_6_axuser_3_reg
				      ,input [31:0] rd_req_desc_6_axuser_4_reg
				      ,input [31:0] rd_req_desc_6_axuser_5_reg
				      ,input [31:0] rd_req_desc_6_axuser_6_reg
				      ,input [31:0] rd_req_desc_6_axuser_7_reg
				      ,input [31:0] rd_req_desc_6_axuser_8_reg
				      ,input [31:0] rd_req_desc_6_axuser_9_reg
				      ,input [31:0] rd_req_desc_6_axuser_10_reg
				      ,input [31:0] rd_req_desc_6_axuser_11_reg
				      ,input [31:0] rd_req_desc_6_axuser_12_reg
				      ,input [31:0] rd_req_desc_6_axuser_13_reg
				      ,input [31:0] rd_req_desc_6_axuser_14_reg
				      ,input [31:0] rd_req_desc_6_axuser_15_reg
				      ,input [31:0] rd_resp_desc_6_data_offset_reg
				      ,input [31:0] rd_resp_desc_6_data_size_reg
				      ,input [31:0] rd_resp_desc_6_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_6_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_6_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_6_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_6_resp_reg
				      ,input [31:0] rd_resp_desc_6_xid_0_reg
				      ,input [31:0] rd_resp_desc_6_xid_1_reg
				      ,input [31:0] rd_resp_desc_6_xid_2_reg
				      ,input [31:0] rd_resp_desc_6_xid_3_reg
				      ,input [31:0] rd_resp_desc_6_xuser_0_reg
				      ,input [31:0] rd_resp_desc_6_xuser_1_reg
				      ,input [31:0] rd_resp_desc_6_xuser_2_reg
				      ,input [31:0] rd_resp_desc_6_xuser_3_reg
				      ,input [31:0] rd_resp_desc_6_xuser_4_reg
				      ,input [31:0] rd_resp_desc_6_xuser_5_reg
				      ,input [31:0] rd_resp_desc_6_xuser_6_reg
				      ,input [31:0] rd_resp_desc_6_xuser_7_reg
				      ,input [31:0] rd_resp_desc_6_xuser_8_reg
				      ,input [31:0] rd_resp_desc_6_xuser_9_reg
				      ,input [31:0] rd_resp_desc_6_xuser_10_reg
				      ,input [31:0] rd_resp_desc_6_xuser_11_reg
				      ,input [31:0] rd_resp_desc_6_xuser_12_reg
				      ,input [31:0] rd_resp_desc_6_xuser_13_reg
				      ,input [31:0] rd_resp_desc_6_xuser_14_reg
				      ,input [31:0] rd_resp_desc_6_xuser_15_reg
				      ,input [31:0] wr_req_desc_6_txn_type_reg
				      ,input [31:0] wr_req_desc_6_size_reg
				      ,input [31:0] wr_req_desc_6_data_offset_reg
				      ,input [31:0] wr_req_desc_6_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_6_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_6_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_6_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_6_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_6_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_6_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_6_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_6_axsize_reg
				      ,input [31:0] wr_req_desc_6_attr_reg
				      ,input [31:0] wr_req_desc_6_axaddr_0_reg
				      ,input [31:0] wr_req_desc_6_axaddr_1_reg
				      ,input [31:0] wr_req_desc_6_axaddr_2_reg
				      ,input [31:0] wr_req_desc_6_axaddr_3_reg
				      ,input [31:0] wr_req_desc_6_axid_0_reg
				      ,input [31:0] wr_req_desc_6_axid_1_reg
				      ,input [31:0] wr_req_desc_6_axid_2_reg
				      ,input [31:0] wr_req_desc_6_axid_3_reg
				      ,input [31:0] wr_req_desc_6_axuser_0_reg
				      ,input [31:0] wr_req_desc_6_axuser_1_reg
				      ,input [31:0] wr_req_desc_6_axuser_2_reg
				      ,input [31:0] wr_req_desc_6_axuser_3_reg
				      ,input [31:0] wr_req_desc_6_axuser_4_reg
				      ,input [31:0] wr_req_desc_6_axuser_5_reg
				      ,input [31:0] wr_req_desc_6_axuser_6_reg
				      ,input [31:0] wr_req_desc_6_axuser_7_reg
				      ,input [31:0] wr_req_desc_6_axuser_8_reg
				      ,input [31:0] wr_req_desc_6_axuser_9_reg
				      ,input [31:0] wr_req_desc_6_axuser_10_reg
				      ,input [31:0] wr_req_desc_6_axuser_11_reg
				      ,input [31:0] wr_req_desc_6_axuser_12_reg
				      ,input [31:0] wr_req_desc_6_axuser_13_reg
				      ,input [31:0] wr_req_desc_6_axuser_14_reg
				      ,input [31:0] wr_req_desc_6_axuser_15_reg
				      ,input [31:0] wr_req_desc_6_wuser_0_reg
				      ,input [31:0] wr_req_desc_6_wuser_1_reg
				      ,input [31:0] wr_req_desc_6_wuser_2_reg
				      ,input [31:0] wr_req_desc_6_wuser_3_reg
				      ,input [31:0] wr_req_desc_6_wuser_4_reg
				      ,input [31:0] wr_req_desc_6_wuser_5_reg
				      ,input [31:0] wr_req_desc_6_wuser_6_reg
				      ,input [31:0] wr_req_desc_6_wuser_7_reg
				      ,input [31:0] wr_req_desc_6_wuser_8_reg
				      ,input [31:0] wr_req_desc_6_wuser_9_reg
				      ,input [31:0] wr_req_desc_6_wuser_10_reg
				      ,input [31:0] wr_req_desc_6_wuser_11_reg
				      ,input [31:0] wr_req_desc_6_wuser_12_reg
				      ,input [31:0] wr_req_desc_6_wuser_13_reg
				      ,input [31:0] wr_req_desc_6_wuser_14_reg
				      ,input [31:0] wr_req_desc_6_wuser_15_reg
				      ,input [31:0] wr_resp_desc_6_resp_reg
				      ,input [31:0] wr_resp_desc_6_xid_0_reg
				      ,input [31:0] wr_resp_desc_6_xid_1_reg
				      ,input [31:0] wr_resp_desc_6_xid_2_reg
				      ,input [31:0] wr_resp_desc_6_xid_3_reg
				      ,input [31:0] wr_resp_desc_6_xuser_0_reg
				      ,input [31:0] wr_resp_desc_6_xuser_1_reg
				      ,input [31:0] wr_resp_desc_6_xuser_2_reg
				      ,input [31:0] wr_resp_desc_6_xuser_3_reg
				      ,input [31:0] wr_resp_desc_6_xuser_4_reg
				      ,input [31:0] wr_resp_desc_6_xuser_5_reg
				      ,input [31:0] wr_resp_desc_6_xuser_6_reg
				      ,input [31:0] wr_resp_desc_6_xuser_7_reg
				      ,input [31:0] wr_resp_desc_6_xuser_8_reg
				      ,input [31:0] wr_resp_desc_6_xuser_9_reg
				      ,input [31:0] wr_resp_desc_6_xuser_10_reg
				      ,input [31:0] wr_resp_desc_6_xuser_11_reg
				      ,input [31:0] wr_resp_desc_6_xuser_12_reg
				      ,input [31:0] wr_resp_desc_6_xuser_13_reg
				      ,input [31:0] wr_resp_desc_6_xuser_14_reg
				      ,input [31:0] wr_resp_desc_6_xuser_15_reg
				      ,input [31:0] sn_req_desc_6_attr_reg
				      ,input [31:0] sn_req_desc_6_acaddr_0_reg
				      ,input [31:0] sn_req_desc_6_acaddr_1_reg
				      ,input [31:0] sn_req_desc_6_acaddr_2_reg
				      ,input [31:0] sn_req_desc_6_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_6_resp_reg
				      ,input [31:0] rd_req_desc_7_txn_type_reg
				      ,input [31:0] rd_req_desc_7_size_reg
				      ,input [31:0] rd_req_desc_7_axsize_reg
				      ,input [31:0] rd_req_desc_7_attr_reg
				      ,input [31:0] rd_req_desc_7_axaddr_0_reg
				      ,input [31:0] rd_req_desc_7_axaddr_1_reg
				      ,input [31:0] rd_req_desc_7_axaddr_2_reg
				      ,input [31:0] rd_req_desc_7_axaddr_3_reg
				      ,input [31:0] rd_req_desc_7_axid_0_reg
				      ,input [31:0] rd_req_desc_7_axid_1_reg
				      ,input [31:0] rd_req_desc_7_axid_2_reg
				      ,input [31:0] rd_req_desc_7_axid_3_reg
				      ,input [31:0] rd_req_desc_7_axuser_0_reg
				      ,input [31:0] rd_req_desc_7_axuser_1_reg
				      ,input [31:0] rd_req_desc_7_axuser_2_reg
				      ,input [31:0] rd_req_desc_7_axuser_3_reg
				      ,input [31:0] rd_req_desc_7_axuser_4_reg
				      ,input [31:0] rd_req_desc_7_axuser_5_reg
				      ,input [31:0] rd_req_desc_7_axuser_6_reg
				      ,input [31:0] rd_req_desc_7_axuser_7_reg
				      ,input [31:0] rd_req_desc_7_axuser_8_reg
				      ,input [31:0] rd_req_desc_7_axuser_9_reg
				      ,input [31:0] rd_req_desc_7_axuser_10_reg
				      ,input [31:0] rd_req_desc_7_axuser_11_reg
				      ,input [31:0] rd_req_desc_7_axuser_12_reg
				      ,input [31:0] rd_req_desc_7_axuser_13_reg
				      ,input [31:0] rd_req_desc_7_axuser_14_reg
				      ,input [31:0] rd_req_desc_7_axuser_15_reg
				      ,input [31:0] rd_resp_desc_7_data_offset_reg
				      ,input [31:0] rd_resp_desc_7_data_size_reg
				      ,input [31:0] rd_resp_desc_7_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_7_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_7_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_7_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_7_resp_reg
				      ,input [31:0] rd_resp_desc_7_xid_0_reg
				      ,input [31:0] rd_resp_desc_7_xid_1_reg
				      ,input [31:0] rd_resp_desc_7_xid_2_reg
				      ,input [31:0] rd_resp_desc_7_xid_3_reg
				      ,input [31:0] rd_resp_desc_7_xuser_0_reg
				      ,input [31:0] rd_resp_desc_7_xuser_1_reg
				      ,input [31:0] rd_resp_desc_7_xuser_2_reg
				      ,input [31:0] rd_resp_desc_7_xuser_3_reg
				      ,input [31:0] rd_resp_desc_7_xuser_4_reg
				      ,input [31:0] rd_resp_desc_7_xuser_5_reg
				      ,input [31:0] rd_resp_desc_7_xuser_6_reg
				      ,input [31:0] rd_resp_desc_7_xuser_7_reg
				      ,input [31:0] rd_resp_desc_7_xuser_8_reg
				      ,input [31:0] rd_resp_desc_7_xuser_9_reg
				      ,input [31:0] rd_resp_desc_7_xuser_10_reg
				      ,input [31:0] rd_resp_desc_7_xuser_11_reg
				      ,input [31:0] rd_resp_desc_7_xuser_12_reg
				      ,input [31:0] rd_resp_desc_7_xuser_13_reg
				      ,input [31:0] rd_resp_desc_7_xuser_14_reg
				      ,input [31:0] rd_resp_desc_7_xuser_15_reg
				      ,input [31:0] wr_req_desc_7_txn_type_reg
				      ,input [31:0] wr_req_desc_7_size_reg
				      ,input [31:0] wr_req_desc_7_data_offset_reg
				      ,input [31:0] wr_req_desc_7_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_7_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_7_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_7_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_7_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_7_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_7_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_7_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_7_axsize_reg
				      ,input [31:0] wr_req_desc_7_attr_reg
				      ,input [31:0] wr_req_desc_7_axaddr_0_reg
				      ,input [31:0] wr_req_desc_7_axaddr_1_reg
				      ,input [31:0] wr_req_desc_7_axaddr_2_reg
				      ,input [31:0] wr_req_desc_7_axaddr_3_reg
				      ,input [31:0] wr_req_desc_7_axid_0_reg
				      ,input [31:0] wr_req_desc_7_axid_1_reg
				      ,input [31:0] wr_req_desc_7_axid_2_reg
				      ,input [31:0] wr_req_desc_7_axid_3_reg
				      ,input [31:0] wr_req_desc_7_axuser_0_reg
				      ,input [31:0] wr_req_desc_7_axuser_1_reg
				      ,input [31:0] wr_req_desc_7_axuser_2_reg
				      ,input [31:0] wr_req_desc_7_axuser_3_reg
				      ,input [31:0] wr_req_desc_7_axuser_4_reg
				      ,input [31:0] wr_req_desc_7_axuser_5_reg
				      ,input [31:0] wr_req_desc_7_axuser_6_reg
				      ,input [31:0] wr_req_desc_7_axuser_7_reg
				      ,input [31:0] wr_req_desc_7_axuser_8_reg
				      ,input [31:0] wr_req_desc_7_axuser_9_reg
				      ,input [31:0] wr_req_desc_7_axuser_10_reg
				      ,input [31:0] wr_req_desc_7_axuser_11_reg
				      ,input [31:0] wr_req_desc_7_axuser_12_reg
				      ,input [31:0] wr_req_desc_7_axuser_13_reg
				      ,input [31:0] wr_req_desc_7_axuser_14_reg
				      ,input [31:0] wr_req_desc_7_axuser_15_reg
				      ,input [31:0] wr_req_desc_7_wuser_0_reg
				      ,input [31:0] wr_req_desc_7_wuser_1_reg
				      ,input [31:0] wr_req_desc_7_wuser_2_reg
				      ,input [31:0] wr_req_desc_7_wuser_3_reg
				      ,input [31:0] wr_req_desc_7_wuser_4_reg
				      ,input [31:0] wr_req_desc_7_wuser_5_reg
				      ,input [31:0] wr_req_desc_7_wuser_6_reg
				      ,input [31:0] wr_req_desc_7_wuser_7_reg
				      ,input [31:0] wr_req_desc_7_wuser_8_reg
				      ,input [31:0] wr_req_desc_7_wuser_9_reg
				      ,input [31:0] wr_req_desc_7_wuser_10_reg
				      ,input [31:0] wr_req_desc_7_wuser_11_reg
				      ,input [31:0] wr_req_desc_7_wuser_12_reg
				      ,input [31:0] wr_req_desc_7_wuser_13_reg
				      ,input [31:0] wr_req_desc_7_wuser_14_reg
				      ,input [31:0] wr_req_desc_7_wuser_15_reg
				      ,input [31:0] wr_resp_desc_7_resp_reg
				      ,input [31:0] wr_resp_desc_7_xid_0_reg
				      ,input [31:0] wr_resp_desc_7_xid_1_reg
				      ,input [31:0] wr_resp_desc_7_xid_2_reg
				      ,input [31:0] wr_resp_desc_7_xid_3_reg
				      ,input [31:0] wr_resp_desc_7_xuser_0_reg
				      ,input [31:0] wr_resp_desc_7_xuser_1_reg
				      ,input [31:0] wr_resp_desc_7_xuser_2_reg
				      ,input [31:0] wr_resp_desc_7_xuser_3_reg
				      ,input [31:0] wr_resp_desc_7_xuser_4_reg
				      ,input [31:0] wr_resp_desc_7_xuser_5_reg
				      ,input [31:0] wr_resp_desc_7_xuser_6_reg
				      ,input [31:0] wr_resp_desc_7_xuser_7_reg
				      ,input [31:0] wr_resp_desc_7_xuser_8_reg
				      ,input [31:0] wr_resp_desc_7_xuser_9_reg
				      ,input [31:0] wr_resp_desc_7_xuser_10_reg
				      ,input [31:0] wr_resp_desc_7_xuser_11_reg
				      ,input [31:0] wr_resp_desc_7_xuser_12_reg
				      ,input [31:0] wr_resp_desc_7_xuser_13_reg
				      ,input [31:0] wr_resp_desc_7_xuser_14_reg
				      ,input [31:0] wr_resp_desc_7_xuser_15_reg
				      ,input [31:0] sn_req_desc_7_attr_reg
				      ,input [31:0] sn_req_desc_7_acaddr_0_reg
				      ,input [31:0] sn_req_desc_7_acaddr_1_reg
				      ,input [31:0] sn_req_desc_7_acaddr_2_reg
				      ,input [31:0] sn_req_desc_7_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_7_resp_reg
				      ,input [31:0] rd_req_desc_8_txn_type_reg
				      ,input [31:0] rd_req_desc_8_size_reg
				      ,input [31:0] rd_req_desc_8_axsize_reg
				      ,input [31:0] rd_req_desc_8_attr_reg
				      ,input [31:0] rd_req_desc_8_axaddr_0_reg
				      ,input [31:0] rd_req_desc_8_axaddr_1_reg
				      ,input [31:0] rd_req_desc_8_axaddr_2_reg
				      ,input [31:0] rd_req_desc_8_axaddr_3_reg
				      ,input [31:0] rd_req_desc_8_axid_0_reg
				      ,input [31:0] rd_req_desc_8_axid_1_reg
				      ,input [31:0] rd_req_desc_8_axid_2_reg
				      ,input [31:0] rd_req_desc_8_axid_3_reg
				      ,input [31:0] rd_req_desc_8_axuser_0_reg
				      ,input [31:0] rd_req_desc_8_axuser_1_reg
				      ,input [31:0] rd_req_desc_8_axuser_2_reg
				      ,input [31:0] rd_req_desc_8_axuser_3_reg
				      ,input [31:0] rd_req_desc_8_axuser_4_reg
				      ,input [31:0] rd_req_desc_8_axuser_5_reg
				      ,input [31:0] rd_req_desc_8_axuser_6_reg
				      ,input [31:0] rd_req_desc_8_axuser_7_reg
				      ,input [31:0] rd_req_desc_8_axuser_8_reg
				      ,input [31:0] rd_req_desc_8_axuser_9_reg
				      ,input [31:0] rd_req_desc_8_axuser_10_reg
				      ,input [31:0] rd_req_desc_8_axuser_11_reg
				      ,input [31:0] rd_req_desc_8_axuser_12_reg
				      ,input [31:0] rd_req_desc_8_axuser_13_reg
				      ,input [31:0] rd_req_desc_8_axuser_14_reg
				      ,input [31:0] rd_req_desc_8_axuser_15_reg
				      ,input [31:0] rd_resp_desc_8_data_offset_reg
				      ,input [31:0] rd_resp_desc_8_data_size_reg
				      ,input [31:0] rd_resp_desc_8_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_8_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_8_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_8_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_8_resp_reg
				      ,input [31:0] rd_resp_desc_8_xid_0_reg
				      ,input [31:0] rd_resp_desc_8_xid_1_reg
				      ,input [31:0] rd_resp_desc_8_xid_2_reg
				      ,input [31:0] rd_resp_desc_8_xid_3_reg
				      ,input [31:0] rd_resp_desc_8_xuser_0_reg
				      ,input [31:0] rd_resp_desc_8_xuser_1_reg
				      ,input [31:0] rd_resp_desc_8_xuser_2_reg
				      ,input [31:0] rd_resp_desc_8_xuser_3_reg
				      ,input [31:0] rd_resp_desc_8_xuser_4_reg
				      ,input [31:0] rd_resp_desc_8_xuser_5_reg
				      ,input [31:0] rd_resp_desc_8_xuser_6_reg
				      ,input [31:0] rd_resp_desc_8_xuser_7_reg
				      ,input [31:0] rd_resp_desc_8_xuser_8_reg
				      ,input [31:0] rd_resp_desc_8_xuser_9_reg
				      ,input [31:0] rd_resp_desc_8_xuser_10_reg
				      ,input [31:0] rd_resp_desc_8_xuser_11_reg
				      ,input [31:0] rd_resp_desc_8_xuser_12_reg
				      ,input [31:0] rd_resp_desc_8_xuser_13_reg
				      ,input [31:0] rd_resp_desc_8_xuser_14_reg
				      ,input [31:0] rd_resp_desc_8_xuser_15_reg
				      ,input [31:0] wr_req_desc_8_txn_type_reg
				      ,input [31:0] wr_req_desc_8_size_reg
				      ,input [31:0] wr_req_desc_8_data_offset_reg
				      ,input [31:0] wr_req_desc_8_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_8_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_8_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_8_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_8_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_8_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_8_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_8_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_8_axsize_reg
				      ,input [31:0] wr_req_desc_8_attr_reg
				      ,input [31:0] wr_req_desc_8_axaddr_0_reg
				      ,input [31:0] wr_req_desc_8_axaddr_1_reg
				      ,input [31:0] wr_req_desc_8_axaddr_2_reg
				      ,input [31:0] wr_req_desc_8_axaddr_3_reg
				      ,input [31:0] wr_req_desc_8_axid_0_reg
				      ,input [31:0] wr_req_desc_8_axid_1_reg
				      ,input [31:0] wr_req_desc_8_axid_2_reg
				      ,input [31:0] wr_req_desc_8_axid_3_reg
				      ,input [31:0] wr_req_desc_8_axuser_0_reg
				      ,input [31:0] wr_req_desc_8_axuser_1_reg
				      ,input [31:0] wr_req_desc_8_axuser_2_reg
				      ,input [31:0] wr_req_desc_8_axuser_3_reg
				      ,input [31:0] wr_req_desc_8_axuser_4_reg
				      ,input [31:0] wr_req_desc_8_axuser_5_reg
				      ,input [31:0] wr_req_desc_8_axuser_6_reg
				      ,input [31:0] wr_req_desc_8_axuser_7_reg
				      ,input [31:0] wr_req_desc_8_axuser_8_reg
				      ,input [31:0] wr_req_desc_8_axuser_9_reg
				      ,input [31:0] wr_req_desc_8_axuser_10_reg
				      ,input [31:0] wr_req_desc_8_axuser_11_reg
				      ,input [31:0] wr_req_desc_8_axuser_12_reg
				      ,input [31:0] wr_req_desc_8_axuser_13_reg
				      ,input [31:0] wr_req_desc_8_axuser_14_reg
				      ,input [31:0] wr_req_desc_8_axuser_15_reg
				      ,input [31:0] wr_req_desc_8_wuser_0_reg
				      ,input [31:0] wr_req_desc_8_wuser_1_reg
				      ,input [31:0] wr_req_desc_8_wuser_2_reg
				      ,input [31:0] wr_req_desc_8_wuser_3_reg
				      ,input [31:0] wr_req_desc_8_wuser_4_reg
				      ,input [31:0] wr_req_desc_8_wuser_5_reg
				      ,input [31:0] wr_req_desc_8_wuser_6_reg
				      ,input [31:0] wr_req_desc_8_wuser_7_reg
				      ,input [31:0] wr_req_desc_8_wuser_8_reg
				      ,input [31:0] wr_req_desc_8_wuser_9_reg
				      ,input [31:0] wr_req_desc_8_wuser_10_reg
				      ,input [31:0] wr_req_desc_8_wuser_11_reg
				      ,input [31:0] wr_req_desc_8_wuser_12_reg
				      ,input [31:0] wr_req_desc_8_wuser_13_reg
				      ,input [31:0] wr_req_desc_8_wuser_14_reg
				      ,input [31:0] wr_req_desc_8_wuser_15_reg
				      ,input [31:0] wr_resp_desc_8_resp_reg
				      ,input [31:0] wr_resp_desc_8_xid_0_reg
				      ,input [31:0] wr_resp_desc_8_xid_1_reg
				      ,input [31:0] wr_resp_desc_8_xid_2_reg
				      ,input [31:0] wr_resp_desc_8_xid_3_reg
				      ,input [31:0] wr_resp_desc_8_xuser_0_reg
				      ,input [31:0] wr_resp_desc_8_xuser_1_reg
				      ,input [31:0] wr_resp_desc_8_xuser_2_reg
				      ,input [31:0] wr_resp_desc_8_xuser_3_reg
				      ,input [31:0] wr_resp_desc_8_xuser_4_reg
				      ,input [31:0] wr_resp_desc_8_xuser_5_reg
				      ,input [31:0] wr_resp_desc_8_xuser_6_reg
				      ,input [31:0] wr_resp_desc_8_xuser_7_reg
				      ,input [31:0] wr_resp_desc_8_xuser_8_reg
				      ,input [31:0] wr_resp_desc_8_xuser_9_reg
				      ,input [31:0] wr_resp_desc_8_xuser_10_reg
				      ,input [31:0] wr_resp_desc_8_xuser_11_reg
				      ,input [31:0] wr_resp_desc_8_xuser_12_reg
				      ,input [31:0] wr_resp_desc_8_xuser_13_reg
				      ,input [31:0] wr_resp_desc_8_xuser_14_reg
				      ,input [31:0] wr_resp_desc_8_xuser_15_reg
				      ,input [31:0] sn_req_desc_8_attr_reg
				      ,input [31:0] sn_req_desc_8_acaddr_0_reg
				      ,input [31:0] sn_req_desc_8_acaddr_1_reg
				      ,input [31:0] sn_req_desc_8_acaddr_2_reg
				      ,input [31:0] sn_req_desc_8_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_8_resp_reg
				      ,input [31:0] rd_req_desc_9_txn_type_reg
				      ,input [31:0] rd_req_desc_9_size_reg
				      ,input [31:0] rd_req_desc_9_axsize_reg
				      ,input [31:0] rd_req_desc_9_attr_reg
				      ,input [31:0] rd_req_desc_9_axaddr_0_reg
				      ,input [31:0] rd_req_desc_9_axaddr_1_reg
				      ,input [31:0] rd_req_desc_9_axaddr_2_reg
				      ,input [31:0] rd_req_desc_9_axaddr_3_reg
				      ,input [31:0] rd_req_desc_9_axid_0_reg
				      ,input [31:0] rd_req_desc_9_axid_1_reg
				      ,input [31:0] rd_req_desc_9_axid_2_reg
				      ,input [31:0] rd_req_desc_9_axid_3_reg
				      ,input [31:0] rd_req_desc_9_axuser_0_reg
				      ,input [31:0] rd_req_desc_9_axuser_1_reg
				      ,input [31:0] rd_req_desc_9_axuser_2_reg
				      ,input [31:0] rd_req_desc_9_axuser_3_reg
				      ,input [31:0] rd_req_desc_9_axuser_4_reg
				      ,input [31:0] rd_req_desc_9_axuser_5_reg
				      ,input [31:0] rd_req_desc_9_axuser_6_reg
				      ,input [31:0] rd_req_desc_9_axuser_7_reg
				      ,input [31:0] rd_req_desc_9_axuser_8_reg
				      ,input [31:0] rd_req_desc_9_axuser_9_reg
				      ,input [31:0] rd_req_desc_9_axuser_10_reg
				      ,input [31:0] rd_req_desc_9_axuser_11_reg
				      ,input [31:0] rd_req_desc_9_axuser_12_reg
				      ,input [31:0] rd_req_desc_9_axuser_13_reg
				      ,input [31:0] rd_req_desc_9_axuser_14_reg
				      ,input [31:0] rd_req_desc_9_axuser_15_reg
				      ,input [31:0] rd_resp_desc_9_data_offset_reg
				      ,input [31:0] rd_resp_desc_9_data_size_reg
				      ,input [31:0] rd_resp_desc_9_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_9_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_9_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_9_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_9_resp_reg
				      ,input [31:0] rd_resp_desc_9_xid_0_reg
				      ,input [31:0] rd_resp_desc_9_xid_1_reg
				      ,input [31:0] rd_resp_desc_9_xid_2_reg
				      ,input [31:0] rd_resp_desc_9_xid_3_reg
				      ,input [31:0] rd_resp_desc_9_xuser_0_reg
				      ,input [31:0] rd_resp_desc_9_xuser_1_reg
				      ,input [31:0] rd_resp_desc_9_xuser_2_reg
				      ,input [31:0] rd_resp_desc_9_xuser_3_reg
				      ,input [31:0] rd_resp_desc_9_xuser_4_reg
				      ,input [31:0] rd_resp_desc_9_xuser_5_reg
				      ,input [31:0] rd_resp_desc_9_xuser_6_reg
				      ,input [31:0] rd_resp_desc_9_xuser_7_reg
				      ,input [31:0] rd_resp_desc_9_xuser_8_reg
				      ,input [31:0] rd_resp_desc_9_xuser_9_reg
				      ,input [31:0] rd_resp_desc_9_xuser_10_reg
				      ,input [31:0] rd_resp_desc_9_xuser_11_reg
				      ,input [31:0] rd_resp_desc_9_xuser_12_reg
				      ,input [31:0] rd_resp_desc_9_xuser_13_reg
				      ,input [31:0] rd_resp_desc_9_xuser_14_reg
				      ,input [31:0] rd_resp_desc_9_xuser_15_reg
				      ,input [31:0] wr_req_desc_9_txn_type_reg
				      ,input [31:0] wr_req_desc_9_size_reg
				      ,input [31:0] wr_req_desc_9_data_offset_reg
				      ,input [31:0] wr_req_desc_9_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_9_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_9_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_9_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_9_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_9_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_9_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_9_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_9_axsize_reg
				      ,input [31:0] wr_req_desc_9_attr_reg
				      ,input [31:0] wr_req_desc_9_axaddr_0_reg
				      ,input [31:0] wr_req_desc_9_axaddr_1_reg
				      ,input [31:0] wr_req_desc_9_axaddr_2_reg
				      ,input [31:0] wr_req_desc_9_axaddr_3_reg
				      ,input [31:0] wr_req_desc_9_axid_0_reg
				      ,input [31:0] wr_req_desc_9_axid_1_reg
				      ,input [31:0] wr_req_desc_9_axid_2_reg
				      ,input [31:0] wr_req_desc_9_axid_3_reg
				      ,input [31:0] wr_req_desc_9_axuser_0_reg
				      ,input [31:0] wr_req_desc_9_axuser_1_reg
				      ,input [31:0] wr_req_desc_9_axuser_2_reg
				      ,input [31:0] wr_req_desc_9_axuser_3_reg
				      ,input [31:0] wr_req_desc_9_axuser_4_reg
				      ,input [31:0] wr_req_desc_9_axuser_5_reg
				      ,input [31:0] wr_req_desc_9_axuser_6_reg
				      ,input [31:0] wr_req_desc_9_axuser_7_reg
				      ,input [31:0] wr_req_desc_9_axuser_8_reg
				      ,input [31:0] wr_req_desc_9_axuser_9_reg
				      ,input [31:0] wr_req_desc_9_axuser_10_reg
				      ,input [31:0] wr_req_desc_9_axuser_11_reg
				      ,input [31:0] wr_req_desc_9_axuser_12_reg
				      ,input [31:0] wr_req_desc_9_axuser_13_reg
				      ,input [31:0] wr_req_desc_9_axuser_14_reg
				      ,input [31:0] wr_req_desc_9_axuser_15_reg
				      ,input [31:0] wr_req_desc_9_wuser_0_reg
				      ,input [31:0] wr_req_desc_9_wuser_1_reg
				      ,input [31:0] wr_req_desc_9_wuser_2_reg
				      ,input [31:0] wr_req_desc_9_wuser_3_reg
				      ,input [31:0] wr_req_desc_9_wuser_4_reg
				      ,input [31:0] wr_req_desc_9_wuser_5_reg
				      ,input [31:0] wr_req_desc_9_wuser_6_reg
				      ,input [31:0] wr_req_desc_9_wuser_7_reg
				      ,input [31:0] wr_req_desc_9_wuser_8_reg
				      ,input [31:0] wr_req_desc_9_wuser_9_reg
				      ,input [31:0] wr_req_desc_9_wuser_10_reg
				      ,input [31:0] wr_req_desc_9_wuser_11_reg
				      ,input [31:0] wr_req_desc_9_wuser_12_reg
				      ,input [31:0] wr_req_desc_9_wuser_13_reg
				      ,input [31:0] wr_req_desc_9_wuser_14_reg
				      ,input [31:0] wr_req_desc_9_wuser_15_reg
				      ,input [31:0] wr_resp_desc_9_resp_reg
				      ,input [31:0] wr_resp_desc_9_xid_0_reg
				      ,input [31:0] wr_resp_desc_9_xid_1_reg
				      ,input [31:0] wr_resp_desc_9_xid_2_reg
				      ,input [31:0] wr_resp_desc_9_xid_3_reg
				      ,input [31:0] wr_resp_desc_9_xuser_0_reg
				      ,input [31:0] wr_resp_desc_9_xuser_1_reg
				      ,input [31:0] wr_resp_desc_9_xuser_2_reg
				      ,input [31:0] wr_resp_desc_9_xuser_3_reg
				      ,input [31:0] wr_resp_desc_9_xuser_4_reg
				      ,input [31:0] wr_resp_desc_9_xuser_5_reg
				      ,input [31:0] wr_resp_desc_9_xuser_6_reg
				      ,input [31:0] wr_resp_desc_9_xuser_7_reg
				      ,input [31:0] wr_resp_desc_9_xuser_8_reg
				      ,input [31:0] wr_resp_desc_9_xuser_9_reg
				      ,input [31:0] wr_resp_desc_9_xuser_10_reg
				      ,input [31:0] wr_resp_desc_9_xuser_11_reg
				      ,input [31:0] wr_resp_desc_9_xuser_12_reg
				      ,input [31:0] wr_resp_desc_9_xuser_13_reg
				      ,input [31:0] wr_resp_desc_9_xuser_14_reg
				      ,input [31:0] wr_resp_desc_9_xuser_15_reg
				      ,input [31:0] sn_req_desc_9_attr_reg
				      ,input [31:0] sn_req_desc_9_acaddr_0_reg
				      ,input [31:0] sn_req_desc_9_acaddr_1_reg
				      ,input [31:0] sn_req_desc_9_acaddr_2_reg
				      ,input [31:0] sn_req_desc_9_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_9_resp_reg
				      ,input [31:0] rd_req_desc_a_txn_type_reg
				      ,input [31:0] rd_req_desc_a_size_reg
				      ,input [31:0] rd_req_desc_a_axsize_reg
				      ,input [31:0] rd_req_desc_a_attr_reg
				      ,input [31:0] rd_req_desc_a_axaddr_0_reg
				      ,input [31:0] rd_req_desc_a_axaddr_1_reg
				      ,input [31:0] rd_req_desc_a_axaddr_2_reg
				      ,input [31:0] rd_req_desc_a_axaddr_3_reg
				      ,input [31:0] rd_req_desc_a_axid_0_reg
				      ,input [31:0] rd_req_desc_a_axid_1_reg
				      ,input [31:0] rd_req_desc_a_axid_2_reg
				      ,input [31:0] rd_req_desc_a_axid_3_reg
				      ,input [31:0] rd_req_desc_a_axuser_0_reg
				      ,input [31:0] rd_req_desc_a_axuser_1_reg
				      ,input [31:0] rd_req_desc_a_axuser_2_reg
				      ,input [31:0] rd_req_desc_a_axuser_3_reg
				      ,input [31:0] rd_req_desc_a_axuser_4_reg
				      ,input [31:0] rd_req_desc_a_axuser_5_reg
				      ,input [31:0] rd_req_desc_a_axuser_6_reg
				      ,input [31:0] rd_req_desc_a_axuser_7_reg
				      ,input [31:0] rd_req_desc_a_axuser_8_reg
				      ,input [31:0] rd_req_desc_a_axuser_9_reg
				      ,input [31:0] rd_req_desc_a_axuser_10_reg
				      ,input [31:0] rd_req_desc_a_axuser_11_reg
				      ,input [31:0] rd_req_desc_a_axuser_12_reg
				      ,input [31:0] rd_req_desc_a_axuser_13_reg
				      ,input [31:0] rd_req_desc_a_axuser_14_reg
				      ,input [31:0] rd_req_desc_a_axuser_15_reg
				      ,input [31:0] rd_resp_desc_a_data_offset_reg
				      ,input [31:0] rd_resp_desc_a_data_size_reg
				      ,input [31:0] rd_resp_desc_a_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_a_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_a_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_a_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_a_resp_reg
				      ,input [31:0] rd_resp_desc_a_xid_0_reg
				      ,input [31:0] rd_resp_desc_a_xid_1_reg
				      ,input [31:0] rd_resp_desc_a_xid_2_reg
				      ,input [31:0] rd_resp_desc_a_xid_3_reg
				      ,input [31:0] rd_resp_desc_a_xuser_0_reg
				      ,input [31:0] rd_resp_desc_a_xuser_1_reg
				      ,input [31:0] rd_resp_desc_a_xuser_2_reg
				      ,input [31:0] rd_resp_desc_a_xuser_3_reg
				      ,input [31:0] rd_resp_desc_a_xuser_4_reg
				      ,input [31:0] rd_resp_desc_a_xuser_5_reg
				      ,input [31:0] rd_resp_desc_a_xuser_6_reg
				      ,input [31:0] rd_resp_desc_a_xuser_7_reg
				      ,input [31:0] rd_resp_desc_a_xuser_8_reg
				      ,input [31:0] rd_resp_desc_a_xuser_9_reg
				      ,input [31:0] rd_resp_desc_a_xuser_10_reg
				      ,input [31:0] rd_resp_desc_a_xuser_11_reg
				      ,input [31:0] rd_resp_desc_a_xuser_12_reg
				      ,input [31:0] rd_resp_desc_a_xuser_13_reg
				      ,input [31:0] rd_resp_desc_a_xuser_14_reg
				      ,input [31:0] rd_resp_desc_a_xuser_15_reg
				      ,input [31:0] wr_req_desc_a_txn_type_reg
				      ,input [31:0] wr_req_desc_a_size_reg
				      ,input [31:0] wr_req_desc_a_data_offset_reg
				      ,input [31:0] wr_req_desc_a_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_a_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_a_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_a_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_a_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_a_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_a_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_a_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_a_axsize_reg
				      ,input [31:0] wr_req_desc_a_attr_reg
				      ,input [31:0] wr_req_desc_a_axaddr_0_reg
				      ,input [31:0] wr_req_desc_a_axaddr_1_reg
				      ,input [31:0] wr_req_desc_a_axaddr_2_reg
				      ,input [31:0] wr_req_desc_a_axaddr_3_reg
				      ,input [31:0] wr_req_desc_a_axid_0_reg
				      ,input [31:0] wr_req_desc_a_axid_1_reg
				      ,input [31:0] wr_req_desc_a_axid_2_reg
				      ,input [31:0] wr_req_desc_a_axid_3_reg
				      ,input [31:0] wr_req_desc_a_axuser_0_reg
				      ,input [31:0] wr_req_desc_a_axuser_1_reg
				      ,input [31:0] wr_req_desc_a_axuser_2_reg
				      ,input [31:0] wr_req_desc_a_axuser_3_reg
				      ,input [31:0] wr_req_desc_a_axuser_4_reg
				      ,input [31:0] wr_req_desc_a_axuser_5_reg
				      ,input [31:0] wr_req_desc_a_axuser_6_reg
				      ,input [31:0] wr_req_desc_a_axuser_7_reg
				      ,input [31:0] wr_req_desc_a_axuser_8_reg
				      ,input [31:0] wr_req_desc_a_axuser_9_reg
				      ,input [31:0] wr_req_desc_a_axuser_10_reg
				      ,input [31:0] wr_req_desc_a_axuser_11_reg
				      ,input [31:0] wr_req_desc_a_axuser_12_reg
				      ,input [31:0] wr_req_desc_a_axuser_13_reg
				      ,input [31:0] wr_req_desc_a_axuser_14_reg
				      ,input [31:0] wr_req_desc_a_axuser_15_reg
				      ,input [31:0] wr_req_desc_a_wuser_0_reg
				      ,input [31:0] wr_req_desc_a_wuser_1_reg
				      ,input [31:0] wr_req_desc_a_wuser_2_reg
				      ,input [31:0] wr_req_desc_a_wuser_3_reg
				      ,input [31:0] wr_req_desc_a_wuser_4_reg
				      ,input [31:0] wr_req_desc_a_wuser_5_reg
				      ,input [31:0] wr_req_desc_a_wuser_6_reg
				      ,input [31:0] wr_req_desc_a_wuser_7_reg
				      ,input [31:0] wr_req_desc_a_wuser_8_reg
				      ,input [31:0] wr_req_desc_a_wuser_9_reg
				      ,input [31:0] wr_req_desc_a_wuser_10_reg
				      ,input [31:0] wr_req_desc_a_wuser_11_reg
				      ,input [31:0] wr_req_desc_a_wuser_12_reg
				      ,input [31:0] wr_req_desc_a_wuser_13_reg
				      ,input [31:0] wr_req_desc_a_wuser_14_reg
				      ,input [31:0] wr_req_desc_a_wuser_15_reg
				      ,input [31:0] wr_resp_desc_a_resp_reg
				      ,input [31:0] wr_resp_desc_a_xid_0_reg
				      ,input [31:0] wr_resp_desc_a_xid_1_reg
				      ,input [31:0] wr_resp_desc_a_xid_2_reg
				      ,input [31:0] wr_resp_desc_a_xid_3_reg
				      ,input [31:0] wr_resp_desc_a_xuser_0_reg
				      ,input [31:0] wr_resp_desc_a_xuser_1_reg
				      ,input [31:0] wr_resp_desc_a_xuser_2_reg
				      ,input [31:0] wr_resp_desc_a_xuser_3_reg
				      ,input [31:0] wr_resp_desc_a_xuser_4_reg
				      ,input [31:0] wr_resp_desc_a_xuser_5_reg
				      ,input [31:0] wr_resp_desc_a_xuser_6_reg
				      ,input [31:0] wr_resp_desc_a_xuser_7_reg
				      ,input [31:0] wr_resp_desc_a_xuser_8_reg
				      ,input [31:0] wr_resp_desc_a_xuser_9_reg
				      ,input [31:0] wr_resp_desc_a_xuser_10_reg
				      ,input [31:0] wr_resp_desc_a_xuser_11_reg
				      ,input [31:0] wr_resp_desc_a_xuser_12_reg
				      ,input [31:0] wr_resp_desc_a_xuser_13_reg
				      ,input [31:0] wr_resp_desc_a_xuser_14_reg
				      ,input [31:0] wr_resp_desc_a_xuser_15_reg
				      ,input [31:0] sn_req_desc_a_attr_reg
				      ,input [31:0] sn_req_desc_a_acaddr_0_reg
				      ,input [31:0] sn_req_desc_a_acaddr_1_reg
				      ,input [31:0] sn_req_desc_a_acaddr_2_reg
				      ,input [31:0] sn_req_desc_a_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_a_resp_reg
				      ,input [31:0] rd_req_desc_b_txn_type_reg
				      ,input [31:0] rd_req_desc_b_size_reg
				      ,input [31:0] rd_req_desc_b_axsize_reg
				      ,input [31:0] rd_req_desc_b_attr_reg
				      ,input [31:0] rd_req_desc_b_axaddr_0_reg
				      ,input [31:0] rd_req_desc_b_axaddr_1_reg
				      ,input [31:0] rd_req_desc_b_axaddr_2_reg
				      ,input [31:0] rd_req_desc_b_axaddr_3_reg
				      ,input [31:0] rd_req_desc_b_axid_0_reg
				      ,input [31:0] rd_req_desc_b_axid_1_reg
				      ,input [31:0] rd_req_desc_b_axid_2_reg
				      ,input [31:0] rd_req_desc_b_axid_3_reg
				      ,input [31:0] rd_req_desc_b_axuser_0_reg
				      ,input [31:0] rd_req_desc_b_axuser_1_reg
				      ,input [31:0] rd_req_desc_b_axuser_2_reg
				      ,input [31:0] rd_req_desc_b_axuser_3_reg
				      ,input [31:0] rd_req_desc_b_axuser_4_reg
				      ,input [31:0] rd_req_desc_b_axuser_5_reg
				      ,input [31:0] rd_req_desc_b_axuser_6_reg
				      ,input [31:0] rd_req_desc_b_axuser_7_reg
				      ,input [31:0] rd_req_desc_b_axuser_8_reg
				      ,input [31:0] rd_req_desc_b_axuser_9_reg
				      ,input [31:0] rd_req_desc_b_axuser_10_reg
				      ,input [31:0] rd_req_desc_b_axuser_11_reg
				      ,input [31:0] rd_req_desc_b_axuser_12_reg
				      ,input [31:0] rd_req_desc_b_axuser_13_reg
				      ,input [31:0] rd_req_desc_b_axuser_14_reg
				      ,input [31:0] rd_req_desc_b_axuser_15_reg
				      ,input [31:0] rd_resp_desc_b_data_offset_reg
				      ,input [31:0] rd_resp_desc_b_data_size_reg
				      ,input [31:0] rd_resp_desc_b_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_b_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_b_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_b_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_b_resp_reg
				      ,input [31:0] rd_resp_desc_b_xid_0_reg
				      ,input [31:0] rd_resp_desc_b_xid_1_reg
				      ,input [31:0] rd_resp_desc_b_xid_2_reg
				      ,input [31:0] rd_resp_desc_b_xid_3_reg
				      ,input [31:0] rd_resp_desc_b_xuser_0_reg
				      ,input [31:0] rd_resp_desc_b_xuser_1_reg
				      ,input [31:0] rd_resp_desc_b_xuser_2_reg
				      ,input [31:0] rd_resp_desc_b_xuser_3_reg
				      ,input [31:0] rd_resp_desc_b_xuser_4_reg
				      ,input [31:0] rd_resp_desc_b_xuser_5_reg
				      ,input [31:0] rd_resp_desc_b_xuser_6_reg
				      ,input [31:0] rd_resp_desc_b_xuser_7_reg
				      ,input [31:0] rd_resp_desc_b_xuser_8_reg
				      ,input [31:0] rd_resp_desc_b_xuser_9_reg
				      ,input [31:0] rd_resp_desc_b_xuser_10_reg
				      ,input [31:0] rd_resp_desc_b_xuser_11_reg
				      ,input [31:0] rd_resp_desc_b_xuser_12_reg
				      ,input [31:0] rd_resp_desc_b_xuser_13_reg
				      ,input [31:0] rd_resp_desc_b_xuser_14_reg
				      ,input [31:0] rd_resp_desc_b_xuser_15_reg
				      ,input [31:0] wr_req_desc_b_txn_type_reg
				      ,input [31:0] wr_req_desc_b_size_reg
				      ,input [31:0] wr_req_desc_b_data_offset_reg
				      ,input [31:0] wr_req_desc_b_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_b_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_b_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_b_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_b_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_b_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_b_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_b_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_b_axsize_reg
				      ,input [31:0] wr_req_desc_b_attr_reg
				      ,input [31:0] wr_req_desc_b_axaddr_0_reg
				      ,input [31:0] wr_req_desc_b_axaddr_1_reg
				      ,input [31:0] wr_req_desc_b_axaddr_2_reg
				      ,input [31:0] wr_req_desc_b_axaddr_3_reg
				      ,input [31:0] wr_req_desc_b_axid_0_reg
				      ,input [31:0] wr_req_desc_b_axid_1_reg
				      ,input [31:0] wr_req_desc_b_axid_2_reg
				      ,input [31:0] wr_req_desc_b_axid_3_reg
				      ,input [31:0] wr_req_desc_b_axuser_0_reg
				      ,input [31:0] wr_req_desc_b_axuser_1_reg
				      ,input [31:0] wr_req_desc_b_axuser_2_reg
				      ,input [31:0] wr_req_desc_b_axuser_3_reg
				      ,input [31:0] wr_req_desc_b_axuser_4_reg
				      ,input [31:0] wr_req_desc_b_axuser_5_reg
				      ,input [31:0] wr_req_desc_b_axuser_6_reg
				      ,input [31:0] wr_req_desc_b_axuser_7_reg
				      ,input [31:0] wr_req_desc_b_axuser_8_reg
				      ,input [31:0] wr_req_desc_b_axuser_9_reg
				      ,input [31:0] wr_req_desc_b_axuser_10_reg
				      ,input [31:0] wr_req_desc_b_axuser_11_reg
				      ,input [31:0] wr_req_desc_b_axuser_12_reg
				      ,input [31:0] wr_req_desc_b_axuser_13_reg
				      ,input [31:0] wr_req_desc_b_axuser_14_reg
				      ,input [31:0] wr_req_desc_b_axuser_15_reg
				      ,input [31:0] wr_req_desc_b_wuser_0_reg
				      ,input [31:0] wr_req_desc_b_wuser_1_reg
				      ,input [31:0] wr_req_desc_b_wuser_2_reg
				      ,input [31:0] wr_req_desc_b_wuser_3_reg
				      ,input [31:0] wr_req_desc_b_wuser_4_reg
				      ,input [31:0] wr_req_desc_b_wuser_5_reg
				      ,input [31:0] wr_req_desc_b_wuser_6_reg
				      ,input [31:0] wr_req_desc_b_wuser_7_reg
				      ,input [31:0] wr_req_desc_b_wuser_8_reg
				      ,input [31:0] wr_req_desc_b_wuser_9_reg
				      ,input [31:0] wr_req_desc_b_wuser_10_reg
				      ,input [31:0] wr_req_desc_b_wuser_11_reg
				      ,input [31:0] wr_req_desc_b_wuser_12_reg
				      ,input [31:0] wr_req_desc_b_wuser_13_reg
				      ,input [31:0] wr_req_desc_b_wuser_14_reg
				      ,input [31:0] wr_req_desc_b_wuser_15_reg
				      ,input [31:0] wr_resp_desc_b_resp_reg
				      ,input [31:0] wr_resp_desc_b_xid_0_reg
				      ,input [31:0] wr_resp_desc_b_xid_1_reg
				      ,input [31:0] wr_resp_desc_b_xid_2_reg
				      ,input [31:0] wr_resp_desc_b_xid_3_reg
				      ,input [31:0] wr_resp_desc_b_xuser_0_reg
				      ,input [31:0] wr_resp_desc_b_xuser_1_reg
				      ,input [31:0] wr_resp_desc_b_xuser_2_reg
				      ,input [31:0] wr_resp_desc_b_xuser_3_reg
				      ,input [31:0] wr_resp_desc_b_xuser_4_reg
				      ,input [31:0] wr_resp_desc_b_xuser_5_reg
				      ,input [31:0] wr_resp_desc_b_xuser_6_reg
				      ,input [31:0] wr_resp_desc_b_xuser_7_reg
				      ,input [31:0] wr_resp_desc_b_xuser_8_reg
				      ,input [31:0] wr_resp_desc_b_xuser_9_reg
				      ,input [31:0] wr_resp_desc_b_xuser_10_reg
				      ,input [31:0] wr_resp_desc_b_xuser_11_reg
				      ,input [31:0] wr_resp_desc_b_xuser_12_reg
				      ,input [31:0] wr_resp_desc_b_xuser_13_reg
				      ,input [31:0] wr_resp_desc_b_xuser_14_reg
				      ,input [31:0] wr_resp_desc_b_xuser_15_reg
				      ,input [31:0] sn_req_desc_b_attr_reg
				      ,input [31:0] sn_req_desc_b_acaddr_0_reg
				      ,input [31:0] sn_req_desc_b_acaddr_1_reg
				      ,input [31:0] sn_req_desc_b_acaddr_2_reg
				      ,input [31:0] sn_req_desc_b_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_b_resp_reg
				      ,input [31:0] rd_req_desc_c_txn_type_reg
				      ,input [31:0] rd_req_desc_c_size_reg
				      ,input [31:0] rd_req_desc_c_axsize_reg
				      ,input [31:0] rd_req_desc_c_attr_reg
				      ,input [31:0] rd_req_desc_c_axaddr_0_reg
				      ,input [31:0] rd_req_desc_c_axaddr_1_reg
				      ,input [31:0] rd_req_desc_c_axaddr_2_reg
				      ,input [31:0] rd_req_desc_c_axaddr_3_reg
				      ,input [31:0] rd_req_desc_c_axid_0_reg
				      ,input [31:0] rd_req_desc_c_axid_1_reg
				      ,input [31:0] rd_req_desc_c_axid_2_reg
				      ,input [31:0] rd_req_desc_c_axid_3_reg
				      ,input [31:0] rd_req_desc_c_axuser_0_reg
				      ,input [31:0] rd_req_desc_c_axuser_1_reg
				      ,input [31:0] rd_req_desc_c_axuser_2_reg
				      ,input [31:0] rd_req_desc_c_axuser_3_reg
				      ,input [31:0] rd_req_desc_c_axuser_4_reg
				      ,input [31:0] rd_req_desc_c_axuser_5_reg
				      ,input [31:0] rd_req_desc_c_axuser_6_reg
				      ,input [31:0] rd_req_desc_c_axuser_7_reg
				      ,input [31:0] rd_req_desc_c_axuser_8_reg
				      ,input [31:0] rd_req_desc_c_axuser_9_reg
				      ,input [31:0] rd_req_desc_c_axuser_10_reg
				      ,input [31:0] rd_req_desc_c_axuser_11_reg
				      ,input [31:0] rd_req_desc_c_axuser_12_reg
				      ,input [31:0] rd_req_desc_c_axuser_13_reg
				      ,input [31:0] rd_req_desc_c_axuser_14_reg
				      ,input [31:0] rd_req_desc_c_axuser_15_reg
				      ,input [31:0] rd_resp_desc_c_data_offset_reg
				      ,input [31:0] rd_resp_desc_c_data_size_reg
				      ,input [31:0] rd_resp_desc_c_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_c_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_c_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_c_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_c_resp_reg
				      ,input [31:0] rd_resp_desc_c_xid_0_reg
				      ,input [31:0] rd_resp_desc_c_xid_1_reg
				      ,input [31:0] rd_resp_desc_c_xid_2_reg
				      ,input [31:0] rd_resp_desc_c_xid_3_reg
				      ,input [31:0] rd_resp_desc_c_xuser_0_reg
				      ,input [31:0] rd_resp_desc_c_xuser_1_reg
				      ,input [31:0] rd_resp_desc_c_xuser_2_reg
				      ,input [31:0] rd_resp_desc_c_xuser_3_reg
				      ,input [31:0] rd_resp_desc_c_xuser_4_reg
				      ,input [31:0] rd_resp_desc_c_xuser_5_reg
				      ,input [31:0] rd_resp_desc_c_xuser_6_reg
				      ,input [31:0] rd_resp_desc_c_xuser_7_reg
				      ,input [31:0] rd_resp_desc_c_xuser_8_reg
				      ,input [31:0] rd_resp_desc_c_xuser_9_reg
				      ,input [31:0] rd_resp_desc_c_xuser_10_reg
				      ,input [31:0] rd_resp_desc_c_xuser_11_reg
				      ,input [31:0] rd_resp_desc_c_xuser_12_reg
				      ,input [31:0] rd_resp_desc_c_xuser_13_reg
				      ,input [31:0] rd_resp_desc_c_xuser_14_reg
				      ,input [31:0] rd_resp_desc_c_xuser_15_reg
				      ,input [31:0] wr_req_desc_c_txn_type_reg
				      ,input [31:0] wr_req_desc_c_size_reg
				      ,input [31:0] wr_req_desc_c_data_offset_reg
				      ,input [31:0] wr_req_desc_c_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_c_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_c_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_c_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_c_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_c_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_c_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_c_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_c_axsize_reg
				      ,input [31:0] wr_req_desc_c_attr_reg
				      ,input [31:0] wr_req_desc_c_axaddr_0_reg
				      ,input [31:0] wr_req_desc_c_axaddr_1_reg
				      ,input [31:0] wr_req_desc_c_axaddr_2_reg
				      ,input [31:0] wr_req_desc_c_axaddr_3_reg
				      ,input [31:0] wr_req_desc_c_axid_0_reg
				      ,input [31:0] wr_req_desc_c_axid_1_reg
				      ,input [31:0] wr_req_desc_c_axid_2_reg
				      ,input [31:0] wr_req_desc_c_axid_3_reg
				      ,input [31:0] wr_req_desc_c_axuser_0_reg
				      ,input [31:0] wr_req_desc_c_axuser_1_reg
				      ,input [31:0] wr_req_desc_c_axuser_2_reg
				      ,input [31:0] wr_req_desc_c_axuser_3_reg
				      ,input [31:0] wr_req_desc_c_axuser_4_reg
				      ,input [31:0] wr_req_desc_c_axuser_5_reg
				      ,input [31:0] wr_req_desc_c_axuser_6_reg
				      ,input [31:0] wr_req_desc_c_axuser_7_reg
				      ,input [31:0] wr_req_desc_c_axuser_8_reg
				      ,input [31:0] wr_req_desc_c_axuser_9_reg
				      ,input [31:0] wr_req_desc_c_axuser_10_reg
				      ,input [31:0] wr_req_desc_c_axuser_11_reg
				      ,input [31:0] wr_req_desc_c_axuser_12_reg
				      ,input [31:0] wr_req_desc_c_axuser_13_reg
				      ,input [31:0] wr_req_desc_c_axuser_14_reg
				      ,input [31:0] wr_req_desc_c_axuser_15_reg
				      ,input [31:0] wr_req_desc_c_wuser_0_reg
				      ,input [31:0] wr_req_desc_c_wuser_1_reg
				      ,input [31:0] wr_req_desc_c_wuser_2_reg
				      ,input [31:0] wr_req_desc_c_wuser_3_reg
				      ,input [31:0] wr_req_desc_c_wuser_4_reg
				      ,input [31:0] wr_req_desc_c_wuser_5_reg
				      ,input [31:0] wr_req_desc_c_wuser_6_reg
				      ,input [31:0] wr_req_desc_c_wuser_7_reg
				      ,input [31:0] wr_req_desc_c_wuser_8_reg
				      ,input [31:0] wr_req_desc_c_wuser_9_reg
				      ,input [31:0] wr_req_desc_c_wuser_10_reg
				      ,input [31:0] wr_req_desc_c_wuser_11_reg
				      ,input [31:0] wr_req_desc_c_wuser_12_reg
				      ,input [31:0] wr_req_desc_c_wuser_13_reg
				      ,input [31:0] wr_req_desc_c_wuser_14_reg
				      ,input [31:0] wr_req_desc_c_wuser_15_reg
				      ,input [31:0] wr_resp_desc_c_resp_reg
				      ,input [31:0] wr_resp_desc_c_xid_0_reg
				      ,input [31:0] wr_resp_desc_c_xid_1_reg
				      ,input [31:0] wr_resp_desc_c_xid_2_reg
				      ,input [31:0] wr_resp_desc_c_xid_3_reg
				      ,input [31:0] wr_resp_desc_c_xuser_0_reg
				      ,input [31:0] wr_resp_desc_c_xuser_1_reg
				      ,input [31:0] wr_resp_desc_c_xuser_2_reg
				      ,input [31:0] wr_resp_desc_c_xuser_3_reg
				      ,input [31:0] wr_resp_desc_c_xuser_4_reg
				      ,input [31:0] wr_resp_desc_c_xuser_5_reg
				      ,input [31:0] wr_resp_desc_c_xuser_6_reg
				      ,input [31:0] wr_resp_desc_c_xuser_7_reg
				      ,input [31:0] wr_resp_desc_c_xuser_8_reg
				      ,input [31:0] wr_resp_desc_c_xuser_9_reg
				      ,input [31:0] wr_resp_desc_c_xuser_10_reg
				      ,input [31:0] wr_resp_desc_c_xuser_11_reg
				      ,input [31:0] wr_resp_desc_c_xuser_12_reg
				      ,input [31:0] wr_resp_desc_c_xuser_13_reg
				      ,input [31:0] wr_resp_desc_c_xuser_14_reg
				      ,input [31:0] wr_resp_desc_c_xuser_15_reg
				      ,input [31:0] sn_req_desc_c_attr_reg
				      ,input [31:0] sn_req_desc_c_acaddr_0_reg
				      ,input [31:0] sn_req_desc_c_acaddr_1_reg
				      ,input [31:0] sn_req_desc_c_acaddr_2_reg
				      ,input [31:0] sn_req_desc_c_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_c_resp_reg
				      ,input [31:0] rd_req_desc_d_txn_type_reg
				      ,input [31:0] rd_req_desc_d_size_reg
				      ,input [31:0] rd_req_desc_d_axsize_reg
				      ,input [31:0] rd_req_desc_d_attr_reg
				      ,input [31:0] rd_req_desc_d_axaddr_0_reg
				      ,input [31:0] rd_req_desc_d_axaddr_1_reg
				      ,input [31:0] rd_req_desc_d_axaddr_2_reg
				      ,input [31:0] rd_req_desc_d_axaddr_3_reg
				      ,input [31:0] rd_req_desc_d_axid_0_reg
				      ,input [31:0] rd_req_desc_d_axid_1_reg
				      ,input [31:0] rd_req_desc_d_axid_2_reg
				      ,input [31:0] rd_req_desc_d_axid_3_reg
				      ,input [31:0] rd_req_desc_d_axuser_0_reg
				      ,input [31:0] rd_req_desc_d_axuser_1_reg
				      ,input [31:0] rd_req_desc_d_axuser_2_reg
				      ,input [31:0] rd_req_desc_d_axuser_3_reg
				      ,input [31:0] rd_req_desc_d_axuser_4_reg
				      ,input [31:0] rd_req_desc_d_axuser_5_reg
				      ,input [31:0] rd_req_desc_d_axuser_6_reg
				      ,input [31:0] rd_req_desc_d_axuser_7_reg
				      ,input [31:0] rd_req_desc_d_axuser_8_reg
				      ,input [31:0] rd_req_desc_d_axuser_9_reg
				      ,input [31:0] rd_req_desc_d_axuser_10_reg
				      ,input [31:0] rd_req_desc_d_axuser_11_reg
				      ,input [31:0] rd_req_desc_d_axuser_12_reg
				      ,input [31:0] rd_req_desc_d_axuser_13_reg
				      ,input [31:0] rd_req_desc_d_axuser_14_reg
				      ,input [31:0] rd_req_desc_d_axuser_15_reg
				      ,input [31:0] rd_resp_desc_d_data_offset_reg
				      ,input [31:0] rd_resp_desc_d_data_size_reg
				      ,input [31:0] rd_resp_desc_d_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_d_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_d_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_d_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_d_resp_reg
				      ,input [31:0] rd_resp_desc_d_xid_0_reg
				      ,input [31:0] rd_resp_desc_d_xid_1_reg
				      ,input [31:0] rd_resp_desc_d_xid_2_reg
				      ,input [31:0] rd_resp_desc_d_xid_3_reg
				      ,input [31:0] rd_resp_desc_d_xuser_0_reg
				      ,input [31:0] rd_resp_desc_d_xuser_1_reg
				      ,input [31:0] rd_resp_desc_d_xuser_2_reg
				      ,input [31:0] rd_resp_desc_d_xuser_3_reg
				      ,input [31:0] rd_resp_desc_d_xuser_4_reg
				      ,input [31:0] rd_resp_desc_d_xuser_5_reg
				      ,input [31:0] rd_resp_desc_d_xuser_6_reg
				      ,input [31:0] rd_resp_desc_d_xuser_7_reg
				      ,input [31:0] rd_resp_desc_d_xuser_8_reg
				      ,input [31:0] rd_resp_desc_d_xuser_9_reg
				      ,input [31:0] rd_resp_desc_d_xuser_10_reg
				      ,input [31:0] rd_resp_desc_d_xuser_11_reg
				      ,input [31:0] rd_resp_desc_d_xuser_12_reg
				      ,input [31:0] rd_resp_desc_d_xuser_13_reg
				      ,input [31:0] rd_resp_desc_d_xuser_14_reg
				      ,input [31:0] rd_resp_desc_d_xuser_15_reg
				      ,input [31:0] wr_req_desc_d_txn_type_reg
				      ,input [31:0] wr_req_desc_d_size_reg
				      ,input [31:0] wr_req_desc_d_data_offset_reg
				      ,input [31:0] wr_req_desc_d_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_d_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_d_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_d_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_d_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_d_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_d_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_d_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_d_axsize_reg
				      ,input [31:0] wr_req_desc_d_attr_reg
				      ,input [31:0] wr_req_desc_d_axaddr_0_reg
				      ,input [31:0] wr_req_desc_d_axaddr_1_reg
				      ,input [31:0] wr_req_desc_d_axaddr_2_reg
				      ,input [31:0] wr_req_desc_d_axaddr_3_reg
				      ,input [31:0] wr_req_desc_d_axid_0_reg
				      ,input [31:0] wr_req_desc_d_axid_1_reg
				      ,input [31:0] wr_req_desc_d_axid_2_reg
				      ,input [31:0] wr_req_desc_d_axid_3_reg
				      ,input [31:0] wr_req_desc_d_axuser_0_reg
				      ,input [31:0] wr_req_desc_d_axuser_1_reg
				      ,input [31:0] wr_req_desc_d_axuser_2_reg
				      ,input [31:0] wr_req_desc_d_axuser_3_reg
				      ,input [31:0] wr_req_desc_d_axuser_4_reg
				      ,input [31:0] wr_req_desc_d_axuser_5_reg
				      ,input [31:0] wr_req_desc_d_axuser_6_reg
				      ,input [31:0] wr_req_desc_d_axuser_7_reg
				      ,input [31:0] wr_req_desc_d_axuser_8_reg
				      ,input [31:0] wr_req_desc_d_axuser_9_reg
				      ,input [31:0] wr_req_desc_d_axuser_10_reg
				      ,input [31:0] wr_req_desc_d_axuser_11_reg
				      ,input [31:0] wr_req_desc_d_axuser_12_reg
				      ,input [31:0] wr_req_desc_d_axuser_13_reg
				      ,input [31:0] wr_req_desc_d_axuser_14_reg
				      ,input [31:0] wr_req_desc_d_axuser_15_reg
				      ,input [31:0] wr_req_desc_d_wuser_0_reg
				      ,input [31:0] wr_req_desc_d_wuser_1_reg
				      ,input [31:0] wr_req_desc_d_wuser_2_reg
				      ,input [31:0] wr_req_desc_d_wuser_3_reg
				      ,input [31:0] wr_req_desc_d_wuser_4_reg
				      ,input [31:0] wr_req_desc_d_wuser_5_reg
				      ,input [31:0] wr_req_desc_d_wuser_6_reg
				      ,input [31:0] wr_req_desc_d_wuser_7_reg
				      ,input [31:0] wr_req_desc_d_wuser_8_reg
				      ,input [31:0] wr_req_desc_d_wuser_9_reg
				      ,input [31:0] wr_req_desc_d_wuser_10_reg
				      ,input [31:0] wr_req_desc_d_wuser_11_reg
				      ,input [31:0] wr_req_desc_d_wuser_12_reg
				      ,input [31:0] wr_req_desc_d_wuser_13_reg
				      ,input [31:0] wr_req_desc_d_wuser_14_reg
				      ,input [31:0] wr_req_desc_d_wuser_15_reg
				      ,input [31:0] wr_resp_desc_d_resp_reg
				      ,input [31:0] wr_resp_desc_d_xid_0_reg
				      ,input [31:0] wr_resp_desc_d_xid_1_reg
				      ,input [31:0] wr_resp_desc_d_xid_2_reg
				      ,input [31:0] wr_resp_desc_d_xid_3_reg
				      ,input [31:0] wr_resp_desc_d_xuser_0_reg
				      ,input [31:0] wr_resp_desc_d_xuser_1_reg
				      ,input [31:0] wr_resp_desc_d_xuser_2_reg
				      ,input [31:0] wr_resp_desc_d_xuser_3_reg
				      ,input [31:0] wr_resp_desc_d_xuser_4_reg
				      ,input [31:0] wr_resp_desc_d_xuser_5_reg
				      ,input [31:0] wr_resp_desc_d_xuser_6_reg
				      ,input [31:0] wr_resp_desc_d_xuser_7_reg
				      ,input [31:0] wr_resp_desc_d_xuser_8_reg
				      ,input [31:0] wr_resp_desc_d_xuser_9_reg
				      ,input [31:0] wr_resp_desc_d_xuser_10_reg
				      ,input [31:0] wr_resp_desc_d_xuser_11_reg
				      ,input [31:0] wr_resp_desc_d_xuser_12_reg
				      ,input [31:0] wr_resp_desc_d_xuser_13_reg
				      ,input [31:0] wr_resp_desc_d_xuser_14_reg
				      ,input [31:0] wr_resp_desc_d_xuser_15_reg
				      ,input [31:0] sn_req_desc_d_attr_reg
				      ,input [31:0] sn_req_desc_d_acaddr_0_reg
				      ,input [31:0] sn_req_desc_d_acaddr_1_reg
				      ,input [31:0] sn_req_desc_d_acaddr_2_reg
				      ,input [31:0] sn_req_desc_d_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_d_resp_reg
				      ,input [31:0] rd_req_desc_e_txn_type_reg
				      ,input [31:0] rd_req_desc_e_size_reg
				      ,input [31:0] rd_req_desc_e_axsize_reg
				      ,input [31:0] rd_req_desc_e_attr_reg
				      ,input [31:0] rd_req_desc_e_axaddr_0_reg
				      ,input [31:0] rd_req_desc_e_axaddr_1_reg
				      ,input [31:0] rd_req_desc_e_axaddr_2_reg
				      ,input [31:0] rd_req_desc_e_axaddr_3_reg
				      ,input [31:0] rd_req_desc_e_axid_0_reg
				      ,input [31:0] rd_req_desc_e_axid_1_reg
				      ,input [31:0] rd_req_desc_e_axid_2_reg
				      ,input [31:0] rd_req_desc_e_axid_3_reg
				      ,input [31:0] rd_req_desc_e_axuser_0_reg
				      ,input [31:0] rd_req_desc_e_axuser_1_reg
				      ,input [31:0] rd_req_desc_e_axuser_2_reg
				      ,input [31:0] rd_req_desc_e_axuser_3_reg
				      ,input [31:0] rd_req_desc_e_axuser_4_reg
				      ,input [31:0] rd_req_desc_e_axuser_5_reg
				      ,input [31:0] rd_req_desc_e_axuser_6_reg
				      ,input [31:0] rd_req_desc_e_axuser_7_reg
				      ,input [31:0] rd_req_desc_e_axuser_8_reg
				      ,input [31:0] rd_req_desc_e_axuser_9_reg
				      ,input [31:0] rd_req_desc_e_axuser_10_reg
				      ,input [31:0] rd_req_desc_e_axuser_11_reg
				      ,input [31:0] rd_req_desc_e_axuser_12_reg
				      ,input [31:0] rd_req_desc_e_axuser_13_reg
				      ,input [31:0] rd_req_desc_e_axuser_14_reg
				      ,input [31:0] rd_req_desc_e_axuser_15_reg
				      ,input [31:0] rd_resp_desc_e_data_offset_reg
				      ,input [31:0] rd_resp_desc_e_data_size_reg
				      ,input [31:0] rd_resp_desc_e_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_e_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_e_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_e_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_e_resp_reg
				      ,input [31:0] rd_resp_desc_e_xid_0_reg
				      ,input [31:0] rd_resp_desc_e_xid_1_reg
				      ,input [31:0] rd_resp_desc_e_xid_2_reg
				      ,input [31:0] rd_resp_desc_e_xid_3_reg
				      ,input [31:0] rd_resp_desc_e_xuser_0_reg
				      ,input [31:0] rd_resp_desc_e_xuser_1_reg
				      ,input [31:0] rd_resp_desc_e_xuser_2_reg
				      ,input [31:0] rd_resp_desc_e_xuser_3_reg
				      ,input [31:0] rd_resp_desc_e_xuser_4_reg
				      ,input [31:0] rd_resp_desc_e_xuser_5_reg
				      ,input [31:0] rd_resp_desc_e_xuser_6_reg
				      ,input [31:0] rd_resp_desc_e_xuser_7_reg
				      ,input [31:0] rd_resp_desc_e_xuser_8_reg
				      ,input [31:0] rd_resp_desc_e_xuser_9_reg
				      ,input [31:0] rd_resp_desc_e_xuser_10_reg
				      ,input [31:0] rd_resp_desc_e_xuser_11_reg
				      ,input [31:0] rd_resp_desc_e_xuser_12_reg
				      ,input [31:0] rd_resp_desc_e_xuser_13_reg
				      ,input [31:0] rd_resp_desc_e_xuser_14_reg
				      ,input [31:0] rd_resp_desc_e_xuser_15_reg
				      ,input [31:0] wr_req_desc_e_txn_type_reg
				      ,input [31:0] wr_req_desc_e_size_reg
				      ,input [31:0] wr_req_desc_e_data_offset_reg
				      ,input [31:0] wr_req_desc_e_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_e_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_e_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_e_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_e_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_e_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_e_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_e_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_e_axsize_reg
				      ,input [31:0] wr_req_desc_e_attr_reg
				      ,input [31:0] wr_req_desc_e_axaddr_0_reg
				      ,input [31:0] wr_req_desc_e_axaddr_1_reg
				      ,input [31:0] wr_req_desc_e_axaddr_2_reg
				      ,input [31:0] wr_req_desc_e_axaddr_3_reg
				      ,input [31:0] wr_req_desc_e_axid_0_reg
				      ,input [31:0] wr_req_desc_e_axid_1_reg
				      ,input [31:0] wr_req_desc_e_axid_2_reg
				      ,input [31:0] wr_req_desc_e_axid_3_reg
				      ,input [31:0] wr_req_desc_e_axuser_0_reg
				      ,input [31:0] wr_req_desc_e_axuser_1_reg
				      ,input [31:0] wr_req_desc_e_axuser_2_reg
				      ,input [31:0] wr_req_desc_e_axuser_3_reg
				      ,input [31:0] wr_req_desc_e_axuser_4_reg
				      ,input [31:0] wr_req_desc_e_axuser_5_reg
				      ,input [31:0] wr_req_desc_e_axuser_6_reg
				      ,input [31:0] wr_req_desc_e_axuser_7_reg
				      ,input [31:0] wr_req_desc_e_axuser_8_reg
				      ,input [31:0] wr_req_desc_e_axuser_9_reg
				      ,input [31:0] wr_req_desc_e_axuser_10_reg
				      ,input [31:0] wr_req_desc_e_axuser_11_reg
				      ,input [31:0] wr_req_desc_e_axuser_12_reg
				      ,input [31:0] wr_req_desc_e_axuser_13_reg
				      ,input [31:0] wr_req_desc_e_axuser_14_reg
				      ,input [31:0] wr_req_desc_e_axuser_15_reg
				      ,input [31:0] wr_req_desc_e_wuser_0_reg
				      ,input [31:0] wr_req_desc_e_wuser_1_reg
				      ,input [31:0] wr_req_desc_e_wuser_2_reg
				      ,input [31:0] wr_req_desc_e_wuser_3_reg
				      ,input [31:0] wr_req_desc_e_wuser_4_reg
				      ,input [31:0] wr_req_desc_e_wuser_5_reg
				      ,input [31:0] wr_req_desc_e_wuser_6_reg
				      ,input [31:0] wr_req_desc_e_wuser_7_reg
				      ,input [31:0] wr_req_desc_e_wuser_8_reg
				      ,input [31:0] wr_req_desc_e_wuser_9_reg
				      ,input [31:0] wr_req_desc_e_wuser_10_reg
				      ,input [31:0] wr_req_desc_e_wuser_11_reg
				      ,input [31:0] wr_req_desc_e_wuser_12_reg
				      ,input [31:0] wr_req_desc_e_wuser_13_reg
				      ,input [31:0] wr_req_desc_e_wuser_14_reg
				      ,input [31:0] wr_req_desc_e_wuser_15_reg
				      ,input [31:0] wr_resp_desc_e_resp_reg
				      ,input [31:0] wr_resp_desc_e_xid_0_reg
				      ,input [31:0] wr_resp_desc_e_xid_1_reg
				      ,input [31:0] wr_resp_desc_e_xid_2_reg
				      ,input [31:0] wr_resp_desc_e_xid_3_reg
				      ,input [31:0] wr_resp_desc_e_xuser_0_reg
				      ,input [31:0] wr_resp_desc_e_xuser_1_reg
				      ,input [31:0] wr_resp_desc_e_xuser_2_reg
				      ,input [31:0] wr_resp_desc_e_xuser_3_reg
				      ,input [31:0] wr_resp_desc_e_xuser_4_reg
				      ,input [31:0] wr_resp_desc_e_xuser_5_reg
				      ,input [31:0] wr_resp_desc_e_xuser_6_reg
				      ,input [31:0] wr_resp_desc_e_xuser_7_reg
				      ,input [31:0] wr_resp_desc_e_xuser_8_reg
				      ,input [31:0] wr_resp_desc_e_xuser_9_reg
				      ,input [31:0] wr_resp_desc_e_xuser_10_reg
				      ,input [31:0] wr_resp_desc_e_xuser_11_reg
				      ,input [31:0] wr_resp_desc_e_xuser_12_reg
				      ,input [31:0] wr_resp_desc_e_xuser_13_reg
				      ,input [31:0] wr_resp_desc_e_xuser_14_reg
				      ,input [31:0] wr_resp_desc_e_xuser_15_reg
				      ,input [31:0] sn_req_desc_e_attr_reg
				      ,input [31:0] sn_req_desc_e_acaddr_0_reg
				      ,input [31:0] sn_req_desc_e_acaddr_1_reg
				      ,input [31:0] sn_req_desc_e_acaddr_2_reg
				      ,input [31:0] sn_req_desc_e_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_e_resp_reg
				      ,input [31:0] rd_req_desc_f_txn_type_reg
				      ,input [31:0] rd_req_desc_f_size_reg
				      ,input [31:0] rd_req_desc_f_axsize_reg
				      ,input [31:0] rd_req_desc_f_attr_reg
				      ,input [31:0] rd_req_desc_f_axaddr_0_reg
				      ,input [31:0] rd_req_desc_f_axaddr_1_reg
				      ,input [31:0] rd_req_desc_f_axaddr_2_reg
				      ,input [31:0] rd_req_desc_f_axaddr_3_reg
				      ,input [31:0] rd_req_desc_f_axid_0_reg
				      ,input [31:0] rd_req_desc_f_axid_1_reg
				      ,input [31:0] rd_req_desc_f_axid_2_reg
				      ,input [31:0] rd_req_desc_f_axid_3_reg
				      ,input [31:0] rd_req_desc_f_axuser_0_reg
				      ,input [31:0] rd_req_desc_f_axuser_1_reg
				      ,input [31:0] rd_req_desc_f_axuser_2_reg
				      ,input [31:0] rd_req_desc_f_axuser_3_reg
				      ,input [31:0] rd_req_desc_f_axuser_4_reg
				      ,input [31:0] rd_req_desc_f_axuser_5_reg
				      ,input [31:0] rd_req_desc_f_axuser_6_reg
				      ,input [31:0] rd_req_desc_f_axuser_7_reg
				      ,input [31:0] rd_req_desc_f_axuser_8_reg
				      ,input [31:0] rd_req_desc_f_axuser_9_reg
				      ,input [31:0] rd_req_desc_f_axuser_10_reg
				      ,input [31:0] rd_req_desc_f_axuser_11_reg
				      ,input [31:0] rd_req_desc_f_axuser_12_reg
				      ,input [31:0] rd_req_desc_f_axuser_13_reg
				      ,input [31:0] rd_req_desc_f_axuser_14_reg
				      ,input [31:0] rd_req_desc_f_axuser_15_reg
				      ,input [31:0] rd_resp_desc_f_data_offset_reg
				      ,input [31:0] rd_resp_desc_f_data_size_reg
				      ,input [31:0] rd_resp_desc_f_data_host_addr_0_reg
				      ,input [31:0] rd_resp_desc_f_data_host_addr_1_reg
				      ,input [31:0] rd_resp_desc_f_data_host_addr_2_reg
				      ,input [31:0] rd_resp_desc_f_data_host_addr_3_reg
				      ,input [31:0] rd_resp_desc_f_resp_reg
				      ,input [31:0] rd_resp_desc_f_xid_0_reg
				      ,input [31:0] rd_resp_desc_f_xid_1_reg
				      ,input [31:0] rd_resp_desc_f_xid_2_reg
				      ,input [31:0] rd_resp_desc_f_xid_3_reg
				      ,input [31:0] rd_resp_desc_f_xuser_0_reg
				      ,input [31:0] rd_resp_desc_f_xuser_1_reg
				      ,input [31:0] rd_resp_desc_f_xuser_2_reg
				      ,input [31:0] rd_resp_desc_f_xuser_3_reg
				      ,input [31:0] rd_resp_desc_f_xuser_4_reg
				      ,input [31:0] rd_resp_desc_f_xuser_5_reg
				      ,input [31:0] rd_resp_desc_f_xuser_6_reg
				      ,input [31:0] rd_resp_desc_f_xuser_7_reg
				      ,input [31:0] rd_resp_desc_f_xuser_8_reg
				      ,input [31:0] rd_resp_desc_f_xuser_9_reg
				      ,input [31:0] rd_resp_desc_f_xuser_10_reg
				      ,input [31:0] rd_resp_desc_f_xuser_11_reg
				      ,input [31:0] rd_resp_desc_f_xuser_12_reg
				      ,input [31:0] rd_resp_desc_f_xuser_13_reg
				      ,input [31:0] rd_resp_desc_f_xuser_14_reg
				      ,input [31:0] rd_resp_desc_f_xuser_15_reg
				      ,input [31:0] wr_req_desc_f_txn_type_reg
				      ,input [31:0] wr_req_desc_f_size_reg
				      ,input [31:0] wr_req_desc_f_data_offset_reg
				      ,input [31:0] wr_req_desc_f_data_host_addr_0_reg
				      ,input [31:0] wr_req_desc_f_data_host_addr_1_reg
				      ,input [31:0] wr_req_desc_f_data_host_addr_2_reg
				      ,input [31:0] wr_req_desc_f_data_host_addr_3_reg
				      ,input [31:0] wr_req_desc_f_wstrb_host_addr_0_reg
				      ,input [31:0] wr_req_desc_f_wstrb_host_addr_1_reg
				      ,input [31:0] wr_req_desc_f_wstrb_host_addr_2_reg
				      ,input [31:0] wr_req_desc_f_wstrb_host_addr_3_reg
				      ,input [31:0] wr_req_desc_f_axsize_reg
				      ,input [31:0] wr_req_desc_f_attr_reg
				      ,input [31:0] wr_req_desc_f_axaddr_0_reg
				      ,input [31:0] wr_req_desc_f_axaddr_1_reg
				      ,input [31:0] wr_req_desc_f_axaddr_2_reg
				      ,input [31:0] wr_req_desc_f_axaddr_3_reg
				      ,input [31:0] wr_req_desc_f_axid_0_reg
				      ,input [31:0] wr_req_desc_f_axid_1_reg
				      ,input [31:0] wr_req_desc_f_axid_2_reg
				      ,input [31:0] wr_req_desc_f_axid_3_reg
				      ,input [31:0] wr_req_desc_f_axuser_0_reg
				      ,input [31:0] wr_req_desc_f_axuser_1_reg
				      ,input [31:0] wr_req_desc_f_axuser_2_reg
				      ,input [31:0] wr_req_desc_f_axuser_3_reg
				      ,input [31:0] wr_req_desc_f_axuser_4_reg
				      ,input [31:0] wr_req_desc_f_axuser_5_reg
				      ,input [31:0] wr_req_desc_f_axuser_6_reg
				      ,input [31:0] wr_req_desc_f_axuser_7_reg
				      ,input [31:0] wr_req_desc_f_axuser_8_reg
				      ,input [31:0] wr_req_desc_f_axuser_9_reg
				      ,input [31:0] wr_req_desc_f_axuser_10_reg
				      ,input [31:0] wr_req_desc_f_axuser_11_reg
				      ,input [31:0] wr_req_desc_f_axuser_12_reg
				      ,input [31:0] wr_req_desc_f_axuser_13_reg
				      ,input [31:0] wr_req_desc_f_axuser_14_reg
				      ,input [31:0] wr_req_desc_f_axuser_15_reg
				      ,input [31:0] wr_req_desc_f_wuser_0_reg
				      ,input [31:0] wr_req_desc_f_wuser_1_reg
				      ,input [31:0] wr_req_desc_f_wuser_2_reg
				      ,input [31:0] wr_req_desc_f_wuser_3_reg
				      ,input [31:0] wr_req_desc_f_wuser_4_reg
				      ,input [31:0] wr_req_desc_f_wuser_5_reg
				      ,input [31:0] wr_req_desc_f_wuser_6_reg
				      ,input [31:0] wr_req_desc_f_wuser_7_reg
				      ,input [31:0] wr_req_desc_f_wuser_8_reg
				      ,input [31:0] wr_req_desc_f_wuser_9_reg
				      ,input [31:0] wr_req_desc_f_wuser_10_reg
				      ,input [31:0] wr_req_desc_f_wuser_11_reg
				      ,input [31:0] wr_req_desc_f_wuser_12_reg
				      ,input [31:0] wr_req_desc_f_wuser_13_reg
				      ,input [31:0] wr_req_desc_f_wuser_14_reg
				      ,input [31:0] wr_req_desc_f_wuser_15_reg
				      ,input [31:0] wr_resp_desc_f_resp_reg
				      ,input [31:0] wr_resp_desc_f_xid_0_reg
				      ,input [31:0] wr_resp_desc_f_xid_1_reg
				      ,input [31:0] wr_resp_desc_f_xid_2_reg
				      ,input [31:0] wr_resp_desc_f_xid_3_reg
				      ,input [31:0] wr_resp_desc_f_xuser_0_reg
				      ,input [31:0] wr_resp_desc_f_xuser_1_reg
				      ,input [31:0] wr_resp_desc_f_xuser_2_reg
				      ,input [31:0] wr_resp_desc_f_xuser_3_reg
				      ,input [31:0] wr_resp_desc_f_xuser_4_reg
				      ,input [31:0] wr_resp_desc_f_xuser_5_reg
				      ,input [31:0] wr_resp_desc_f_xuser_6_reg
				      ,input [31:0] wr_resp_desc_f_xuser_7_reg
				      ,input [31:0] wr_resp_desc_f_xuser_8_reg
				      ,input [31:0] wr_resp_desc_f_xuser_9_reg
				      ,input [31:0] wr_resp_desc_f_xuser_10_reg
				      ,input [31:0] wr_resp_desc_f_xuser_11_reg
				      ,input [31:0] wr_resp_desc_f_xuser_12_reg
				      ,input [31:0] wr_resp_desc_f_xuser_13_reg
				      ,input [31:0] wr_resp_desc_f_xuser_14_reg
				      ,input [31:0] wr_resp_desc_f_xuser_15_reg
				      ,input [31:0] sn_req_desc_f_attr_reg
				      ,input [31:0] sn_req_desc_f_acaddr_0_reg
				      ,input [31:0] sn_req_desc_f_acaddr_1_reg
				      ,input [31:0] sn_req_desc_f_acaddr_2_reg
				      ,input [31:0] sn_req_desc_f_acaddr_3_reg
				      ,input [31:0] sn_resp_desc_f_resp_reg
   
   
				      ,output [31:0] uc2rb_intr_error_status_reg
				      ,output [31:0] uc2rb_rd_req_fifo_pop_desc_reg
				      ,output [31:0] uc2rb_rd_req_fifo_fill_level_reg
				      ,output [31:0] uc2rb_rd_resp_fifo_free_level_reg
				      ,output [31:0] uc2rb_rd_resp_intr_comp_status_reg
				      ,output [31:0] uc2rb_wr_req_fifo_pop_desc_reg
				      ,output [31:0] uc2rb_wr_req_fifo_fill_level_reg
				      ,output [31:0] uc2rb_wr_resp_fifo_free_level_reg
				      ,output [31:0] uc2rb_wr_resp_intr_comp_status_reg
				      ,output [31:0] uc2rb_sn_req_fifo_free_level_reg
				      ,output [31:0] uc2rb_sn_req_intr_comp_status_reg
				      ,output [31:0] uc2rb_sn_resp_fifo_pop_desc_reg
				      ,output [31:0] uc2rb_sn_resp_fifo_fill_level_reg
				      ,output [31:0] uc2rb_sn_data_fifo_pop_desc_reg
				      ,output [31:0] uc2rb_sn_data_fifo_fill_level_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_0_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_1_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_2_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_3_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_4_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_5_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_6_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_7_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_8_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_9_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_a_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_b_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_c_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_d_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_e_resp_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_txn_type_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_size_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axsize_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_attr_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_0_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_1_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_2_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_3_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_4_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_5_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_6_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_7_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_8_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_9_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_10_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_11_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_12_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_13_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_14_reg
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_txn_type_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_size_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_data_offset_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axsize_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_attr_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_15_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_0_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_1_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_2_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_3_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_4_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_5_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_6_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_7_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_8_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_9_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_10_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_11_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_12_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_13_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_14_reg
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_15_reg
				      ,output [31:0] uc2rb_sn_resp_desc_f_resp_reg
   
   
				      ,output [31:0] uc2rb_intr_error_status_reg_we
				      ,output [31:0] uc2rb_rd_req_fifo_pop_desc_reg_we
				      ,output [31:0] uc2rb_rd_req_fifo_fill_level_reg_we
				      ,output [31:0] uc2rb_rd_resp_fifo_free_level_reg_we
				      ,output [31:0] uc2rb_rd_resp_intr_comp_status_reg_we
				      ,output [31:0] uc2rb_wr_req_fifo_pop_desc_reg_we
				      ,output [31:0] uc2rb_wr_req_fifo_fill_level_reg_we
				      ,output [31:0] uc2rb_wr_resp_fifo_free_level_reg_we
				      ,output [31:0] uc2rb_wr_resp_intr_comp_status_reg_we
				      ,output [31:0] uc2rb_sn_req_fifo_free_level_reg_we
				      ,output [31:0] uc2rb_sn_req_intr_comp_status_reg_we
				      ,output [31:0] uc2rb_sn_resp_fifo_pop_desc_reg_we
				      ,output [31:0] uc2rb_sn_resp_fifo_fill_level_reg_we
				      ,output [31:0] uc2rb_sn_data_fifo_pop_desc_reg_we
				      ,output [31:0] uc2rb_sn_data_fifo_fill_level_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_0_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_0_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_0_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_1_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_1_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_1_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_2_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_2_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_2_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_3_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_3_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_3_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_4_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_4_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_4_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_5_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_5_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_5_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_6_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_6_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_6_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_7_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_7_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_7_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_8_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_8_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_8_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_9_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_9_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_9_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_a_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_a_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_a_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_b_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_b_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_b_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_c_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_c_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_c_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_d_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_d_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_d_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_e_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_e_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_e_resp_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_txn_type_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_size_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axsize_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_attr_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axaddr_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axid_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_0_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_1_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_2_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_3_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_4_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_5_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_6_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_7_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_8_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_9_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_10_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_11_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_12_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_13_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_14_reg_we
				      ,output [31:0] uc2rb_rd_req_desc_f_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_txn_type_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_size_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_data_offset_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axsize_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_attr_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axaddr_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axid_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_axuser_15_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_0_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_1_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_2_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_3_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_4_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_5_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_6_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_7_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_8_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_9_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_10_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_11_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_12_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_13_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_14_reg_we
				      ,output [31:0] uc2rb_wr_req_desc_f_wuser_15_reg_we
				      ,output [31:0] uc2rb_sn_resp_desc_f_resp_reg_we
   
   
				      //RAM commands  
				      //RDATA_RAM
				      ,output [(`CLOG2((XX_RAM_SIZE*8)/XX_DATA_WIDTH))-1:0] uc2rb_rd_addr 
				      ,input [XX_DATA_WIDTH-1:0] rb2uc_rd_data 
   
				      //WDATA_RAM and WSTRB_RAM                               
				      ,output uc2rb_wr_we 
				      ,output [(XX_DATA_WIDTH/8)-1:0] uc2rb_wr_bwe //Generate all 1s always.     
				      ,output [(`CLOG2((XX_RAM_SIZE*8)/XX_DATA_WIDTH))-1:0] uc2rb_wr_addr 
				      ,output [XX_DATA_WIDTH-1:0] uc2rb_wr_data 
				      ,output [(XX_DATA_WIDTH/8)-1:0] uc2rb_wr_wstrb 
   
				      //CDDATA_RAM                               
				      ,output uc2rb_sn_we 
				      ,output [(SN_DATA_WIDTH/8)-1:0] uc2rb_sn_bwe //Generate all 1s always.     
				      ,output [(`CLOG2((SN_RAM_SIZE*8)/SN_DATA_WIDTH))-1:0] uc2rb_sn_addr 
				      ,output [SN_DATA_WIDTH-1:0] uc2rb_sn_data 
   
				      ,output [XX_MAX_DESC-1:0] rd_uc2hm_trig 
				      ,input [XX_MAX_DESC-1:0] rd_hm2uc_done
				      ,output [XX_MAX_DESC-1:0] wr_uc2hm_trig 
				      ,input [XX_MAX_DESC-1:0] wr_hm2uc_done
   
				      //pop request to FIFO
				      ,input rd_req_fifo_pop_desc_conn 
				      ,input wr_req_fifo_pop_desc_conn 
				      ,input sn_resp_fifo_pop_desc_conn
				      ,input sn_data_fifo_pop_desc_conn
   
				      //output from FIFO
				      ,output [(`CLOG2(XX_MAX_DESC))-1:0] rd_req_fifo_out
				      ,output rd_req_fifo_out_valid //it is one clock cycle pulse
				      ,output [(`CLOG2(XX_MAX_DESC))-1:0] wr_req_fifo_out
				      ,output wr_req_fifo_out_valid //it is one clock cycle pulse
				      ,output [(`CLOG2(SN_MAX_DESC))-1:0] sn_resp_fifo_out
				      ,output sn_resp_fifo_out_valid //it is one clock cycle pulse
				      ,output [(`CLOG2(SN_MAX_DESC))-1:0] sn_data_fifo_out
				      ,output sn_data_fifo_out_valid  //it is one clock cycle pulse


				      );
   
   localparam XX_DESC_IDX_WIDTH                                            = `CLOG2(XX_MAX_DESC);
   localparam XX_RAM_OFFSET_WIDTH                                          = `CLOG2((XX_RAM_SIZE*8)/XX_DATA_WIDTH);

   //Declare all fields ( <reg>_<field>_f )

   wire [0:0] 				    bridge_identification_last_bridge_f;
   wire [7:0] 				    version_major_ver_f;
   wire [7:0] 				    version_minor_ver_f;
   wire [7:0] 				    bridge_type_type_f;
   wire [0:0] 				    bridge_config_extend_wstrb_f;
   wire [7:0] 				    bridge_config_id_width_f;
   wire [2:0] 				    bridge_config_data_width_f;
   wire [9:0] 				    bridge_rd_user_config_ruser_width_f;
   wire [9:0] 				    bridge_rd_user_config_aruser_width_f;
   wire [9:0] 				    bridge_wr_user_config_buser_width_f;
   wire [9:0] 				    bridge_wr_user_config_wuser_width_f;
   wire [9:0] 				    bridge_wr_user_config_awuser_width_f;
   wire [7:0] 				    rd_max_desc_resp_max_desc_f;
   wire [7:0] 				    rd_max_desc_req_max_desc_f;
   wire [7:0] 				    wr_max_desc_resp_max_desc_f;
   wire [7:0] 				    wr_max_desc_req_max_desc_f;
   wire [7:0] 				    sn_max_desc_data_max_desc_f;
   wire [7:0] 				    sn_max_desc_resp_max_desc_f;
   wire [7:0] 				    sn_max_desc_req_max_desc_f;
   wire [0:0] 				    reset_dut_srst_3_f;
   wire [0:0] 				    reset_dut_srst_2_f;
   wire [0:0] 				    reset_dut_srst_1_f;
   wire [0:0] 				    reset_dut_srst_0_f;
   wire [0:0] 				    reset_srst_f;
   wire [0:0] 				    mode_select_mode_0_1_f;
   wire [0:0] 				    intr_status_sn_data_fifo_nonempty_f;
   wire [0:0] 				    intr_status_sn_resp_fifo_nonempty_f;
   wire [0:0] 				    intr_status_sn_req_comp_f;
   wire [0:0] 				    intr_status_wr_resp_comp_f;
   wire [0:0] 				    intr_status_wr_req_fifo_nonempty_f;
   wire [0:0] 				    intr_status_rd_resp_comp_f;
   wire [0:0] 				    intr_status_rd_req_fifo_nonempty_f;
   wire [0:0] 				    intr_status_c2h_f;
   wire [0:0] 				    intr_status_error_f;
   wire [0:0] 				    intr_error_status_err_1_f;
   wire [0:0] 				    intr_error_status_err_0_f;
   wire [0:0] 				    intr_error_clear_clr_err_2_f;
   wire [0:0] 				    intr_error_clear_clr_err_1_f;
   wire [0:0] 				    intr_error_clear_clr_err_0_f;
   wire [0:0] 				    intr_error_enable_en_err_2_f;
   wire [0:0] 				    intr_error_enable_en_err_1_f;
   wire [0:0] 				    intr_error_enable_en_err_0_f;
   wire [15:0] 				    rd_req_free_desc_desc_f;
   wire [0:0] 				    rd_req_fifo_pop_desc_valid_f;
   wire [3:0] 				    rd_req_fifo_pop_desc_desc_index_f;
   wire [4:0] 				    rd_req_fifo_fill_level_fill_f;
   wire [0:0] 				    rd_resp_fifo_push_desc_valid_f;
   wire [3:0] 				    rd_resp_fifo_push_desc_desc_index_f;
   wire [4:0] 				    rd_resp_fifo_free_level_free_f;
   wire [15:0] 				    rd_resp_intr_comp_status_comp_f;
   wire [15:0] 				    rd_resp_intr_comp_clear_clr_comp_f;
   wire [15:0] 				    rd_resp_intr_comp_enable_en_comp_f;
   wire [15:0] 				    wr_req_free_desc_desc_f;
   wire [0:0] 				    wr_req_fifo_pop_desc_valid_f;
   wire [3:0] 				    wr_req_fifo_pop_desc_desc_index_f;
   wire [4:0] 				    wr_req_fifo_fill_level_fill_f;
   wire [0:0] 				    wr_resp_fifo_push_desc_valid_f;
   wire [3:0] 				    wr_resp_fifo_push_desc_desc_index_f;
   wire [4:0] 				    wr_resp_fifo_free_level_free_f;
   wire [15:0] 				    wr_resp_intr_comp_status_comp_f;
   wire [15:0] 				    wr_resp_intr_comp_clear_clr_comp_f;
   wire [15:0] 				    wr_resp_intr_comp_enable_en_comp_f;
   wire [0:0] 				    sn_req_fifo_push_desc_valid_f;
   wire [3:0] 				    sn_req_fifo_push_desc_desc_index_f;
   wire [4:0] 				    sn_req_fifo_free_level_free_f;
   wire [15:0] 				    sn_req_intr_comp_status_comp_f;
   wire [15:0] 				    sn_req_intr_comp_clear_clr_comp_f;
   wire [15:0] 				    sn_req_intr_comp_enable_en_comp_f;
   wire [15:0] 				    sn_resp_free_desc_desc_f;
   wire [0:0] 				    sn_resp_fifo_pop_desc_valid_f;
   wire [3:0] 				    sn_resp_fifo_pop_desc_desc_index_f;
   wire [4:0] 				    sn_resp_fifo_fill_level_fill_f;
   wire [15:0] 				    sn_data_free_desc_desc_f;
   wire [0:0] 				    sn_data_fifo_pop_desc_valid_f;
   wire [3:0] 				    sn_data_fifo_pop_desc_desc_index_f;
   wire [4:0] 				    sn_data_fifo_fill_level_fill_f;
   wire [0:0] 				    intr_fifo_enable_en_sn_data_fifo_nonempty_f;
   wire [0:0] 				    intr_fifo_enable_en_sn_resp_fifo_nonempty_f;
   wire [0:0] 				    intr_fifo_enable_en_wr_req_fifo_nonempty_f;
   wire [0:0] 				    intr_fifo_enable_en_rd_req_fifo_nonempty_f;
   wire [0:0] 				    h2c_intr_0_h2c_31_f;
   wire [0:0] 				    h2c_intr_0_h2c_30_f;
   wire [0:0] 				    h2c_intr_0_h2c_29_f;
   wire [0:0] 				    h2c_intr_0_h2c_28_f;
   wire [0:0] 				    h2c_intr_0_h2c_27_f;
   wire [0:0] 				    h2c_intr_0_h2c_26_f;
   wire [0:0] 				    h2c_intr_0_h2c_25_f;
   wire [0:0] 				    h2c_intr_0_h2c_24_f;
   wire [0:0] 				    h2c_intr_0_h2c_23_f;
   wire [0:0] 				    h2c_intr_0_h2c_22_f;
   wire [0:0] 				    h2c_intr_0_h2c_21_f;
   wire [0:0] 				    h2c_intr_0_h2c_20_f;
   wire [0:0] 				    h2c_intr_0_h2c_19_f;
   wire [0:0] 				    h2c_intr_0_h2c_18_f;
   wire [0:0] 				    h2c_intr_0_h2c_17_f;
   wire [0:0] 				    h2c_intr_0_h2c_16_f;
   wire [0:0] 				    h2c_intr_0_h2c_15_f;
   wire [0:0] 				    h2c_intr_0_h2c_14_f;
   wire [0:0] 				    h2c_intr_0_h2c_13_f;
   wire [0:0] 				    h2c_intr_0_h2c_12_f;
   wire [0:0] 				    h2c_intr_0_h2c_11_f;
   wire [0:0] 				    h2c_intr_0_h2c_10_f;
   wire [0:0] 				    h2c_intr_0_h2c_9_f;
   wire [0:0] 				    h2c_intr_0_h2c_8_f;
   wire [0:0] 				    h2c_intr_0_h2c_7_f;
   wire [0:0] 				    h2c_intr_0_h2c_6_f;
   wire [0:0] 				    h2c_intr_0_h2c_5_f;
   wire [0:0] 				    h2c_intr_0_h2c_4_f;
   wire [0:0] 				    h2c_intr_0_h2c_3_f;
   wire [0:0] 				    h2c_intr_0_h2c_2_f;
   wire [0:0] 				    h2c_intr_0_h2c_1_f;
   wire [0:0] 				    h2c_intr_0_h2c_0_f;
   wire [0:0] 				    h2c_intr_1_h2c_31_f;
   wire [0:0] 				    h2c_intr_1_h2c_30_f;
   wire [0:0] 				    h2c_intr_1_h2c_29_f;
   wire [0:0] 				    h2c_intr_1_h2c_28_f;
   wire [0:0] 				    h2c_intr_1_h2c_27_f;
   wire [0:0] 				    h2c_intr_1_h2c_26_f;
   wire [0:0] 				    h2c_intr_1_h2c_25_f;
   wire [0:0] 				    h2c_intr_1_h2c_24_f;
   wire [0:0] 				    h2c_intr_1_h2c_23_f;
   wire [0:0] 				    h2c_intr_1_h2c_22_f;
   wire [0:0] 				    h2c_intr_1_h2c_21_f;
   wire [0:0] 				    h2c_intr_1_h2c_20_f;
   wire [0:0] 				    h2c_intr_1_h2c_19_f;
   wire [0:0] 				    h2c_intr_1_h2c_18_f;
   wire [0:0] 				    h2c_intr_1_h2c_17_f;
   wire [0:0] 				    h2c_intr_1_h2c_16_f;
   wire [0:0] 				    h2c_intr_1_h2c_15_f;
   wire [0:0] 				    h2c_intr_1_h2c_14_f;
   wire [0:0] 				    h2c_intr_1_h2c_13_f;
   wire [0:0] 				    h2c_intr_1_h2c_12_f;
   wire [0:0] 				    h2c_intr_1_h2c_11_f;
   wire [0:0] 				    h2c_intr_1_h2c_10_f;
   wire [0:0] 				    h2c_intr_1_h2c_9_f;
   wire [0:0] 				    h2c_intr_1_h2c_8_f;
   wire [0:0] 				    h2c_intr_1_h2c_7_f;
   wire [0:0] 				    h2c_intr_1_h2c_6_f;
   wire [0:0] 				    h2c_intr_1_h2c_5_f;
   wire [0:0] 				    h2c_intr_1_h2c_4_f;
   wire [0:0] 				    h2c_intr_1_h2c_3_f;
   wire [0:0] 				    h2c_intr_1_h2c_2_f;
   wire [0:0] 				    h2c_intr_1_h2c_1_f;
   wire [0:0] 				    h2c_intr_1_h2c_0_f;
   wire [0:0] 				    h2c_intr_2_h2c_31_f;
   wire [0:0] 				    h2c_intr_2_h2c_30_f;
   wire [0:0] 				    h2c_intr_2_h2c_29_f;
   wire [0:0] 				    h2c_intr_2_h2c_28_f;
   wire [0:0] 				    h2c_intr_2_h2c_27_f;
   wire [0:0] 				    h2c_intr_2_h2c_26_f;
   wire [0:0] 				    h2c_intr_2_h2c_25_f;
   wire [0:0] 				    h2c_intr_2_h2c_24_f;
   wire [0:0] 				    h2c_intr_2_h2c_23_f;
   wire [0:0] 				    h2c_intr_2_h2c_22_f;
   wire [0:0] 				    h2c_intr_2_h2c_21_f;
   wire [0:0] 				    h2c_intr_2_h2c_20_f;
   wire [0:0] 				    h2c_intr_2_h2c_19_f;
   wire [0:0] 				    h2c_intr_2_h2c_18_f;
   wire [0:0] 				    h2c_intr_2_h2c_17_f;
   wire [0:0] 				    h2c_intr_2_h2c_16_f;
   wire [0:0] 				    h2c_intr_2_h2c_15_f;
   wire [0:0] 				    h2c_intr_2_h2c_14_f;
   wire [0:0] 				    h2c_intr_2_h2c_13_f;
   wire [0:0] 				    h2c_intr_2_h2c_12_f;
   wire [0:0] 				    h2c_intr_2_h2c_11_f;
   wire [0:0] 				    h2c_intr_2_h2c_10_f;
   wire [0:0] 				    h2c_intr_2_h2c_9_f;
   wire [0:0] 				    h2c_intr_2_h2c_8_f;
   wire [0:0] 				    h2c_intr_2_h2c_7_f;
   wire [0:0] 				    h2c_intr_2_h2c_6_f;
   wire [0:0] 				    h2c_intr_2_h2c_5_f;
   wire [0:0] 				    h2c_intr_2_h2c_4_f;
   wire [0:0] 				    h2c_intr_2_h2c_3_f;
   wire [0:0] 				    h2c_intr_2_h2c_2_f;
   wire [0:0] 				    h2c_intr_2_h2c_1_f;
   wire [0:0] 				    h2c_intr_2_h2c_0_f;
   wire [0:0] 				    h2c_intr_3_h2c_31_f;
   wire [0:0] 				    h2c_intr_3_h2c_30_f;
   wire [0:0] 				    h2c_intr_3_h2c_29_f;
   wire [0:0] 				    h2c_intr_3_h2c_28_f;
   wire [0:0] 				    h2c_intr_3_h2c_27_f;
   wire [0:0] 				    h2c_intr_3_h2c_26_f;
   wire [0:0] 				    h2c_intr_3_h2c_25_f;
   wire [0:0] 				    h2c_intr_3_h2c_24_f;
   wire [0:0] 				    h2c_intr_3_h2c_23_f;
   wire [0:0] 				    h2c_intr_3_h2c_22_f;
   wire [0:0] 				    h2c_intr_3_h2c_21_f;
   wire [0:0] 				    h2c_intr_3_h2c_20_f;
   wire [0:0] 				    h2c_intr_3_h2c_19_f;
   wire [0:0] 				    h2c_intr_3_h2c_18_f;
   wire [0:0] 				    h2c_intr_3_h2c_17_f;
   wire [0:0] 				    h2c_intr_3_h2c_16_f;
   wire [0:0] 				    h2c_intr_3_h2c_15_f;
   wire [0:0] 				    h2c_intr_3_h2c_14_f;
   wire [0:0] 				    h2c_intr_3_h2c_13_f;
   wire [0:0] 				    h2c_intr_3_h2c_12_f;
   wire [0:0] 				    h2c_intr_3_h2c_11_f;
   wire [0:0] 				    h2c_intr_3_h2c_10_f;
   wire [0:0] 				    h2c_intr_3_h2c_9_f;
   wire [0:0] 				    h2c_intr_3_h2c_8_f;
   wire [0:0] 				    h2c_intr_3_h2c_7_f;
   wire [0:0] 				    h2c_intr_3_h2c_6_f;
   wire [0:0] 				    h2c_intr_3_h2c_5_f;
   wire [0:0] 				    h2c_intr_3_h2c_4_f;
   wire [0:0] 				    h2c_intr_3_h2c_3_f;
   wire [0:0] 				    h2c_intr_3_h2c_2_f;
   wire [0:0] 				    h2c_intr_3_h2c_1_f;
   wire [0:0] 				    h2c_intr_3_h2c_0_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_31_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_30_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_29_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_28_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_27_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_26_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_25_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_24_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_23_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_22_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_21_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_20_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_19_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_18_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_17_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_16_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_15_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_14_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_13_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_12_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_11_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_10_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_9_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_8_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_7_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_6_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_5_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_4_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_3_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_2_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_1_f;
   wire [0:0] 				    c2h_intr_status_0_c2h_0_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_31_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_30_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_29_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_28_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_27_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_26_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_25_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_24_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_23_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_22_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_21_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_20_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_19_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_18_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_17_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_16_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_15_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_14_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_13_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_12_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_11_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_10_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_9_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_8_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_7_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_6_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_5_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_4_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_3_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_2_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_1_f;
   wire [0:0] 				    intr_c2h_toggle_status_0_t_c2h_0_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_31_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_30_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_29_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_28_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_27_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_26_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_25_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_24_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_23_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_22_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_21_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_20_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_19_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_18_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_17_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_16_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_15_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_14_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_13_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_12_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_11_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_10_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_9_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_8_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_7_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_6_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_5_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_4_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_3_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_2_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_1_f;
   wire [0:0] 				    intr_c2h_toggle_clear_0_clr_t_c2h_0_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_31_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_30_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_29_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_28_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_27_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_26_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_25_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_24_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_23_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_22_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_21_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_20_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_19_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_18_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_17_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_16_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_15_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_14_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_13_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_12_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_11_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_10_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_9_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_8_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_7_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_6_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_5_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_4_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_3_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_2_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_1_f;
   wire [0:0] 				    intr_c2h_toggle_enable_0_en_t_c2h_0_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_31_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_30_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_29_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_28_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_27_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_26_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_25_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_24_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_23_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_22_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_21_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_20_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_19_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_18_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_17_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_16_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_15_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_14_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_13_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_12_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_11_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_10_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_9_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_8_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_7_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_6_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_5_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_4_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_3_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_2_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_1_f;
   wire [0:0] 				    c2h_intr_status_1_c2h_0_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_31_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_30_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_29_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_28_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_27_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_26_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_25_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_24_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_23_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_22_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_21_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_20_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_19_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_18_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_17_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_16_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_15_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_14_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_13_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_12_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_11_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_10_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_9_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_8_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_7_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_6_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_5_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_4_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_3_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_2_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_1_f;
   wire [0:0] 				    intr_c2h_toggle_status_1_t_c2h_0_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_31_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_30_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_29_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_28_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_27_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_26_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_25_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_24_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_23_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_22_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_21_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_20_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_19_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_18_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_17_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_16_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_15_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_14_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_13_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_12_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_11_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_10_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_9_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_8_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_7_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_6_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_5_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_4_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_3_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_2_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_1_f;
   wire [0:0] 				    intr_c2h_toggle_clear_1_clr_t_c2h_0_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_31_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_30_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_29_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_28_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_27_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_26_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_25_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_24_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_23_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_22_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_21_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_20_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_19_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_18_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_17_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_16_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_15_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_14_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_13_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_12_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_11_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_10_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_9_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_8_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_7_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_6_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_5_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_4_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_3_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_2_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_1_f;
   wire [0:0] 				    intr_c2h_toggle_enable_1_en_t_c2h_0_f;
   wire [0:0] 				    c2h_gpio_0_gpio_31_f;
   wire [0:0] 				    c2h_gpio_0_gpio_30_f;
   wire [0:0] 				    c2h_gpio_0_gpio_29_f;
   wire [0:0] 				    c2h_gpio_0_gpio_28_f;
   wire [0:0] 				    c2h_gpio_0_gpio_27_f;
   wire [0:0] 				    c2h_gpio_0_gpio_26_f;
   wire [0:0] 				    c2h_gpio_0_gpio_25_f;
   wire [0:0] 				    c2h_gpio_0_gpio_24_f;
   wire [0:0] 				    c2h_gpio_0_gpio_23_f;
   wire [0:0] 				    c2h_gpio_0_gpio_22_f;
   wire [0:0] 				    c2h_gpio_0_gpio_21_f;
   wire [0:0] 				    c2h_gpio_0_gpio_20_f;
   wire [0:0] 				    c2h_gpio_0_gpio_19_f;
   wire [0:0] 				    c2h_gpio_0_gpio_18_f;
   wire [0:0] 				    c2h_gpio_0_gpio_17_f;
   wire [0:0] 				    c2h_gpio_0_gpio_16_f;
   wire [0:0] 				    c2h_gpio_0_gpio_15_f;
   wire [0:0] 				    c2h_gpio_0_gpio_14_f;
   wire [0:0] 				    c2h_gpio_0_gpio_13_f;
   wire [0:0] 				    c2h_gpio_0_gpio_12_f;
   wire [0:0] 				    c2h_gpio_0_gpio_11_f;
   wire [0:0] 				    c2h_gpio_0_gpio_10_f;
   wire [0:0] 				    c2h_gpio_0_gpio_9_f;
   wire [0:0] 				    c2h_gpio_0_gpio_8_f;
   wire [0:0] 				    c2h_gpio_0_gpio_7_f;
   wire [0:0] 				    c2h_gpio_0_gpio_6_f;
   wire [0:0] 				    c2h_gpio_0_gpio_5_f;
   wire [0:0] 				    c2h_gpio_0_gpio_4_f;
   wire [0:0] 				    c2h_gpio_0_gpio_3_f;
   wire [0:0] 				    c2h_gpio_0_gpio_2_f;
   wire [0:0] 				    c2h_gpio_0_gpio_1_f;
   wire [0:0] 				    c2h_gpio_0_gpio_0_f;
   wire [0:0] 				    c2h_gpio_1_gpio_31_f;
   wire [0:0] 				    c2h_gpio_1_gpio_30_f;
   wire [0:0] 				    c2h_gpio_1_gpio_29_f;
   wire [0:0] 				    c2h_gpio_1_gpio_28_f;
   wire [0:0] 				    c2h_gpio_1_gpio_27_f;
   wire [0:0] 				    c2h_gpio_1_gpio_26_f;
   wire [0:0] 				    c2h_gpio_1_gpio_25_f;
   wire [0:0] 				    c2h_gpio_1_gpio_24_f;
   wire [0:0] 				    c2h_gpio_1_gpio_23_f;
   wire [0:0] 				    c2h_gpio_1_gpio_22_f;
   wire [0:0] 				    c2h_gpio_1_gpio_21_f;
   wire [0:0] 				    c2h_gpio_1_gpio_20_f;
   wire [0:0] 				    c2h_gpio_1_gpio_19_f;
   wire [0:0] 				    c2h_gpio_1_gpio_18_f;
   wire [0:0] 				    c2h_gpio_1_gpio_17_f;
   wire [0:0] 				    c2h_gpio_1_gpio_16_f;
   wire [0:0] 				    c2h_gpio_1_gpio_15_f;
   wire [0:0] 				    c2h_gpio_1_gpio_14_f;
   wire [0:0] 				    c2h_gpio_1_gpio_13_f;
   wire [0:0] 				    c2h_gpio_1_gpio_12_f;
   wire [0:0] 				    c2h_gpio_1_gpio_11_f;
   wire [0:0] 				    c2h_gpio_1_gpio_10_f;
   wire [0:0] 				    c2h_gpio_1_gpio_9_f;
   wire [0:0] 				    c2h_gpio_1_gpio_8_f;
   wire [0:0] 				    c2h_gpio_1_gpio_7_f;
   wire [0:0] 				    c2h_gpio_1_gpio_6_f;
   wire [0:0] 				    c2h_gpio_1_gpio_5_f;
   wire [0:0] 				    c2h_gpio_1_gpio_4_f;
   wire [0:0] 				    c2h_gpio_1_gpio_3_f;
   wire [0:0] 				    c2h_gpio_1_gpio_2_f;
   wire [0:0] 				    c2h_gpio_1_gpio_1_f;
   wire [0:0] 				    c2h_gpio_1_gpio_0_f;
   wire [0:0] 				    c2h_gpio_2_gpio_31_f;
   wire [0:0] 				    c2h_gpio_2_gpio_30_f;
   wire [0:0] 				    c2h_gpio_2_gpio_29_f;
   wire [0:0] 				    c2h_gpio_2_gpio_28_f;
   wire [0:0] 				    c2h_gpio_2_gpio_27_f;
   wire [0:0] 				    c2h_gpio_2_gpio_26_f;
   wire [0:0] 				    c2h_gpio_2_gpio_25_f;
   wire [0:0] 				    c2h_gpio_2_gpio_24_f;
   wire [0:0] 				    c2h_gpio_2_gpio_23_f;
   wire [0:0] 				    c2h_gpio_2_gpio_22_f;
   wire [0:0] 				    c2h_gpio_2_gpio_21_f;
   wire [0:0] 				    c2h_gpio_2_gpio_20_f;
   wire [0:0] 				    c2h_gpio_2_gpio_19_f;
   wire [0:0] 				    c2h_gpio_2_gpio_18_f;
   wire [0:0] 				    c2h_gpio_2_gpio_17_f;
   wire [0:0] 				    c2h_gpio_2_gpio_16_f;
   wire [0:0] 				    c2h_gpio_2_gpio_15_f;
   wire [0:0] 				    c2h_gpio_2_gpio_14_f;
   wire [0:0] 				    c2h_gpio_2_gpio_13_f;
   wire [0:0] 				    c2h_gpio_2_gpio_12_f;
   wire [0:0] 				    c2h_gpio_2_gpio_11_f;
   wire [0:0] 				    c2h_gpio_2_gpio_10_f;
   wire [0:0] 				    c2h_gpio_2_gpio_9_f;
   wire [0:0] 				    c2h_gpio_2_gpio_8_f;
   wire [0:0] 				    c2h_gpio_2_gpio_7_f;
   wire [0:0] 				    c2h_gpio_2_gpio_6_f;
   wire [0:0] 				    c2h_gpio_2_gpio_5_f;
   wire [0:0] 				    c2h_gpio_2_gpio_4_f;
   wire [0:0] 				    c2h_gpio_2_gpio_3_f;
   wire [0:0] 				    c2h_gpio_2_gpio_2_f;
   wire [0:0] 				    c2h_gpio_2_gpio_1_f;
   wire [0:0] 				    c2h_gpio_2_gpio_0_f;
   wire [0:0] 				    c2h_gpio_3_gpio_31_f;
   wire [0:0] 				    c2h_gpio_3_gpio_30_f;
   wire [0:0] 				    c2h_gpio_3_gpio_29_f;
   wire [0:0] 				    c2h_gpio_3_gpio_28_f;
   wire [0:0] 				    c2h_gpio_3_gpio_27_f;
   wire [0:0] 				    c2h_gpio_3_gpio_26_f;
   wire [0:0] 				    c2h_gpio_3_gpio_25_f;
   wire [0:0] 				    c2h_gpio_3_gpio_24_f;
   wire [0:0] 				    c2h_gpio_3_gpio_23_f;
   wire [0:0] 				    c2h_gpio_3_gpio_22_f;
   wire [0:0] 				    c2h_gpio_3_gpio_21_f;
   wire [0:0] 				    c2h_gpio_3_gpio_20_f;
   wire [0:0] 				    c2h_gpio_3_gpio_19_f;
   wire [0:0] 				    c2h_gpio_3_gpio_18_f;
   wire [0:0] 				    c2h_gpio_3_gpio_17_f;
   wire [0:0] 				    c2h_gpio_3_gpio_16_f;
   wire [0:0] 				    c2h_gpio_3_gpio_15_f;
   wire [0:0] 				    c2h_gpio_3_gpio_14_f;
   wire [0:0] 				    c2h_gpio_3_gpio_13_f;
   wire [0:0] 				    c2h_gpio_3_gpio_12_f;
   wire [0:0] 				    c2h_gpio_3_gpio_11_f;
   wire [0:0] 				    c2h_gpio_3_gpio_10_f;
   wire [0:0] 				    c2h_gpio_3_gpio_9_f;
   wire [0:0] 				    c2h_gpio_3_gpio_8_f;
   wire [0:0] 				    c2h_gpio_3_gpio_7_f;
   wire [0:0] 				    c2h_gpio_3_gpio_6_f;
   wire [0:0] 				    c2h_gpio_3_gpio_5_f;
   wire [0:0] 				    c2h_gpio_3_gpio_4_f;
   wire [0:0] 				    c2h_gpio_3_gpio_3_f;
   wire [0:0] 				    c2h_gpio_3_gpio_2_f;
   wire [0:0] 				    c2h_gpio_3_gpio_1_f;
   wire [0:0] 				    c2h_gpio_3_gpio_0_f;
   wire [0:0] 				    c2h_gpio_4_gpio_31_f;
   wire [0:0] 				    c2h_gpio_4_gpio_30_f;
   wire [0:0] 				    c2h_gpio_4_gpio_29_f;
   wire [0:0] 				    c2h_gpio_4_gpio_28_f;
   wire [0:0] 				    c2h_gpio_4_gpio_27_f;
   wire [0:0] 				    c2h_gpio_4_gpio_26_f;
   wire [0:0] 				    c2h_gpio_4_gpio_25_f;
   wire [0:0] 				    c2h_gpio_4_gpio_24_f;
   wire [0:0] 				    c2h_gpio_4_gpio_23_f;
   wire [0:0] 				    c2h_gpio_4_gpio_22_f;
   wire [0:0] 				    c2h_gpio_4_gpio_21_f;
   wire [0:0] 				    c2h_gpio_4_gpio_20_f;
   wire [0:0] 				    c2h_gpio_4_gpio_19_f;
   wire [0:0] 				    c2h_gpio_4_gpio_18_f;
   wire [0:0] 				    c2h_gpio_4_gpio_17_f;
   wire [0:0] 				    c2h_gpio_4_gpio_16_f;
   wire [0:0] 				    c2h_gpio_4_gpio_15_f;
   wire [0:0] 				    c2h_gpio_4_gpio_14_f;
   wire [0:0] 				    c2h_gpio_4_gpio_13_f;
   wire [0:0] 				    c2h_gpio_4_gpio_12_f;
   wire [0:0] 				    c2h_gpio_4_gpio_11_f;
   wire [0:0] 				    c2h_gpio_4_gpio_10_f;
   wire [0:0] 				    c2h_gpio_4_gpio_9_f;
   wire [0:0] 				    c2h_gpio_4_gpio_8_f;
   wire [0:0] 				    c2h_gpio_4_gpio_7_f;
   wire [0:0] 				    c2h_gpio_4_gpio_6_f;
   wire [0:0] 				    c2h_gpio_4_gpio_5_f;
   wire [0:0] 				    c2h_gpio_4_gpio_4_f;
   wire [0:0] 				    c2h_gpio_4_gpio_3_f;
   wire [0:0] 				    c2h_gpio_4_gpio_2_f;
   wire [0:0] 				    c2h_gpio_4_gpio_1_f;
   wire [0:0] 				    c2h_gpio_4_gpio_0_f;
   wire [0:0] 				    c2h_gpio_5_gpio_31_f;
   wire [0:0] 				    c2h_gpio_5_gpio_30_f;
   wire [0:0] 				    c2h_gpio_5_gpio_29_f;
   wire [0:0] 				    c2h_gpio_5_gpio_28_f;
   wire [0:0] 				    c2h_gpio_5_gpio_27_f;
   wire [0:0] 				    c2h_gpio_5_gpio_26_f;
   wire [0:0] 				    c2h_gpio_5_gpio_25_f;
   wire [0:0] 				    c2h_gpio_5_gpio_24_f;
   wire [0:0] 				    c2h_gpio_5_gpio_23_f;
   wire [0:0] 				    c2h_gpio_5_gpio_22_f;
   wire [0:0] 				    c2h_gpio_5_gpio_21_f;
   wire [0:0] 				    c2h_gpio_5_gpio_20_f;
   wire [0:0] 				    c2h_gpio_5_gpio_19_f;
   wire [0:0] 				    c2h_gpio_5_gpio_18_f;
   wire [0:0] 				    c2h_gpio_5_gpio_17_f;
   wire [0:0] 				    c2h_gpio_5_gpio_16_f;
   wire [0:0] 				    c2h_gpio_5_gpio_15_f;
   wire [0:0] 				    c2h_gpio_5_gpio_14_f;
   wire [0:0] 				    c2h_gpio_5_gpio_13_f;
   wire [0:0] 				    c2h_gpio_5_gpio_12_f;
   wire [0:0] 				    c2h_gpio_5_gpio_11_f;
   wire [0:0] 				    c2h_gpio_5_gpio_10_f;
   wire [0:0] 				    c2h_gpio_5_gpio_9_f;
   wire [0:0] 				    c2h_gpio_5_gpio_8_f;
   wire [0:0] 				    c2h_gpio_5_gpio_7_f;
   wire [0:0] 				    c2h_gpio_5_gpio_6_f;
   wire [0:0] 				    c2h_gpio_5_gpio_5_f;
   wire [0:0] 				    c2h_gpio_5_gpio_4_f;
   wire [0:0] 				    c2h_gpio_5_gpio_3_f;
   wire [0:0] 				    c2h_gpio_5_gpio_2_f;
   wire [0:0] 				    c2h_gpio_5_gpio_1_f;
   wire [0:0] 				    c2h_gpio_5_gpio_0_f;
   wire [0:0] 				    c2h_gpio_6_gpio_31_f;
   wire [0:0] 				    c2h_gpio_6_gpio_30_f;
   wire [0:0] 				    c2h_gpio_6_gpio_29_f;
   wire [0:0] 				    c2h_gpio_6_gpio_28_f;
   wire [0:0] 				    c2h_gpio_6_gpio_27_f;
   wire [0:0] 				    c2h_gpio_6_gpio_26_f;
   wire [0:0] 				    c2h_gpio_6_gpio_25_f;
   wire [0:0] 				    c2h_gpio_6_gpio_24_f;
   wire [0:0] 				    c2h_gpio_6_gpio_23_f;
   wire [0:0] 				    c2h_gpio_6_gpio_22_f;
   wire [0:0] 				    c2h_gpio_6_gpio_21_f;
   wire [0:0] 				    c2h_gpio_6_gpio_20_f;
   wire [0:0] 				    c2h_gpio_6_gpio_19_f;
   wire [0:0] 				    c2h_gpio_6_gpio_18_f;
   wire [0:0] 				    c2h_gpio_6_gpio_17_f;
   wire [0:0] 				    c2h_gpio_6_gpio_16_f;
   wire [0:0] 				    c2h_gpio_6_gpio_15_f;
   wire [0:0] 				    c2h_gpio_6_gpio_14_f;
   wire [0:0] 				    c2h_gpio_6_gpio_13_f;
   wire [0:0] 				    c2h_gpio_6_gpio_12_f;
   wire [0:0] 				    c2h_gpio_6_gpio_11_f;
   wire [0:0] 				    c2h_gpio_6_gpio_10_f;
   wire [0:0] 				    c2h_gpio_6_gpio_9_f;
   wire [0:0] 				    c2h_gpio_6_gpio_8_f;
   wire [0:0] 				    c2h_gpio_6_gpio_7_f;
   wire [0:0] 				    c2h_gpio_6_gpio_6_f;
   wire [0:0] 				    c2h_gpio_6_gpio_5_f;
   wire [0:0] 				    c2h_gpio_6_gpio_4_f;
   wire [0:0] 				    c2h_gpio_6_gpio_3_f;
   wire [0:0] 				    c2h_gpio_6_gpio_2_f;
   wire [0:0] 				    c2h_gpio_6_gpio_1_f;
   wire [0:0] 				    c2h_gpio_6_gpio_0_f;
   wire [0:0] 				    c2h_gpio_7_gpio_31_f;
   wire [0:0] 				    c2h_gpio_7_gpio_30_f;
   wire [0:0] 				    c2h_gpio_7_gpio_29_f;
   wire [0:0] 				    c2h_gpio_7_gpio_28_f;
   wire [0:0] 				    c2h_gpio_7_gpio_27_f;
   wire [0:0] 				    c2h_gpio_7_gpio_26_f;
   wire [0:0] 				    c2h_gpio_7_gpio_25_f;
   wire [0:0] 				    c2h_gpio_7_gpio_24_f;
   wire [0:0] 				    c2h_gpio_7_gpio_23_f;
   wire [0:0] 				    c2h_gpio_7_gpio_22_f;
   wire [0:0] 				    c2h_gpio_7_gpio_21_f;
   wire [0:0] 				    c2h_gpio_7_gpio_20_f;
   wire [0:0] 				    c2h_gpio_7_gpio_19_f;
   wire [0:0] 				    c2h_gpio_7_gpio_18_f;
   wire [0:0] 				    c2h_gpio_7_gpio_17_f;
   wire [0:0] 				    c2h_gpio_7_gpio_16_f;
   wire [0:0] 				    c2h_gpio_7_gpio_15_f;
   wire [0:0] 				    c2h_gpio_7_gpio_14_f;
   wire [0:0] 				    c2h_gpio_7_gpio_13_f;
   wire [0:0] 				    c2h_gpio_7_gpio_12_f;
   wire [0:0] 				    c2h_gpio_7_gpio_11_f;
   wire [0:0] 				    c2h_gpio_7_gpio_10_f;
   wire [0:0] 				    c2h_gpio_7_gpio_9_f;
   wire [0:0] 				    c2h_gpio_7_gpio_8_f;
   wire [0:0] 				    c2h_gpio_7_gpio_7_f;
   wire [0:0] 				    c2h_gpio_7_gpio_6_f;
   wire [0:0] 				    c2h_gpio_7_gpio_5_f;
   wire [0:0] 				    c2h_gpio_7_gpio_4_f;
   wire [0:0] 				    c2h_gpio_7_gpio_3_f;
   wire [0:0] 				    c2h_gpio_7_gpio_2_f;
   wire [0:0] 				    c2h_gpio_7_gpio_1_f;
   wire [0:0] 				    c2h_gpio_7_gpio_0_f;
   wire [0:0] 				    c2h_gpio_8_gpio_31_f;
   wire [0:0] 				    c2h_gpio_8_gpio_30_f;
   wire [0:0] 				    c2h_gpio_8_gpio_29_f;
   wire [0:0] 				    c2h_gpio_8_gpio_28_f;
   wire [0:0] 				    c2h_gpio_8_gpio_27_f;
   wire [0:0] 				    c2h_gpio_8_gpio_26_f;
   wire [0:0] 				    c2h_gpio_8_gpio_25_f;
   wire [0:0] 				    c2h_gpio_8_gpio_24_f;
   wire [0:0] 				    c2h_gpio_8_gpio_23_f;
   wire [0:0] 				    c2h_gpio_8_gpio_22_f;
   wire [0:0] 				    c2h_gpio_8_gpio_21_f;
   wire [0:0] 				    c2h_gpio_8_gpio_20_f;
   wire [0:0] 				    c2h_gpio_8_gpio_19_f;
   wire [0:0] 				    c2h_gpio_8_gpio_18_f;
   wire [0:0] 				    c2h_gpio_8_gpio_17_f;
   wire [0:0] 				    c2h_gpio_8_gpio_16_f;
   wire [0:0] 				    c2h_gpio_8_gpio_15_f;
   wire [0:0] 				    c2h_gpio_8_gpio_14_f;
   wire [0:0] 				    c2h_gpio_8_gpio_13_f;
   wire [0:0] 				    c2h_gpio_8_gpio_12_f;
   wire [0:0] 				    c2h_gpio_8_gpio_11_f;
   wire [0:0] 				    c2h_gpio_8_gpio_10_f;
   wire [0:0] 				    c2h_gpio_8_gpio_9_f;
   wire [0:0] 				    c2h_gpio_8_gpio_8_f;
   wire [0:0] 				    c2h_gpio_8_gpio_7_f;
   wire [0:0] 				    c2h_gpio_8_gpio_6_f;
   wire [0:0] 				    c2h_gpio_8_gpio_5_f;
   wire [0:0] 				    c2h_gpio_8_gpio_4_f;
   wire [0:0] 				    c2h_gpio_8_gpio_3_f;
   wire [0:0] 				    c2h_gpio_8_gpio_2_f;
   wire [0:0] 				    c2h_gpio_8_gpio_1_f;
   wire [0:0] 				    c2h_gpio_8_gpio_0_f;
   wire [0:0] 				    c2h_gpio_9_gpio_31_f;
   wire [0:0] 				    c2h_gpio_9_gpio_30_f;
   wire [0:0] 				    c2h_gpio_9_gpio_29_f;
   wire [0:0] 				    c2h_gpio_9_gpio_28_f;
   wire [0:0] 				    c2h_gpio_9_gpio_27_f;
   wire [0:0] 				    c2h_gpio_9_gpio_26_f;
   wire [0:0] 				    c2h_gpio_9_gpio_25_f;
   wire [0:0] 				    c2h_gpio_9_gpio_24_f;
   wire [0:0] 				    c2h_gpio_9_gpio_23_f;
   wire [0:0] 				    c2h_gpio_9_gpio_22_f;
   wire [0:0] 				    c2h_gpio_9_gpio_21_f;
   wire [0:0] 				    c2h_gpio_9_gpio_20_f;
   wire [0:0] 				    c2h_gpio_9_gpio_19_f;
   wire [0:0] 				    c2h_gpio_9_gpio_18_f;
   wire [0:0] 				    c2h_gpio_9_gpio_17_f;
   wire [0:0] 				    c2h_gpio_9_gpio_16_f;
   wire [0:0] 				    c2h_gpio_9_gpio_15_f;
   wire [0:0] 				    c2h_gpio_9_gpio_14_f;
   wire [0:0] 				    c2h_gpio_9_gpio_13_f;
   wire [0:0] 				    c2h_gpio_9_gpio_12_f;
   wire [0:0] 				    c2h_gpio_9_gpio_11_f;
   wire [0:0] 				    c2h_gpio_9_gpio_10_f;
   wire [0:0] 				    c2h_gpio_9_gpio_9_f;
   wire [0:0] 				    c2h_gpio_9_gpio_8_f;
   wire [0:0] 				    c2h_gpio_9_gpio_7_f;
   wire [0:0] 				    c2h_gpio_9_gpio_6_f;
   wire [0:0] 				    c2h_gpio_9_gpio_5_f;
   wire [0:0] 				    c2h_gpio_9_gpio_4_f;
   wire [0:0] 				    c2h_gpio_9_gpio_3_f;
   wire [0:0] 				    c2h_gpio_9_gpio_2_f;
   wire [0:0] 				    c2h_gpio_9_gpio_1_f;
   wire [0:0] 				    c2h_gpio_9_gpio_0_f;
   wire [0:0] 				    c2h_gpio_10_gpio_31_f;
   wire [0:0] 				    c2h_gpio_10_gpio_30_f;
   wire [0:0] 				    c2h_gpio_10_gpio_29_f;
   wire [0:0] 				    c2h_gpio_10_gpio_28_f;
   wire [0:0] 				    c2h_gpio_10_gpio_27_f;
   wire [0:0] 				    c2h_gpio_10_gpio_26_f;
   wire [0:0] 				    c2h_gpio_10_gpio_25_f;
   wire [0:0] 				    c2h_gpio_10_gpio_24_f;
   wire [0:0] 				    c2h_gpio_10_gpio_23_f;
   wire [0:0] 				    c2h_gpio_10_gpio_22_f;
   wire [0:0] 				    c2h_gpio_10_gpio_21_f;
   wire [0:0] 				    c2h_gpio_10_gpio_20_f;
   wire [0:0] 				    c2h_gpio_10_gpio_19_f;
   wire [0:0] 				    c2h_gpio_10_gpio_18_f;
   wire [0:0] 				    c2h_gpio_10_gpio_17_f;
   wire [0:0] 				    c2h_gpio_10_gpio_16_f;
   wire [0:0] 				    c2h_gpio_10_gpio_15_f;
   wire [0:0] 				    c2h_gpio_10_gpio_14_f;
   wire [0:0] 				    c2h_gpio_10_gpio_13_f;
   wire [0:0] 				    c2h_gpio_10_gpio_12_f;
   wire [0:0] 				    c2h_gpio_10_gpio_11_f;
   wire [0:0] 				    c2h_gpio_10_gpio_10_f;
   wire [0:0] 				    c2h_gpio_10_gpio_9_f;
   wire [0:0] 				    c2h_gpio_10_gpio_8_f;
   wire [0:0] 				    c2h_gpio_10_gpio_7_f;
   wire [0:0] 				    c2h_gpio_10_gpio_6_f;
   wire [0:0] 				    c2h_gpio_10_gpio_5_f;
   wire [0:0] 				    c2h_gpio_10_gpio_4_f;
   wire [0:0] 				    c2h_gpio_10_gpio_3_f;
   wire [0:0] 				    c2h_gpio_10_gpio_2_f;
   wire [0:0] 				    c2h_gpio_10_gpio_1_f;
   wire [0:0] 				    c2h_gpio_10_gpio_0_f;
   wire [0:0] 				    c2h_gpio_11_gpio_31_f;
   wire [0:0] 				    c2h_gpio_11_gpio_30_f;
   wire [0:0] 				    c2h_gpio_11_gpio_29_f;
   wire [0:0] 				    c2h_gpio_11_gpio_28_f;
   wire [0:0] 				    c2h_gpio_11_gpio_27_f;
   wire [0:0] 				    c2h_gpio_11_gpio_26_f;
   wire [0:0] 				    c2h_gpio_11_gpio_25_f;
   wire [0:0] 				    c2h_gpio_11_gpio_24_f;
   wire [0:0] 				    c2h_gpio_11_gpio_23_f;
   wire [0:0] 				    c2h_gpio_11_gpio_22_f;
   wire [0:0] 				    c2h_gpio_11_gpio_21_f;
   wire [0:0] 				    c2h_gpio_11_gpio_20_f;
   wire [0:0] 				    c2h_gpio_11_gpio_19_f;
   wire [0:0] 				    c2h_gpio_11_gpio_18_f;
   wire [0:0] 				    c2h_gpio_11_gpio_17_f;
   wire [0:0] 				    c2h_gpio_11_gpio_16_f;
   wire [0:0] 				    c2h_gpio_11_gpio_15_f;
   wire [0:0] 				    c2h_gpio_11_gpio_14_f;
   wire [0:0] 				    c2h_gpio_11_gpio_13_f;
   wire [0:0] 				    c2h_gpio_11_gpio_12_f;
   wire [0:0] 				    c2h_gpio_11_gpio_11_f;
   wire [0:0] 				    c2h_gpio_11_gpio_10_f;
   wire [0:0] 				    c2h_gpio_11_gpio_9_f;
   wire [0:0] 				    c2h_gpio_11_gpio_8_f;
   wire [0:0] 				    c2h_gpio_11_gpio_7_f;
   wire [0:0] 				    c2h_gpio_11_gpio_6_f;
   wire [0:0] 				    c2h_gpio_11_gpio_5_f;
   wire [0:0] 				    c2h_gpio_11_gpio_4_f;
   wire [0:0] 				    c2h_gpio_11_gpio_3_f;
   wire [0:0] 				    c2h_gpio_11_gpio_2_f;
   wire [0:0] 				    c2h_gpio_11_gpio_1_f;
   wire [0:0] 				    c2h_gpio_11_gpio_0_f;
   wire [0:0] 				    c2h_gpio_12_gpio_31_f;
   wire [0:0] 				    c2h_gpio_12_gpio_30_f;
   wire [0:0] 				    c2h_gpio_12_gpio_29_f;
   wire [0:0] 				    c2h_gpio_12_gpio_28_f;
   wire [0:0] 				    c2h_gpio_12_gpio_27_f;
   wire [0:0] 				    c2h_gpio_12_gpio_26_f;
   wire [0:0] 				    c2h_gpio_12_gpio_25_f;
   wire [0:0] 				    c2h_gpio_12_gpio_24_f;
   wire [0:0] 				    c2h_gpio_12_gpio_23_f;
   wire [0:0] 				    c2h_gpio_12_gpio_22_f;
   wire [0:0] 				    c2h_gpio_12_gpio_21_f;
   wire [0:0] 				    c2h_gpio_12_gpio_20_f;
   wire [0:0] 				    c2h_gpio_12_gpio_19_f;
   wire [0:0] 				    c2h_gpio_12_gpio_18_f;
   wire [0:0] 				    c2h_gpio_12_gpio_17_f;
   wire [0:0] 				    c2h_gpio_12_gpio_16_f;
   wire [0:0] 				    c2h_gpio_12_gpio_15_f;
   wire [0:0] 				    c2h_gpio_12_gpio_14_f;
   wire [0:0] 				    c2h_gpio_12_gpio_13_f;
   wire [0:0] 				    c2h_gpio_12_gpio_12_f;
   wire [0:0] 				    c2h_gpio_12_gpio_11_f;
   wire [0:0] 				    c2h_gpio_12_gpio_10_f;
   wire [0:0] 				    c2h_gpio_12_gpio_9_f;
   wire [0:0] 				    c2h_gpio_12_gpio_8_f;
   wire [0:0] 				    c2h_gpio_12_gpio_7_f;
   wire [0:0] 				    c2h_gpio_12_gpio_6_f;
   wire [0:0] 				    c2h_gpio_12_gpio_5_f;
   wire [0:0] 				    c2h_gpio_12_gpio_4_f;
   wire [0:0] 				    c2h_gpio_12_gpio_3_f;
   wire [0:0] 				    c2h_gpio_12_gpio_2_f;
   wire [0:0] 				    c2h_gpio_12_gpio_1_f;
   wire [0:0] 				    c2h_gpio_12_gpio_0_f;
   wire [0:0] 				    c2h_gpio_13_gpio_31_f;
   wire [0:0] 				    c2h_gpio_13_gpio_30_f;
   wire [0:0] 				    c2h_gpio_13_gpio_29_f;
   wire [0:0] 				    c2h_gpio_13_gpio_28_f;
   wire [0:0] 				    c2h_gpio_13_gpio_27_f;
   wire [0:0] 				    c2h_gpio_13_gpio_26_f;
   wire [0:0] 				    c2h_gpio_13_gpio_25_f;
   wire [0:0] 				    c2h_gpio_13_gpio_24_f;
   wire [0:0] 				    c2h_gpio_13_gpio_23_f;
   wire [0:0] 				    c2h_gpio_13_gpio_22_f;
   wire [0:0] 				    c2h_gpio_13_gpio_21_f;
   wire [0:0] 				    c2h_gpio_13_gpio_20_f;
   wire [0:0] 				    c2h_gpio_13_gpio_19_f;
   wire [0:0] 				    c2h_gpio_13_gpio_18_f;
   wire [0:0] 				    c2h_gpio_13_gpio_17_f;
   wire [0:0] 				    c2h_gpio_13_gpio_16_f;
   wire [0:0] 				    c2h_gpio_13_gpio_15_f;
   wire [0:0] 				    c2h_gpio_13_gpio_14_f;
   wire [0:0] 				    c2h_gpio_13_gpio_13_f;
   wire [0:0] 				    c2h_gpio_13_gpio_12_f;
   wire [0:0] 				    c2h_gpio_13_gpio_11_f;
   wire [0:0] 				    c2h_gpio_13_gpio_10_f;
   wire [0:0] 				    c2h_gpio_13_gpio_9_f;
   wire [0:0] 				    c2h_gpio_13_gpio_8_f;
   wire [0:0] 				    c2h_gpio_13_gpio_7_f;
   wire [0:0] 				    c2h_gpio_13_gpio_6_f;
   wire [0:0] 				    c2h_gpio_13_gpio_5_f;
   wire [0:0] 				    c2h_gpio_13_gpio_4_f;
   wire [0:0] 				    c2h_gpio_13_gpio_3_f;
   wire [0:0] 				    c2h_gpio_13_gpio_2_f;
   wire [0:0] 				    c2h_gpio_13_gpio_1_f;
   wire [0:0] 				    c2h_gpio_13_gpio_0_f;
   wire [0:0] 				    c2h_gpio_14_gpio_31_f;
   wire [0:0] 				    c2h_gpio_14_gpio_30_f;
   wire [0:0] 				    c2h_gpio_14_gpio_29_f;
   wire [0:0] 				    c2h_gpio_14_gpio_28_f;
   wire [0:0] 				    c2h_gpio_14_gpio_27_f;
   wire [0:0] 				    c2h_gpio_14_gpio_26_f;
   wire [0:0] 				    c2h_gpio_14_gpio_25_f;
   wire [0:0] 				    c2h_gpio_14_gpio_24_f;
   wire [0:0] 				    c2h_gpio_14_gpio_23_f;
   wire [0:0] 				    c2h_gpio_14_gpio_22_f;
   wire [0:0] 				    c2h_gpio_14_gpio_21_f;
   wire [0:0] 				    c2h_gpio_14_gpio_20_f;
   wire [0:0] 				    c2h_gpio_14_gpio_19_f;
   wire [0:0] 				    c2h_gpio_14_gpio_18_f;
   wire [0:0] 				    c2h_gpio_14_gpio_17_f;
   wire [0:0] 				    c2h_gpio_14_gpio_16_f;
   wire [0:0] 				    c2h_gpio_14_gpio_15_f;
   wire [0:0] 				    c2h_gpio_14_gpio_14_f;
   wire [0:0] 				    c2h_gpio_14_gpio_13_f;
   wire [0:0] 				    c2h_gpio_14_gpio_12_f;
   wire [0:0] 				    c2h_gpio_14_gpio_11_f;
   wire [0:0] 				    c2h_gpio_14_gpio_10_f;
   wire [0:0] 				    c2h_gpio_14_gpio_9_f;
   wire [0:0] 				    c2h_gpio_14_gpio_8_f;
   wire [0:0] 				    c2h_gpio_14_gpio_7_f;
   wire [0:0] 				    c2h_gpio_14_gpio_6_f;
   wire [0:0] 				    c2h_gpio_14_gpio_5_f;
   wire [0:0] 				    c2h_gpio_14_gpio_4_f;
   wire [0:0] 				    c2h_gpio_14_gpio_3_f;
   wire [0:0] 				    c2h_gpio_14_gpio_2_f;
   wire [0:0] 				    c2h_gpio_14_gpio_1_f;
   wire [0:0] 				    c2h_gpio_14_gpio_0_f;
   wire [0:0] 				    c2h_gpio_15_gpio_31_f;
   wire [0:0] 				    c2h_gpio_15_gpio_30_f;
   wire [0:0] 				    c2h_gpio_15_gpio_29_f;
   wire [0:0] 				    c2h_gpio_15_gpio_28_f;
   wire [0:0] 				    c2h_gpio_15_gpio_27_f;
   wire [0:0] 				    c2h_gpio_15_gpio_26_f;
   wire [0:0] 				    c2h_gpio_15_gpio_25_f;
   wire [0:0] 				    c2h_gpio_15_gpio_24_f;
   wire [0:0] 				    c2h_gpio_15_gpio_23_f;
   wire [0:0] 				    c2h_gpio_15_gpio_22_f;
   wire [0:0] 				    c2h_gpio_15_gpio_21_f;
   wire [0:0] 				    c2h_gpio_15_gpio_20_f;
   wire [0:0] 				    c2h_gpio_15_gpio_19_f;
   wire [0:0] 				    c2h_gpio_15_gpio_18_f;
   wire [0:0] 				    c2h_gpio_15_gpio_17_f;
   wire [0:0] 				    c2h_gpio_15_gpio_16_f;
   wire [0:0] 				    c2h_gpio_15_gpio_15_f;
   wire [0:0] 				    c2h_gpio_15_gpio_14_f;
   wire [0:0] 				    c2h_gpio_15_gpio_13_f;
   wire [0:0] 				    c2h_gpio_15_gpio_12_f;
   wire [0:0] 				    c2h_gpio_15_gpio_11_f;
   wire [0:0] 				    c2h_gpio_15_gpio_10_f;
   wire [0:0] 				    c2h_gpio_15_gpio_9_f;
   wire [0:0] 				    c2h_gpio_15_gpio_8_f;
   wire [0:0] 				    c2h_gpio_15_gpio_7_f;
   wire [0:0] 				    c2h_gpio_15_gpio_6_f;
   wire [0:0] 				    c2h_gpio_15_gpio_5_f;
   wire [0:0] 				    c2h_gpio_15_gpio_4_f;
   wire [0:0] 				    c2h_gpio_15_gpio_3_f;
   wire [0:0] 				    c2h_gpio_15_gpio_2_f;
   wire [0:0] 				    c2h_gpio_15_gpio_1_f;
   wire [0:0] 				    c2h_gpio_15_gpio_0_f;
   wire [0:0] 				    h2c_gpio_0_gpio_31_f;
   wire [0:0] 				    h2c_gpio_0_gpio_30_f;
   wire [0:0] 				    h2c_gpio_0_gpio_29_f;
   wire [0:0] 				    h2c_gpio_0_gpio_28_f;
   wire [0:0] 				    h2c_gpio_0_gpio_27_f;
   wire [0:0] 				    h2c_gpio_0_gpio_26_f;
   wire [0:0] 				    h2c_gpio_0_gpio_25_f;
   wire [0:0] 				    h2c_gpio_0_gpio_24_f;
   wire [0:0] 				    h2c_gpio_0_gpio_23_f;
   wire [0:0] 				    h2c_gpio_0_gpio_22_f;
   wire [0:0] 				    h2c_gpio_0_gpio_21_f;
   wire [0:0] 				    h2c_gpio_0_gpio_20_f;
   wire [0:0] 				    h2c_gpio_0_gpio_19_f;
   wire [0:0] 				    h2c_gpio_0_gpio_18_f;
   wire [0:0] 				    h2c_gpio_0_gpio_17_f;
   wire [0:0] 				    h2c_gpio_0_gpio_16_f;
   wire [0:0] 				    h2c_gpio_0_gpio_15_f;
   wire [0:0] 				    h2c_gpio_0_gpio_14_f;
   wire [0:0] 				    h2c_gpio_0_gpio_13_f;
   wire [0:0] 				    h2c_gpio_0_gpio_12_f;
   wire [0:0] 				    h2c_gpio_0_gpio_11_f;
   wire [0:0] 				    h2c_gpio_0_gpio_10_f;
   wire [0:0] 				    h2c_gpio_0_gpio_9_f;
   wire [0:0] 				    h2c_gpio_0_gpio_8_f;
   wire [0:0] 				    h2c_gpio_0_gpio_7_f;
   wire [0:0] 				    h2c_gpio_0_gpio_6_f;
   wire [0:0] 				    h2c_gpio_0_gpio_5_f;
   wire [0:0] 				    h2c_gpio_0_gpio_4_f;
   wire [0:0] 				    h2c_gpio_0_gpio_3_f;
   wire [0:0] 				    h2c_gpio_0_gpio_2_f;
   wire [0:0] 				    h2c_gpio_0_gpio_1_f;
   wire [0:0] 				    h2c_gpio_0_gpio_0_f;
   wire [0:0] 				    h2c_gpio_1_gpio_31_f;
   wire [0:0] 				    h2c_gpio_1_gpio_30_f;
   wire [0:0] 				    h2c_gpio_1_gpio_29_f;
   wire [0:0] 				    h2c_gpio_1_gpio_28_f;
   wire [0:0] 				    h2c_gpio_1_gpio_27_f;
   wire [0:0] 				    h2c_gpio_1_gpio_26_f;
   wire [0:0] 				    h2c_gpio_1_gpio_25_f;
   wire [0:0] 				    h2c_gpio_1_gpio_24_f;
   wire [0:0] 				    h2c_gpio_1_gpio_23_f;
   wire [0:0] 				    h2c_gpio_1_gpio_22_f;
   wire [0:0] 				    h2c_gpio_1_gpio_21_f;
   wire [0:0] 				    h2c_gpio_1_gpio_20_f;
   wire [0:0] 				    h2c_gpio_1_gpio_19_f;
   wire [0:0] 				    h2c_gpio_1_gpio_18_f;
   wire [0:0] 				    h2c_gpio_1_gpio_17_f;
   wire [0:0] 				    h2c_gpio_1_gpio_16_f;
   wire [0:0] 				    h2c_gpio_1_gpio_15_f;
   wire [0:0] 				    h2c_gpio_1_gpio_14_f;
   wire [0:0] 				    h2c_gpio_1_gpio_13_f;
   wire [0:0] 				    h2c_gpio_1_gpio_12_f;
   wire [0:0] 				    h2c_gpio_1_gpio_11_f;
   wire [0:0] 				    h2c_gpio_1_gpio_10_f;
   wire [0:0] 				    h2c_gpio_1_gpio_9_f;
   wire [0:0] 				    h2c_gpio_1_gpio_8_f;
   wire [0:0] 				    h2c_gpio_1_gpio_7_f;
   wire [0:0] 				    h2c_gpio_1_gpio_6_f;
   wire [0:0] 				    h2c_gpio_1_gpio_5_f;
   wire [0:0] 				    h2c_gpio_1_gpio_4_f;
   wire [0:0] 				    h2c_gpio_1_gpio_3_f;
   wire [0:0] 				    h2c_gpio_1_gpio_2_f;
   wire [0:0] 				    h2c_gpio_1_gpio_1_f;
   wire [0:0] 				    h2c_gpio_1_gpio_0_f;
   wire [0:0] 				    h2c_gpio_2_gpio_31_f;
   wire [0:0] 				    h2c_gpio_2_gpio_30_f;
   wire [0:0] 				    h2c_gpio_2_gpio_29_f;
   wire [0:0] 				    h2c_gpio_2_gpio_28_f;
   wire [0:0] 				    h2c_gpio_2_gpio_27_f;
   wire [0:0] 				    h2c_gpio_2_gpio_26_f;
   wire [0:0] 				    h2c_gpio_2_gpio_25_f;
   wire [0:0] 				    h2c_gpio_2_gpio_24_f;
   wire [0:0] 				    h2c_gpio_2_gpio_23_f;
   wire [0:0] 				    h2c_gpio_2_gpio_22_f;
   wire [0:0] 				    h2c_gpio_2_gpio_21_f;
   wire [0:0] 				    h2c_gpio_2_gpio_20_f;
   wire [0:0] 				    h2c_gpio_2_gpio_19_f;
   wire [0:0] 				    h2c_gpio_2_gpio_18_f;
   wire [0:0] 				    h2c_gpio_2_gpio_17_f;
   wire [0:0] 				    h2c_gpio_2_gpio_16_f;
   wire [0:0] 				    h2c_gpio_2_gpio_15_f;
   wire [0:0] 				    h2c_gpio_2_gpio_14_f;
   wire [0:0] 				    h2c_gpio_2_gpio_13_f;
   wire [0:0] 				    h2c_gpio_2_gpio_12_f;
   wire [0:0] 				    h2c_gpio_2_gpio_11_f;
   wire [0:0] 				    h2c_gpio_2_gpio_10_f;
   wire [0:0] 				    h2c_gpio_2_gpio_9_f;
   wire [0:0] 				    h2c_gpio_2_gpio_8_f;
   wire [0:0] 				    h2c_gpio_2_gpio_7_f;
   wire [0:0] 				    h2c_gpio_2_gpio_6_f;
   wire [0:0] 				    h2c_gpio_2_gpio_5_f;
   wire [0:0] 				    h2c_gpio_2_gpio_4_f;
   wire [0:0] 				    h2c_gpio_2_gpio_3_f;
   wire [0:0] 				    h2c_gpio_2_gpio_2_f;
   wire [0:0] 				    h2c_gpio_2_gpio_1_f;
   wire [0:0] 				    h2c_gpio_2_gpio_0_f;
   wire [0:0] 				    h2c_gpio_3_gpio_31_f;
   wire [0:0] 				    h2c_gpio_3_gpio_30_f;
   wire [0:0] 				    h2c_gpio_3_gpio_29_f;
   wire [0:0] 				    h2c_gpio_3_gpio_28_f;
   wire [0:0] 				    h2c_gpio_3_gpio_27_f;
   wire [0:0] 				    h2c_gpio_3_gpio_26_f;
   wire [0:0] 				    h2c_gpio_3_gpio_25_f;
   wire [0:0] 				    h2c_gpio_3_gpio_24_f;
   wire [0:0] 				    h2c_gpio_3_gpio_23_f;
   wire [0:0] 				    h2c_gpio_3_gpio_22_f;
   wire [0:0] 				    h2c_gpio_3_gpio_21_f;
   wire [0:0] 				    h2c_gpio_3_gpio_20_f;
   wire [0:0] 				    h2c_gpio_3_gpio_19_f;
   wire [0:0] 				    h2c_gpio_3_gpio_18_f;
   wire [0:0] 				    h2c_gpio_3_gpio_17_f;
   wire [0:0] 				    h2c_gpio_3_gpio_16_f;
   wire [0:0] 				    h2c_gpio_3_gpio_15_f;
   wire [0:0] 				    h2c_gpio_3_gpio_14_f;
   wire [0:0] 				    h2c_gpio_3_gpio_13_f;
   wire [0:0] 				    h2c_gpio_3_gpio_12_f;
   wire [0:0] 				    h2c_gpio_3_gpio_11_f;
   wire [0:0] 				    h2c_gpio_3_gpio_10_f;
   wire [0:0] 				    h2c_gpio_3_gpio_9_f;
   wire [0:0] 				    h2c_gpio_3_gpio_8_f;
   wire [0:0] 				    h2c_gpio_3_gpio_7_f;
   wire [0:0] 				    h2c_gpio_3_gpio_6_f;
   wire [0:0] 				    h2c_gpio_3_gpio_5_f;
   wire [0:0] 				    h2c_gpio_3_gpio_4_f;
   wire [0:0] 				    h2c_gpio_3_gpio_3_f;
   wire [0:0] 				    h2c_gpio_3_gpio_2_f;
   wire [0:0] 				    h2c_gpio_3_gpio_1_f;
   wire [0:0] 				    h2c_gpio_3_gpio_0_f;
   wire [0:0] 				    h2c_gpio_4_gpio_31_f;
   wire [0:0] 				    h2c_gpio_4_gpio_30_f;
   wire [0:0] 				    h2c_gpio_4_gpio_29_f;
   wire [0:0] 				    h2c_gpio_4_gpio_28_f;
   wire [0:0] 				    h2c_gpio_4_gpio_27_f;
   wire [0:0] 				    h2c_gpio_4_gpio_26_f;
   wire [0:0] 				    h2c_gpio_4_gpio_25_f;
   wire [0:0] 				    h2c_gpio_4_gpio_24_f;
   wire [0:0] 				    h2c_gpio_4_gpio_23_f;
   wire [0:0] 				    h2c_gpio_4_gpio_22_f;
   wire [0:0] 				    h2c_gpio_4_gpio_21_f;
   wire [0:0] 				    h2c_gpio_4_gpio_20_f;
   wire [0:0] 				    h2c_gpio_4_gpio_19_f;
   wire [0:0] 				    h2c_gpio_4_gpio_18_f;
   wire [0:0] 				    h2c_gpio_4_gpio_17_f;
   wire [0:0] 				    h2c_gpio_4_gpio_16_f;
   wire [0:0] 				    h2c_gpio_4_gpio_15_f;
   wire [0:0] 				    h2c_gpio_4_gpio_14_f;
   wire [0:0] 				    h2c_gpio_4_gpio_13_f;
   wire [0:0] 				    h2c_gpio_4_gpio_12_f;
   wire [0:0] 				    h2c_gpio_4_gpio_11_f;
   wire [0:0] 				    h2c_gpio_4_gpio_10_f;
   wire [0:0] 				    h2c_gpio_4_gpio_9_f;
   wire [0:0] 				    h2c_gpio_4_gpio_8_f;
   wire [0:0] 				    h2c_gpio_4_gpio_7_f;
   wire [0:0] 				    h2c_gpio_4_gpio_6_f;
   wire [0:0] 				    h2c_gpio_4_gpio_5_f;
   wire [0:0] 				    h2c_gpio_4_gpio_4_f;
   wire [0:0] 				    h2c_gpio_4_gpio_3_f;
   wire [0:0] 				    h2c_gpio_4_gpio_2_f;
   wire [0:0] 				    h2c_gpio_4_gpio_1_f;
   wire [0:0] 				    h2c_gpio_4_gpio_0_f;
   wire [0:0] 				    h2c_gpio_5_gpio_31_f;
   wire [0:0] 				    h2c_gpio_5_gpio_30_f;
   wire [0:0] 				    h2c_gpio_5_gpio_29_f;
   wire [0:0] 				    h2c_gpio_5_gpio_28_f;
   wire [0:0] 				    h2c_gpio_5_gpio_27_f;
   wire [0:0] 				    h2c_gpio_5_gpio_26_f;
   wire [0:0] 				    h2c_gpio_5_gpio_25_f;
   wire [0:0] 				    h2c_gpio_5_gpio_24_f;
   wire [0:0] 				    h2c_gpio_5_gpio_23_f;
   wire [0:0] 				    h2c_gpio_5_gpio_22_f;
   wire [0:0] 				    h2c_gpio_5_gpio_21_f;
   wire [0:0] 				    h2c_gpio_5_gpio_20_f;
   wire [0:0] 				    h2c_gpio_5_gpio_19_f;
   wire [0:0] 				    h2c_gpio_5_gpio_18_f;
   wire [0:0] 				    h2c_gpio_5_gpio_17_f;
   wire [0:0] 				    h2c_gpio_5_gpio_16_f;
   wire [0:0] 				    h2c_gpio_5_gpio_15_f;
   wire [0:0] 				    h2c_gpio_5_gpio_14_f;
   wire [0:0] 				    h2c_gpio_5_gpio_13_f;
   wire [0:0] 				    h2c_gpio_5_gpio_12_f;
   wire [0:0] 				    h2c_gpio_5_gpio_11_f;
   wire [0:0] 				    h2c_gpio_5_gpio_10_f;
   wire [0:0] 				    h2c_gpio_5_gpio_9_f;
   wire [0:0] 				    h2c_gpio_5_gpio_8_f;
   wire [0:0] 				    h2c_gpio_5_gpio_7_f;
   wire [0:0] 				    h2c_gpio_5_gpio_6_f;
   wire [0:0] 				    h2c_gpio_5_gpio_5_f;
   wire [0:0] 				    h2c_gpio_5_gpio_4_f;
   wire [0:0] 				    h2c_gpio_5_gpio_3_f;
   wire [0:0] 				    h2c_gpio_5_gpio_2_f;
   wire [0:0] 				    h2c_gpio_5_gpio_1_f;
   wire [0:0] 				    h2c_gpio_5_gpio_0_f;
   wire [0:0] 				    h2c_gpio_6_gpio_31_f;
   wire [0:0] 				    h2c_gpio_6_gpio_30_f;
   wire [0:0] 				    h2c_gpio_6_gpio_29_f;
   wire [0:0] 				    h2c_gpio_6_gpio_28_f;
   wire [0:0] 				    h2c_gpio_6_gpio_27_f;
   wire [0:0] 				    h2c_gpio_6_gpio_26_f;
   wire [0:0] 				    h2c_gpio_6_gpio_25_f;
   wire [0:0] 				    h2c_gpio_6_gpio_24_f;
   wire [0:0] 				    h2c_gpio_6_gpio_23_f;
   wire [0:0] 				    h2c_gpio_6_gpio_22_f;
   wire [0:0] 				    h2c_gpio_6_gpio_21_f;
   wire [0:0] 				    h2c_gpio_6_gpio_20_f;
   wire [0:0] 				    h2c_gpio_6_gpio_19_f;
   wire [0:0] 				    h2c_gpio_6_gpio_18_f;
   wire [0:0] 				    h2c_gpio_6_gpio_17_f;
   wire [0:0] 				    h2c_gpio_6_gpio_16_f;
   wire [0:0] 				    h2c_gpio_6_gpio_15_f;
   wire [0:0] 				    h2c_gpio_6_gpio_14_f;
   wire [0:0] 				    h2c_gpio_6_gpio_13_f;
   wire [0:0] 				    h2c_gpio_6_gpio_12_f;
   wire [0:0] 				    h2c_gpio_6_gpio_11_f;
   wire [0:0] 				    h2c_gpio_6_gpio_10_f;
   wire [0:0] 				    h2c_gpio_6_gpio_9_f;
   wire [0:0] 				    h2c_gpio_6_gpio_8_f;
   wire [0:0] 				    h2c_gpio_6_gpio_7_f;
   wire [0:0] 				    h2c_gpio_6_gpio_6_f;
   wire [0:0] 				    h2c_gpio_6_gpio_5_f;
   wire [0:0] 				    h2c_gpio_6_gpio_4_f;
   wire [0:0] 				    h2c_gpio_6_gpio_3_f;
   wire [0:0] 				    h2c_gpio_6_gpio_2_f;
   wire [0:0] 				    h2c_gpio_6_gpio_1_f;
   wire [0:0] 				    h2c_gpio_6_gpio_0_f;
   wire [0:0] 				    h2c_gpio_7_gpio_31_f;
   wire [0:0] 				    h2c_gpio_7_gpio_30_f;
   wire [0:0] 				    h2c_gpio_7_gpio_29_f;
   wire [0:0] 				    h2c_gpio_7_gpio_28_f;
   wire [0:0] 				    h2c_gpio_7_gpio_27_f;
   wire [0:0] 				    h2c_gpio_7_gpio_26_f;
   wire [0:0] 				    h2c_gpio_7_gpio_25_f;
   wire [0:0] 				    h2c_gpio_7_gpio_24_f;
   wire [0:0] 				    h2c_gpio_7_gpio_23_f;
   wire [0:0] 				    h2c_gpio_7_gpio_22_f;
   wire [0:0] 				    h2c_gpio_7_gpio_21_f;
   wire [0:0] 				    h2c_gpio_7_gpio_20_f;
   wire [0:0] 				    h2c_gpio_7_gpio_19_f;
   wire [0:0] 				    h2c_gpio_7_gpio_18_f;
   wire [0:0] 				    h2c_gpio_7_gpio_17_f;
   wire [0:0] 				    h2c_gpio_7_gpio_16_f;
   wire [0:0] 				    h2c_gpio_7_gpio_15_f;
   wire [0:0] 				    h2c_gpio_7_gpio_14_f;
   wire [0:0] 				    h2c_gpio_7_gpio_13_f;
   wire [0:0] 				    h2c_gpio_7_gpio_12_f;
   wire [0:0] 				    h2c_gpio_7_gpio_11_f;
   wire [0:0] 				    h2c_gpio_7_gpio_10_f;
   wire [0:0] 				    h2c_gpio_7_gpio_9_f;
   wire [0:0] 				    h2c_gpio_7_gpio_8_f;
   wire [0:0] 				    h2c_gpio_7_gpio_7_f;
   wire [0:0] 				    h2c_gpio_7_gpio_6_f;
   wire [0:0] 				    h2c_gpio_7_gpio_5_f;
   wire [0:0] 				    h2c_gpio_7_gpio_4_f;
   wire [0:0] 				    h2c_gpio_7_gpio_3_f;
   wire [0:0] 				    h2c_gpio_7_gpio_2_f;
   wire [0:0] 				    h2c_gpio_7_gpio_1_f;
   wire [0:0] 				    h2c_gpio_7_gpio_0_f;
   wire [0:0] 				    h2c_gpio_8_gpio_31_f;
   wire [0:0] 				    h2c_gpio_8_gpio_30_f;
   wire [0:0] 				    h2c_gpio_8_gpio_29_f;
   wire [0:0] 				    h2c_gpio_8_gpio_28_f;
   wire [0:0] 				    h2c_gpio_8_gpio_27_f;
   wire [0:0] 				    h2c_gpio_8_gpio_26_f;
   wire [0:0] 				    h2c_gpio_8_gpio_25_f;
   wire [0:0] 				    h2c_gpio_8_gpio_24_f;
   wire [0:0] 				    h2c_gpio_8_gpio_23_f;
   wire [0:0] 				    h2c_gpio_8_gpio_22_f;
   wire [0:0] 				    h2c_gpio_8_gpio_21_f;
   wire [0:0] 				    h2c_gpio_8_gpio_20_f;
   wire [0:0] 				    h2c_gpio_8_gpio_19_f;
   wire [0:0] 				    h2c_gpio_8_gpio_18_f;
   wire [0:0] 				    h2c_gpio_8_gpio_17_f;
   wire [0:0] 				    h2c_gpio_8_gpio_16_f;
   wire [0:0] 				    h2c_gpio_8_gpio_15_f;
   wire [0:0] 				    h2c_gpio_8_gpio_14_f;
   wire [0:0] 				    h2c_gpio_8_gpio_13_f;
   wire [0:0] 				    h2c_gpio_8_gpio_12_f;
   wire [0:0] 				    h2c_gpio_8_gpio_11_f;
   wire [0:0] 				    h2c_gpio_8_gpio_10_f;
   wire [0:0] 				    h2c_gpio_8_gpio_9_f;
   wire [0:0] 				    h2c_gpio_8_gpio_8_f;
   wire [0:0] 				    h2c_gpio_8_gpio_7_f;
   wire [0:0] 				    h2c_gpio_8_gpio_6_f;
   wire [0:0] 				    h2c_gpio_8_gpio_5_f;
   wire [0:0] 				    h2c_gpio_8_gpio_4_f;
   wire [0:0] 				    h2c_gpio_8_gpio_3_f;
   wire [0:0] 				    h2c_gpio_8_gpio_2_f;
   wire [0:0] 				    h2c_gpio_8_gpio_1_f;
   wire [0:0] 				    h2c_gpio_8_gpio_0_f;
   wire [0:0] 				    h2c_gpio_9_gpio_31_f;
   wire [0:0] 				    h2c_gpio_9_gpio_30_f;
   wire [0:0] 				    h2c_gpio_9_gpio_29_f;
   wire [0:0] 				    h2c_gpio_9_gpio_28_f;
   wire [0:0] 				    h2c_gpio_9_gpio_27_f;
   wire [0:0] 				    h2c_gpio_9_gpio_26_f;
   wire [0:0] 				    h2c_gpio_9_gpio_25_f;
   wire [0:0] 				    h2c_gpio_9_gpio_24_f;
   wire [0:0] 				    h2c_gpio_9_gpio_23_f;
   wire [0:0] 				    h2c_gpio_9_gpio_22_f;
   wire [0:0] 				    h2c_gpio_9_gpio_21_f;
   wire [0:0] 				    h2c_gpio_9_gpio_20_f;
   wire [0:0] 				    h2c_gpio_9_gpio_19_f;
   wire [0:0] 				    h2c_gpio_9_gpio_18_f;
   wire [0:0] 				    h2c_gpio_9_gpio_17_f;
   wire [0:0] 				    h2c_gpio_9_gpio_16_f;
   wire [0:0] 				    h2c_gpio_9_gpio_15_f;
   wire [0:0] 				    h2c_gpio_9_gpio_14_f;
   wire [0:0] 				    h2c_gpio_9_gpio_13_f;
   wire [0:0] 				    h2c_gpio_9_gpio_12_f;
   wire [0:0] 				    h2c_gpio_9_gpio_11_f;
   wire [0:0] 				    h2c_gpio_9_gpio_10_f;
   wire [0:0] 				    h2c_gpio_9_gpio_9_f;
   wire [0:0] 				    h2c_gpio_9_gpio_8_f;
   wire [0:0] 				    h2c_gpio_9_gpio_7_f;
   wire [0:0] 				    h2c_gpio_9_gpio_6_f;
   wire [0:0] 				    h2c_gpio_9_gpio_5_f;
   wire [0:0] 				    h2c_gpio_9_gpio_4_f;
   wire [0:0] 				    h2c_gpio_9_gpio_3_f;
   wire [0:0] 				    h2c_gpio_9_gpio_2_f;
   wire [0:0] 				    h2c_gpio_9_gpio_1_f;
   wire [0:0] 				    h2c_gpio_9_gpio_0_f;
   wire [0:0] 				    h2c_gpio_10_gpio_31_f;
   wire [0:0] 				    h2c_gpio_10_gpio_30_f;
   wire [0:0] 				    h2c_gpio_10_gpio_29_f;
   wire [0:0] 				    h2c_gpio_10_gpio_28_f;
   wire [0:0] 				    h2c_gpio_10_gpio_27_f;
   wire [0:0] 				    h2c_gpio_10_gpio_26_f;
   wire [0:0] 				    h2c_gpio_10_gpio_25_f;
   wire [0:0] 				    h2c_gpio_10_gpio_24_f;
   wire [0:0] 				    h2c_gpio_10_gpio_23_f;
   wire [0:0] 				    h2c_gpio_10_gpio_22_f;
   wire [0:0] 				    h2c_gpio_10_gpio_21_f;
   wire [0:0] 				    h2c_gpio_10_gpio_20_f;
   wire [0:0] 				    h2c_gpio_10_gpio_19_f;
   wire [0:0] 				    h2c_gpio_10_gpio_18_f;
   wire [0:0] 				    h2c_gpio_10_gpio_17_f;
   wire [0:0] 				    h2c_gpio_10_gpio_16_f;
   wire [0:0] 				    h2c_gpio_10_gpio_15_f;
   wire [0:0] 				    h2c_gpio_10_gpio_14_f;
   wire [0:0] 				    h2c_gpio_10_gpio_13_f;
   wire [0:0] 				    h2c_gpio_10_gpio_12_f;
   wire [0:0] 				    h2c_gpio_10_gpio_11_f;
   wire [0:0] 				    h2c_gpio_10_gpio_10_f;
   wire [0:0] 				    h2c_gpio_10_gpio_9_f;
   wire [0:0] 				    h2c_gpio_10_gpio_8_f;
   wire [0:0] 				    h2c_gpio_10_gpio_7_f;
   wire [0:0] 				    h2c_gpio_10_gpio_6_f;
   wire [0:0] 				    h2c_gpio_10_gpio_5_f;
   wire [0:0] 				    h2c_gpio_10_gpio_4_f;
   wire [0:0] 				    h2c_gpio_10_gpio_3_f;
   wire [0:0] 				    h2c_gpio_10_gpio_2_f;
   wire [0:0] 				    h2c_gpio_10_gpio_1_f;
   wire [0:0] 				    h2c_gpio_10_gpio_0_f;
   wire [0:0] 				    h2c_gpio_11_gpio_31_f;
   wire [0:0] 				    h2c_gpio_11_gpio_30_f;
   wire [0:0] 				    h2c_gpio_11_gpio_29_f;
   wire [0:0] 				    h2c_gpio_11_gpio_28_f;
   wire [0:0] 				    h2c_gpio_11_gpio_27_f;
   wire [0:0] 				    h2c_gpio_11_gpio_26_f;
   wire [0:0] 				    h2c_gpio_11_gpio_25_f;
   wire [0:0] 				    h2c_gpio_11_gpio_24_f;
   wire [0:0] 				    h2c_gpio_11_gpio_23_f;
   wire [0:0] 				    h2c_gpio_11_gpio_22_f;
   wire [0:0] 				    h2c_gpio_11_gpio_21_f;
   wire [0:0] 				    h2c_gpio_11_gpio_20_f;
   wire [0:0] 				    h2c_gpio_11_gpio_19_f;
   wire [0:0] 				    h2c_gpio_11_gpio_18_f;
   wire [0:0] 				    h2c_gpio_11_gpio_17_f;
   wire [0:0] 				    h2c_gpio_11_gpio_16_f;
   wire [0:0] 				    h2c_gpio_11_gpio_15_f;
   wire [0:0] 				    h2c_gpio_11_gpio_14_f;
   wire [0:0] 				    h2c_gpio_11_gpio_13_f;
   wire [0:0] 				    h2c_gpio_11_gpio_12_f;
   wire [0:0] 				    h2c_gpio_11_gpio_11_f;
   wire [0:0] 				    h2c_gpio_11_gpio_10_f;
   wire [0:0] 				    h2c_gpio_11_gpio_9_f;
   wire [0:0] 				    h2c_gpio_11_gpio_8_f;
   wire [0:0] 				    h2c_gpio_11_gpio_7_f;
   wire [0:0] 				    h2c_gpio_11_gpio_6_f;
   wire [0:0] 				    h2c_gpio_11_gpio_5_f;
   wire [0:0] 				    h2c_gpio_11_gpio_4_f;
   wire [0:0] 				    h2c_gpio_11_gpio_3_f;
   wire [0:0] 				    h2c_gpio_11_gpio_2_f;
   wire [0:0] 				    h2c_gpio_11_gpio_1_f;
   wire [0:0] 				    h2c_gpio_11_gpio_0_f;
   wire [0:0] 				    h2c_gpio_12_gpio_31_f;
   wire [0:0] 				    h2c_gpio_12_gpio_30_f;
   wire [0:0] 				    h2c_gpio_12_gpio_29_f;
   wire [0:0] 				    h2c_gpio_12_gpio_28_f;
   wire [0:0] 				    h2c_gpio_12_gpio_27_f;
   wire [0:0] 				    h2c_gpio_12_gpio_26_f;
   wire [0:0] 				    h2c_gpio_12_gpio_25_f;
   wire [0:0] 				    h2c_gpio_12_gpio_24_f;
   wire [0:0] 				    h2c_gpio_12_gpio_23_f;
   wire [0:0] 				    h2c_gpio_12_gpio_22_f;
   wire [0:0] 				    h2c_gpio_12_gpio_21_f;
   wire [0:0] 				    h2c_gpio_12_gpio_20_f;
   wire [0:0] 				    h2c_gpio_12_gpio_19_f;
   wire [0:0] 				    h2c_gpio_12_gpio_18_f;
   wire [0:0] 				    h2c_gpio_12_gpio_17_f;
   wire [0:0] 				    h2c_gpio_12_gpio_16_f;
   wire [0:0] 				    h2c_gpio_12_gpio_15_f;
   wire [0:0] 				    h2c_gpio_12_gpio_14_f;
   wire [0:0] 				    h2c_gpio_12_gpio_13_f;
   wire [0:0] 				    h2c_gpio_12_gpio_12_f;
   wire [0:0] 				    h2c_gpio_12_gpio_11_f;
   wire [0:0] 				    h2c_gpio_12_gpio_10_f;
   wire [0:0] 				    h2c_gpio_12_gpio_9_f;
   wire [0:0] 				    h2c_gpio_12_gpio_8_f;
   wire [0:0] 				    h2c_gpio_12_gpio_7_f;
   wire [0:0] 				    h2c_gpio_12_gpio_6_f;
   wire [0:0] 				    h2c_gpio_12_gpio_5_f;
   wire [0:0] 				    h2c_gpio_12_gpio_4_f;
   wire [0:0] 				    h2c_gpio_12_gpio_3_f;
   wire [0:0] 				    h2c_gpio_12_gpio_2_f;
   wire [0:0] 				    h2c_gpio_12_gpio_1_f;
   wire [0:0] 				    h2c_gpio_12_gpio_0_f;
   wire [0:0] 				    h2c_gpio_13_gpio_31_f;
   wire [0:0] 				    h2c_gpio_13_gpio_30_f;
   wire [0:0] 				    h2c_gpio_13_gpio_29_f;
   wire [0:0] 				    h2c_gpio_13_gpio_28_f;
   wire [0:0] 				    h2c_gpio_13_gpio_27_f;
   wire [0:0] 				    h2c_gpio_13_gpio_26_f;
   wire [0:0] 				    h2c_gpio_13_gpio_25_f;
   wire [0:0] 				    h2c_gpio_13_gpio_24_f;
   wire [0:0] 				    h2c_gpio_13_gpio_23_f;
   wire [0:0] 				    h2c_gpio_13_gpio_22_f;
   wire [0:0] 				    h2c_gpio_13_gpio_21_f;
   wire [0:0] 				    h2c_gpio_13_gpio_20_f;
   wire [0:0] 				    h2c_gpio_13_gpio_19_f;
   wire [0:0] 				    h2c_gpio_13_gpio_18_f;
   wire [0:0] 				    h2c_gpio_13_gpio_17_f;
   wire [0:0] 				    h2c_gpio_13_gpio_16_f;
   wire [0:0] 				    h2c_gpio_13_gpio_15_f;
   wire [0:0] 				    h2c_gpio_13_gpio_14_f;
   wire [0:0] 				    h2c_gpio_13_gpio_13_f;
   wire [0:0] 				    h2c_gpio_13_gpio_12_f;
   wire [0:0] 				    h2c_gpio_13_gpio_11_f;
   wire [0:0] 				    h2c_gpio_13_gpio_10_f;
   wire [0:0] 				    h2c_gpio_13_gpio_9_f;
   wire [0:0] 				    h2c_gpio_13_gpio_8_f;
   wire [0:0] 				    h2c_gpio_13_gpio_7_f;
   wire [0:0] 				    h2c_gpio_13_gpio_6_f;
   wire [0:0] 				    h2c_gpio_13_gpio_5_f;
   wire [0:0] 				    h2c_gpio_13_gpio_4_f;
   wire [0:0] 				    h2c_gpio_13_gpio_3_f;
   wire [0:0] 				    h2c_gpio_13_gpio_2_f;
   wire [0:0] 				    h2c_gpio_13_gpio_1_f;
   wire [0:0] 				    h2c_gpio_13_gpio_0_f;
   wire [0:0] 				    h2c_gpio_14_gpio_31_f;
   wire [0:0] 				    h2c_gpio_14_gpio_30_f;
   wire [0:0] 				    h2c_gpio_14_gpio_29_f;
   wire [0:0] 				    h2c_gpio_14_gpio_28_f;
   wire [0:0] 				    h2c_gpio_14_gpio_27_f;
   wire [0:0] 				    h2c_gpio_14_gpio_26_f;
   wire [0:0] 				    h2c_gpio_14_gpio_25_f;
   wire [0:0] 				    h2c_gpio_14_gpio_24_f;
   wire [0:0] 				    h2c_gpio_14_gpio_23_f;
   wire [0:0] 				    h2c_gpio_14_gpio_22_f;
   wire [0:0] 				    h2c_gpio_14_gpio_21_f;
   wire [0:0] 				    h2c_gpio_14_gpio_20_f;
   wire [0:0] 				    h2c_gpio_14_gpio_19_f;
   wire [0:0] 				    h2c_gpio_14_gpio_18_f;
   wire [0:0] 				    h2c_gpio_14_gpio_17_f;
   wire [0:0] 				    h2c_gpio_14_gpio_16_f;
   wire [0:0] 				    h2c_gpio_14_gpio_15_f;
   wire [0:0] 				    h2c_gpio_14_gpio_14_f;
   wire [0:0] 				    h2c_gpio_14_gpio_13_f;
   wire [0:0] 				    h2c_gpio_14_gpio_12_f;
   wire [0:0] 				    h2c_gpio_14_gpio_11_f;
   wire [0:0] 				    h2c_gpio_14_gpio_10_f;
   wire [0:0] 				    h2c_gpio_14_gpio_9_f;
   wire [0:0] 				    h2c_gpio_14_gpio_8_f;
   wire [0:0] 				    h2c_gpio_14_gpio_7_f;
   wire [0:0] 				    h2c_gpio_14_gpio_6_f;
   wire [0:0] 				    h2c_gpio_14_gpio_5_f;
   wire [0:0] 				    h2c_gpio_14_gpio_4_f;
   wire [0:0] 				    h2c_gpio_14_gpio_3_f;
   wire [0:0] 				    h2c_gpio_14_gpio_2_f;
   wire [0:0] 				    h2c_gpio_14_gpio_1_f;
   wire [0:0] 				    h2c_gpio_14_gpio_0_f;
   wire [0:0] 				    h2c_gpio_15_gpio_31_f;
   wire [0:0] 				    h2c_gpio_15_gpio_30_f;
   wire [0:0] 				    h2c_gpio_15_gpio_29_f;
   wire [0:0] 				    h2c_gpio_15_gpio_28_f;
   wire [0:0] 				    h2c_gpio_15_gpio_27_f;
   wire [0:0] 				    h2c_gpio_15_gpio_26_f;
   wire [0:0] 				    h2c_gpio_15_gpio_25_f;
   wire [0:0] 				    h2c_gpio_15_gpio_24_f;
   wire [0:0] 				    h2c_gpio_15_gpio_23_f;
   wire [0:0] 				    h2c_gpio_15_gpio_22_f;
   wire [0:0] 				    h2c_gpio_15_gpio_21_f;
   wire [0:0] 				    h2c_gpio_15_gpio_20_f;
   wire [0:0] 				    h2c_gpio_15_gpio_19_f;
   wire [0:0] 				    h2c_gpio_15_gpio_18_f;
   wire [0:0] 				    h2c_gpio_15_gpio_17_f;
   wire [0:0] 				    h2c_gpio_15_gpio_16_f;
   wire [0:0] 				    h2c_gpio_15_gpio_15_f;
   wire [0:0] 				    h2c_gpio_15_gpio_14_f;
   wire [0:0] 				    h2c_gpio_15_gpio_13_f;
   wire [0:0] 				    h2c_gpio_15_gpio_12_f;
   wire [0:0] 				    h2c_gpio_15_gpio_11_f;
   wire [0:0] 				    h2c_gpio_15_gpio_10_f;
   wire [0:0] 				    h2c_gpio_15_gpio_9_f;
   wire [0:0] 				    h2c_gpio_15_gpio_8_f;
   wire [0:0] 				    h2c_gpio_15_gpio_7_f;
   wire [0:0] 				    h2c_gpio_15_gpio_6_f;
   wire [0:0] 				    h2c_gpio_15_gpio_5_f;
   wire [0:0] 				    h2c_gpio_15_gpio_4_f;
   wire [0:0] 				    h2c_gpio_15_gpio_3_f;
   wire [0:0] 				    h2c_gpio_15_gpio_2_f;
   wire [0:0] 				    h2c_gpio_15_gpio_1_f;
   wire [0:0] 				    h2c_gpio_15_gpio_0_f;
   wire [31:0] 				    rd_req_desc_0_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_0_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_0_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_0_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_0_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_0_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_0_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_0_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_0_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_0_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_0_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_0_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_0_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_0_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_0_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_0_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_0_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_0_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_0_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_0_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_0_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_0_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_0_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_0_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_0_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_0_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_0_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_0_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_0_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_0_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_0_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_0_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_0_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_0_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_0_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_0_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_0_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_0_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_0_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_0_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_0_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_0_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_0_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_0_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_0_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_0_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_0_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_0_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_0_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_0_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_0_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_0_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_0_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_0_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_0_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_0_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_0_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_0_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_0_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_0_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_0_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_0_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_0_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_0_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_0_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_0_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_0_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_0_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_0_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_0_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_0_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_0_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_0_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_0_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_0_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_0_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_0_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_0_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_0_resp_resp_f;
   wire [31:0] 				    rd_req_desc_1_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_1_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_1_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_1_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_1_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_1_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_1_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_1_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_1_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_1_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_1_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_1_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_1_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_1_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_1_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_1_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_1_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_1_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_1_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_1_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_1_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_1_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_1_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_1_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_1_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_1_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_1_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_1_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_1_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_1_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_1_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_1_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_1_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_1_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_1_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_1_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_1_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_1_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_1_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_1_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_1_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_1_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_1_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_1_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_1_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_1_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_1_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_1_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_1_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_1_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_1_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_1_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_1_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_1_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_1_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_1_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_1_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_1_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_1_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_1_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_1_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_1_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_1_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_1_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_1_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_1_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_1_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_1_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_1_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_1_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_1_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_1_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_1_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_1_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_1_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_1_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_1_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_1_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_1_resp_resp_f;
   wire [31:0] 				    rd_req_desc_2_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_2_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_2_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_2_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_2_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_2_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_2_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_2_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_2_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_2_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_2_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_2_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_2_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_2_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_2_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_2_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_2_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_2_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_2_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_2_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_2_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_2_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_2_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_2_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_2_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_2_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_2_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_2_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_2_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_2_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_2_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_2_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_2_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_2_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_2_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_2_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_2_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_2_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_2_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_2_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_2_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_2_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_2_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_2_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_2_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_2_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_2_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_2_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_2_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_2_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_2_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_2_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_2_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_2_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_2_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_2_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_2_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_2_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_2_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_2_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_2_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_2_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_2_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_2_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_2_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_2_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_2_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_2_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_2_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_2_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_2_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_2_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_2_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_2_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_2_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_2_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_2_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_2_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_2_resp_resp_f;
   wire [31:0] 				    rd_req_desc_3_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_3_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_3_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_3_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_3_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_3_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_3_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_3_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_3_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_3_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_3_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_3_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_3_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_3_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_3_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_3_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_3_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_3_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_3_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_3_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_3_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_3_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_3_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_3_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_3_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_3_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_3_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_3_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_3_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_3_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_3_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_3_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_3_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_3_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_3_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_3_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_3_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_3_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_3_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_3_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_3_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_3_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_3_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_3_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_3_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_3_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_3_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_3_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_3_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_3_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_3_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_3_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_3_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_3_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_3_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_3_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_3_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_3_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_3_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_3_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_3_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_3_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_3_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_3_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_3_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_3_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_3_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_3_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_3_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_3_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_3_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_3_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_3_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_3_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_3_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_3_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_3_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_3_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_3_resp_resp_f;
   wire [31:0] 				    rd_req_desc_4_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_4_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_4_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_4_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_4_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_4_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_4_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_4_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_4_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_4_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_4_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_4_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_4_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_4_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_4_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_4_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_4_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_4_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_4_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_4_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_4_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_4_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_4_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_4_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_4_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_4_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_4_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_4_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_4_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_4_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_4_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_4_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_4_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_4_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_4_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_4_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_4_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_4_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_4_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_4_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_4_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_4_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_4_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_4_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_4_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_4_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_4_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_4_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_4_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_4_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_4_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_4_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_4_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_4_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_4_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_4_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_4_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_4_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_4_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_4_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_4_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_4_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_4_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_4_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_4_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_4_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_4_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_4_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_4_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_4_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_4_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_4_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_4_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_4_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_4_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_4_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_4_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_4_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_4_resp_resp_f;
   wire [31:0] 				    rd_req_desc_5_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_5_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_5_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_5_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_5_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_5_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_5_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_5_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_5_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_5_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_5_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_5_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_5_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_5_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_5_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_5_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_5_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_5_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_5_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_5_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_5_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_5_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_5_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_5_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_5_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_5_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_5_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_5_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_5_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_5_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_5_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_5_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_5_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_5_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_5_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_5_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_5_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_5_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_5_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_5_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_5_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_5_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_5_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_5_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_5_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_5_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_5_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_5_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_5_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_5_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_5_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_5_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_5_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_5_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_5_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_5_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_5_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_5_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_5_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_5_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_5_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_5_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_5_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_5_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_5_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_5_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_5_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_5_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_5_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_5_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_5_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_5_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_5_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_5_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_5_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_5_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_5_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_5_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_5_resp_resp_f;
   wire [31:0] 				    rd_req_desc_6_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_6_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_6_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_6_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_6_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_6_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_6_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_6_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_6_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_6_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_6_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_6_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_6_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_6_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_6_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_6_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_6_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_6_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_6_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_6_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_6_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_6_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_6_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_6_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_6_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_6_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_6_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_6_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_6_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_6_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_6_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_6_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_6_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_6_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_6_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_6_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_6_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_6_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_6_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_6_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_6_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_6_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_6_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_6_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_6_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_6_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_6_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_6_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_6_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_6_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_6_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_6_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_6_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_6_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_6_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_6_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_6_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_6_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_6_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_6_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_6_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_6_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_6_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_6_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_6_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_6_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_6_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_6_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_6_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_6_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_6_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_6_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_6_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_6_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_6_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_6_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_6_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_6_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_6_resp_resp_f;
   wire [31:0] 				    rd_req_desc_7_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_7_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_7_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_7_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_7_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_7_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_7_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_7_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_7_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_7_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_7_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_7_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_7_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_7_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_7_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_7_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_7_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_7_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_7_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_7_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_7_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_7_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_7_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_7_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_7_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_7_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_7_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_7_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_7_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_7_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_7_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_7_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_7_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_7_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_7_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_7_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_7_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_7_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_7_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_7_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_7_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_7_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_7_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_7_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_7_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_7_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_7_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_7_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_7_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_7_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_7_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_7_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_7_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_7_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_7_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_7_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_7_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_7_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_7_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_7_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_7_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_7_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_7_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_7_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_7_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_7_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_7_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_7_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_7_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_7_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_7_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_7_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_7_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_7_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_7_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_7_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_7_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_7_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_7_resp_resp_f;
   wire [31:0] 				    rd_req_desc_8_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_8_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_8_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_8_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_8_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_8_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_8_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_8_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_8_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_8_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_8_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_8_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_8_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_8_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_8_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_8_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_8_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_8_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_8_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_8_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_8_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_8_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_8_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_8_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_8_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_8_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_8_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_8_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_8_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_8_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_8_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_8_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_8_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_8_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_8_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_8_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_8_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_8_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_8_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_8_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_8_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_8_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_8_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_8_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_8_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_8_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_8_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_8_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_8_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_8_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_8_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_8_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_8_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_8_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_8_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_8_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_8_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_8_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_8_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_8_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_8_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_8_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_8_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_8_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_8_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_8_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_8_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_8_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_8_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_8_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_8_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_8_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_8_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_8_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_8_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_8_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_8_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_8_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_8_resp_resp_f;
   wire [31:0] 				    rd_req_desc_9_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_9_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_9_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_9_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_9_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_9_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_9_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_9_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_9_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_9_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_9_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_9_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_9_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_9_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_9_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_9_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_9_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_9_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_9_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_9_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_9_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_9_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_9_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_9_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_9_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_9_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_9_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_9_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_9_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_9_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_9_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_9_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_9_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_9_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_9_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_9_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_9_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_9_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_9_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_9_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_9_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_9_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_9_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_9_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_9_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_9_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_9_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_9_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_9_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_9_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_9_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_9_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_9_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_9_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_9_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_9_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_9_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_9_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_9_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_9_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_9_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_9_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_9_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_9_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_9_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_9_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_9_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_9_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_9_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_9_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_9_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_9_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_9_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_9_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_9_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_9_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_9_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_9_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_9_resp_resp_f;
   wire [31:0] 				    rd_req_desc_a_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_a_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_a_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_a_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_a_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_a_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_a_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_a_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_a_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_a_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_a_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_a_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_a_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_a_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_a_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_a_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_a_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_a_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_a_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_a_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_a_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_a_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_a_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_a_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_a_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_a_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_a_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_a_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_a_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_a_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_a_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_a_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_a_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_a_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_a_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_a_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_a_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_a_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_a_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_a_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_a_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_a_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_a_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_a_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_a_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_a_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_a_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_a_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_a_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_a_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_a_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_a_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_a_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_a_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_a_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_a_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_a_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_a_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_a_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_a_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_a_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_a_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_a_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_a_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_a_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_a_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_a_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_a_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_a_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_a_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_a_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_a_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_a_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_a_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_a_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_a_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_a_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_a_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_a_resp_resp_f;
   wire [31:0] 				    rd_req_desc_b_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_b_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_b_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_b_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_b_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_b_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_b_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_b_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_b_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_b_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_b_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_b_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_b_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_b_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_b_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_b_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_b_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_b_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_b_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_b_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_b_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_b_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_b_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_b_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_b_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_b_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_b_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_b_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_b_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_b_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_b_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_b_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_b_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_b_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_b_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_b_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_b_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_b_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_b_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_b_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_b_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_b_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_b_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_b_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_b_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_b_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_b_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_b_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_b_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_b_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_b_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_b_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_b_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_b_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_b_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_b_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_b_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_b_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_b_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_b_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_b_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_b_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_b_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_b_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_b_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_b_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_b_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_b_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_b_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_b_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_b_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_b_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_b_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_b_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_b_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_b_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_b_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_b_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_b_resp_resp_f;
   wire [31:0] 				    rd_req_desc_c_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_c_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_c_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_c_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_c_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_c_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_c_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_c_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_c_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_c_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_c_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_c_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_c_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_c_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_c_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_c_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_c_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_c_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_c_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_c_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_c_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_c_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_c_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_c_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_c_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_c_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_c_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_c_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_c_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_c_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_c_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_c_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_c_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_c_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_c_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_c_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_c_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_c_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_c_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_c_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_c_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_c_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_c_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_c_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_c_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_c_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_c_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_c_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_c_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_c_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_c_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_c_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_c_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_c_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_c_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_c_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_c_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_c_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_c_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_c_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_c_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_c_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_c_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_c_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_c_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_c_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_c_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_c_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_c_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_c_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_c_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_c_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_c_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_c_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_c_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_c_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_c_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_c_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_c_resp_resp_f;
   wire [31:0] 				    rd_req_desc_d_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_d_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_d_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_d_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_d_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_d_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_d_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_d_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_d_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_d_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_d_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_d_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_d_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_d_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_d_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_d_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_d_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_d_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_d_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_d_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_d_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_d_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_d_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_d_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_d_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_d_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_d_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_d_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_d_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_d_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_d_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_d_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_d_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_d_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_d_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_d_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_d_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_d_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_d_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_d_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_d_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_d_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_d_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_d_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_d_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_d_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_d_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_d_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_d_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_d_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_d_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_d_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_d_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_d_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_d_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_d_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_d_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_d_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_d_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_d_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_d_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_d_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_d_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_d_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_d_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_d_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_d_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_d_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_d_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_d_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_d_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_d_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_d_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_d_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_d_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_d_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_d_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_d_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_d_resp_resp_f;
   wire [31:0] 				    rd_req_desc_e_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_e_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_e_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_e_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_e_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_e_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_e_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_e_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_e_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_e_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_e_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_e_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_e_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_e_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_e_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_e_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_e_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_e_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_e_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_e_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_e_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_e_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_e_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_e_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_e_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_e_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_e_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_e_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_e_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_e_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_e_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_e_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_e_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_e_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_e_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_e_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_e_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_e_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_e_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_e_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_e_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_e_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_e_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_e_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_e_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_e_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_e_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_e_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_e_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_e_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_e_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_e_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_e_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_e_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_e_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_e_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_e_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_e_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_e_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_e_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_e_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_e_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_e_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_e_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_e_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_e_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_e_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_e_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_e_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_e_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_e_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_e_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_e_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_e_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_e_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_e_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_e_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_e_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_e_resp_resp_f;
   wire [31:0] 				    rd_req_desc_f_size_txn_size_f;
   wire [2:0] 				    rd_req_desc_f_axsize_axsize_f;
   wire [3:0] 				    rd_req_desc_f_attr_axsnoop_f;
   wire [1:0] 				    rd_req_desc_f_attr_axdomain_f;
   wire [1:0] 				    rd_req_desc_f_attr_axbar_f;
   wire [3:0] 				    rd_req_desc_f_attr_axregion_f;
   wire [3:0] 				    rd_req_desc_f_attr_axqos_f;
   wire [2:0] 				    rd_req_desc_f_attr_axprot_f;
   wire [3:0] 				    rd_req_desc_f_attr_axcache_f;
   wire [0:0] 				    rd_req_desc_f_attr_axlock_f;
   wire [1:0] 				    rd_req_desc_f_attr_axburst_f;
   wire [31:0] 				    rd_req_desc_f_axaddr_0_addr_f;
   wire [31:0] 				    rd_req_desc_f_axaddr_1_addr_f;
   wire [31:0] 				    rd_req_desc_f_axaddr_2_addr_f;
   wire [31:0] 				    rd_req_desc_f_axaddr_3_addr_f;
   wire [31:0] 				    rd_req_desc_f_axid_0_axid_f;
   wire [31:0] 				    rd_req_desc_f_axid_1_axid_f;
   wire [31:0] 				    rd_req_desc_f_axid_2_axid_f;
   wire [31:0] 				    rd_req_desc_f_axid_3_axid_f;
   wire [31:0] 				    rd_req_desc_f_axuser_0_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_1_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_2_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_3_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_4_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_5_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_6_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_7_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_8_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_9_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_10_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_11_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_12_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_13_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_14_axuser_f;
   wire [31:0] 				    rd_req_desc_f_axuser_15_axuser_f;
   wire [13:0] 				    rd_resp_desc_f_data_offset_addr_f;
   wire [31:0] 				    rd_resp_desc_f_data_size_size_f;
   wire [31:0] 				    rd_resp_desc_f_data_host_addr_0_addr_f;
   wire [31:0] 				    rd_resp_desc_f_data_host_addr_1_addr_f;
   wire [31:0] 				    rd_resp_desc_f_data_host_addr_2_addr_f;
   wire [31:0] 				    rd_resp_desc_f_data_host_addr_3_addr_f;
   wire [4:0] 				    rd_resp_desc_f_resp_resp_f;
   wire [31:0] 				    rd_resp_desc_f_xid_0_xid_f;
   wire [31:0] 				    rd_resp_desc_f_xid_1_xid_f;
   wire [31:0] 				    rd_resp_desc_f_xid_2_xid_f;
   wire [31:0] 				    rd_resp_desc_f_xid_3_xid_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_0_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_1_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_2_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_3_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_4_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_5_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_6_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_7_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_8_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_9_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_10_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_11_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_12_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_13_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_14_xuser_f;
   wire [31:0] 				    rd_resp_desc_f_xuser_15_xuser_f;
   wire [0:0] 				    wr_req_desc_f_txn_type_wr_strb_f;
   wire [31:0] 				    wr_req_desc_f_size_txn_size_f;
   wire [13:0] 				    wr_req_desc_f_data_offset_addr_f;
   wire [31:0] 				    wr_req_desc_f_data_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_f_data_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_f_data_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_f_data_host_addr_3_addr_f;
   wire [31:0] 				    wr_req_desc_f_wstrb_host_addr_0_addr_f;
   wire [31:0] 				    wr_req_desc_f_wstrb_host_addr_1_addr_f;
   wire [31:0] 				    wr_req_desc_f_wstrb_host_addr_2_addr_f;
   wire [31:0] 				    wr_req_desc_f_wstrb_host_addr_3_addr_f;
   wire [2:0] 				    wr_req_desc_f_axsize_axsize_f;
   wire [3:0] 				    wr_req_desc_f_attr_axsnoop_f;
   wire [1:0] 				    wr_req_desc_f_attr_axdomain_f;
   wire [1:0] 				    wr_req_desc_f_attr_axbar_f;
   wire [0:0] 				    wr_req_desc_f_attr_awunique_f;
   wire [3:0] 				    wr_req_desc_f_attr_axregion_f;
   wire [3:0] 				    wr_req_desc_f_attr_axqos_f;
   wire [2:0] 				    wr_req_desc_f_attr_axprot_f;
   wire [3:0] 				    wr_req_desc_f_attr_axcache_f;
   wire [0:0] 				    wr_req_desc_f_attr_axlock_f;
   wire [1:0] 				    wr_req_desc_f_attr_axburst_f;
   wire [31:0] 				    wr_req_desc_f_axaddr_0_addr_f;
   wire [31:0] 				    wr_req_desc_f_axaddr_1_addr_f;
   wire [31:0] 				    wr_req_desc_f_axaddr_2_addr_f;
   wire [31:0] 				    wr_req_desc_f_axaddr_3_addr_f;
   wire [31:0] 				    wr_req_desc_f_axid_0_axid_f;
   wire [31:0] 				    wr_req_desc_f_axid_1_axid_f;
   wire [31:0] 				    wr_req_desc_f_axid_2_axid_f;
   wire [31:0] 				    wr_req_desc_f_axid_3_axid_f;
   wire [31:0] 				    wr_req_desc_f_axuser_0_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_1_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_2_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_3_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_4_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_5_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_6_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_7_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_8_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_9_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_10_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_11_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_12_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_13_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_14_axuser_f;
   wire [31:0] 				    wr_req_desc_f_axuser_15_axuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_0_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_1_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_2_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_3_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_4_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_5_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_6_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_7_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_8_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_9_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_10_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_11_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_12_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_13_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_14_wuser_f;
   wire [31:0] 				    wr_req_desc_f_wuser_15_wuser_f;
   wire [4:0] 				    wr_resp_desc_f_resp_resp_f;
   wire [31:0] 				    wr_resp_desc_f_xid_0_xid_f;
   wire [31:0] 				    wr_resp_desc_f_xid_1_xid_f;
   wire [31:0] 				    wr_resp_desc_f_xid_2_xid_f;
   wire [31:0] 				    wr_resp_desc_f_xid_3_xid_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_0_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_1_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_2_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_3_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_4_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_5_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_6_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_7_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_8_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_9_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_10_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_11_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_12_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_13_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_14_xuser_f;
   wire [31:0] 				    wr_resp_desc_f_xuser_15_xuser_f;
   wire [3:0] 				    sn_req_desc_f_attr_acsnoop_f;
   wire [2:0] 				    sn_req_desc_f_attr_acprot_f;
   wire [31:0] 				    sn_req_desc_f_acaddr_0_addr_f;
   wire [31:0] 				    sn_req_desc_f_acaddr_1_addr_f;
   wire [31:0] 				    sn_req_desc_f_acaddr_2_addr_f;
   wire [31:0] 				    sn_req_desc_f_acaddr_3_addr_f;
   wire [4:0] 				    sn_resp_desc_f_resp_resp_f;


   //Fields to use in entire slave RTL ( int_<reg>_<field> )

   wire [0:0] 				    int_bridge_identification_last_bridge;
   wire [7:0] 				    int_version_major_ver;
   wire [7:0] 				    int_version_minor_ver;
   wire [7:0] 				    int_bridge_type_type;
   wire [0:0] 				    int_bridge_config_extend_wstrb;
   wire [7:0] 				    int_bridge_config_id_width;
   wire [2:0] 				    int_bridge_config_data_width;
   wire [9:0] 				    int_bridge_rd_user_config_ruser_width;
   wire [9:0] 				    int_bridge_rd_user_config_aruser_width;
   wire [9:0] 				    int_bridge_wr_user_config_buser_width;
   wire [9:0] 				    int_bridge_wr_user_config_wuser_width;
   wire [9:0] 				    int_bridge_wr_user_config_awuser_width;
   wire [7:0] 				    int_rd_max_desc_resp_max_desc;
   wire [7:0] 				    int_rd_max_desc_req_max_desc;
   wire [7:0] 				    int_wr_max_desc_resp_max_desc;
   wire [7:0] 				    int_wr_max_desc_req_max_desc;
   wire [7:0] 				    int_sn_max_desc_data_max_desc;
   wire [7:0] 				    int_sn_max_desc_resp_max_desc;
   wire [7:0] 				    int_sn_max_desc_req_max_desc;
   wire [0:0] 				    int_reset_dut_srst_3;
   wire [0:0] 				    int_reset_dut_srst_2;
   wire [0:0] 				    int_reset_dut_srst_1;
   wire [0:0] 				    int_reset_dut_srst_0;
   wire [0:0] 				    int_reset_srst;
   wire [0:0] 				    int_mode_select_mode_0_1;
   wire [0:0] 				    int_intr_status_sn_data_fifo_nonempty;
   wire [0:0] 				    int_intr_status_sn_resp_fifo_nonempty;
   wire [0:0] 				    int_intr_status_sn_req_comp;
   wire [0:0] 				    int_intr_status_wr_resp_comp;
   wire [0:0] 				    int_intr_status_wr_req_fifo_nonempty;
   wire [0:0] 				    int_intr_status_rd_resp_comp;
   wire [0:0] 				    int_intr_status_rd_req_fifo_nonempty;
   wire [0:0] 				    int_intr_status_c2h;
   wire [0:0] 				    int_intr_status_error;
   wire [0:0] 				    int_intr_error_status_err_1;
   wire [0:0] 				    int_intr_error_status_err_0;
   wire [0:0] 				    int_intr_error_clear_clr_err_2;
   wire [0:0] 				    int_intr_error_clear_clr_err_1;
   wire [0:0] 				    int_intr_error_clear_clr_err_0;
   wire [0:0] 				    int_intr_error_enable_en_err_2;
   wire [0:0] 				    int_intr_error_enable_en_err_1;
   wire [0:0] 				    int_intr_error_enable_en_err_0;
   wire [15:0] 				    int_rd_req_free_desc_desc;
   wire [0:0] 				    int_rd_req_fifo_pop_desc_valid;
   wire [3:0] 				    int_rd_req_fifo_pop_desc_desc_index;
   wire [4:0] 				    int_rd_req_fifo_fill_level_fill;
   wire [0:0] 				    int_rd_resp_fifo_push_desc_valid;
   wire [3:0] 				    int_rd_resp_fifo_push_desc_desc_index;
   wire [4:0] 				    int_rd_resp_fifo_free_level_free;
   wire [15:0] 				    int_rd_resp_intr_comp_status_comp;
   wire [15:0] 				    int_rd_resp_intr_comp_clear_clr_comp;
   wire [15:0] 				    int_rd_resp_intr_comp_enable_en_comp;
   wire [15:0] 				    int_wr_req_free_desc_desc;
   wire [0:0] 				    int_wr_req_fifo_pop_desc_valid;
   wire [3:0] 				    int_wr_req_fifo_pop_desc_desc_index;
   wire [4:0] 				    int_wr_req_fifo_fill_level_fill;
   wire [0:0] 				    int_wr_resp_fifo_push_desc_valid;
   wire [3:0] 				    int_wr_resp_fifo_push_desc_desc_index;
   wire [4:0] 				    int_wr_resp_fifo_free_level_free;
   wire [15:0] 				    int_wr_resp_intr_comp_status_comp;
   wire [15:0] 				    int_wr_resp_intr_comp_clear_clr_comp;
   wire [15:0] 				    int_wr_resp_intr_comp_enable_en_comp;
   wire [0:0] 				    int_sn_req_fifo_push_desc_valid;
   wire [3:0] 				    int_sn_req_fifo_push_desc_desc_index;
   wire [4:0] 				    int_sn_req_fifo_free_level_free;
   wire [15:0] 				    int_sn_req_intr_comp_status_comp;
   wire [15:0] 				    int_sn_req_intr_comp_clear_clr_comp;
   wire [15:0] 				    int_sn_req_intr_comp_enable_en_comp;
   wire [15:0] 				    int_sn_resp_free_desc_desc;
   wire [0:0] 				    int_sn_resp_fifo_pop_desc_valid;
   wire [3:0] 				    int_sn_resp_fifo_pop_desc_desc_index;
   wire [4:0] 				    int_sn_resp_fifo_fill_level_fill;
   wire [15:0] 				    int_sn_data_free_desc_desc;
   wire [0:0] 				    int_sn_data_fifo_pop_desc_valid;
   wire [3:0] 				    int_sn_data_fifo_pop_desc_desc_index;
   wire [4:0] 				    int_sn_data_fifo_fill_level_fill;
   wire [0:0] 				    int_intr_fifo_enable_en_sn_data_fifo_nonempty;
   wire [0:0] 				    int_intr_fifo_enable_en_sn_resp_fifo_nonempty;
   wire [0:0] 				    int_intr_fifo_enable_en_wr_req_fifo_nonempty;
   wire [0:0] 				    int_intr_fifo_enable_en_rd_req_fifo_nonempty;
   wire [0:0] 				    int_h2c_intr_0_h2c_31;
   wire [0:0] 				    int_h2c_intr_0_h2c_30;
   wire [0:0] 				    int_h2c_intr_0_h2c_29;
   wire [0:0] 				    int_h2c_intr_0_h2c_28;
   wire [0:0] 				    int_h2c_intr_0_h2c_27;
   wire [0:0] 				    int_h2c_intr_0_h2c_26;
   wire [0:0] 				    int_h2c_intr_0_h2c_25;
   wire [0:0] 				    int_h2c_intr_0_h2c_24;
   wire [0:0] 				    int_h2c_intr_0_h2c_23;
   wire [0:0] 				    int_h2c_intr_0_h2c_22;
   wire [0:0] 				    int_h2c_intr_0_h2c_21;
   wire [0:0] 				    int_h2c_intr_0_h2c_20;
   wire [0:0] 				    int_h2c_intr_0_h2c_19;
   wire [0:0] 				    int_h2c_intr_0_h2c_18;
   wire [0:0] 				    int_h2c_intr_0_h2c_17;
   wire [0:0] 				    int_h2c_intr_0_h2c_16;
   wire [0:0] 				    int_h2c_intr_0_h2c_15;
   wire [0:0] 				    int_h2c_intr_0_h2c_14;
   wire [0:0] 				    int_h2c_intr_0_h2c_13;
   wire [0:0] 				    int_h2c_intr_0_h2c_12;
   wire [0:0] 				    int_h2c_intr_0_h2c_11;
   wire [0:0] 				    int_h2c_intr_0_h2c_10;
   wire [0:0] 				    int_h2c_intr_0_h2c_9;
   wire [0:0] 				    int_h2c_intr_0_h2c_8;
   wire [0:0] 				    int_h2c_intr_0_h2c_7;
   wire [0:0] 				    int_h2c_intr_0_h2c_6;
   wire [0:0] 				    int_h2c_intr_0_h2c_5;
   wire [0:0] 				    int_h2c_intr_0_h2c_4;
   wire [0:0] 				    int_h2c_intr_0_h2c_3;
   wire [0:0] 				    int_h2c_intr_0_h2c_2;
   wire [0:0] 				    int_h2c_intr_0_h2c_1;
   wire [0:0] 				    int_h2c_intr_0_h2c_0;
   wire [0:0] 				    int_h2c_intr_1_h2c_31;
   wire [0:0] 				    int_h2c_intr_1_h2c_30;
   wire [0:0] 				    int_h2c_intr_1_h2c_29;
   wire [0:0] 				    int_h2c_intr_1_h2c_28;
   wire [0:0] 				    int_h2c_intr_1_h2c_27;
   wire [0:0] 				    int_h2c_intr_1_h2c_26;
   wire [0:0] 				    int_h2c_intr_1_h2c_25;
   wire [0:0] 				    int_h2c_intr_1_h2c_24;
   wire [0:0] 				    int_h2c_intr_1_h2c_23;
   wire [0:0] 				    int_h2c_intr_1_h2c_22;
   wire [0:0] 				    int_h2c_intr_1_h2c_21;
   wire [0:0] 				    int_h2c_intr_1_h2c_20;
   wire [0:0] 				    int_h2c_intr_1_h2c_19;
   wire [0:0] 				    int_h2c_intr_1_h2c_18;
   wire [0:0] 				    int_h2c_intr_1_h2c_17;
   wire [0:0] 				    int_h2c_intr_1_h2c_16;
   wire [0:0] 				    int_h2c_intr_1_h2c_15;
   wire [0:0] 				    int_h2c_intr_1_h2c_14;
   wire [0:0] 				    int_h2c_intr_1_h2c_13;
   wire [0:0] 				    int_h2c_intr_1_h2c_12;
   wire [0:0] 				    int_h2c_intr_1_h2c_11;
   wire [0:0] 				    int_h2c_intr_1_h2c_10;
   wire [0:0] 				    int_h2c_intr_1_h2c_9;
   wire [0:0] 				    int_h2c_intr_1_h2c_8;
   wire [0:0] 				    int_h2c_intr_1_h2c_7;
   wire [0:0] 				    int_h2c_intr_1_h2c_6;
   wire [0:0] 				    int_h2c_intr_1_h2c_5;
   wire [0:0] 				    int_h2c_intr_1_h2c_4;
   wire [0:0] 				    int_h2c_intr_1_h2c_3;
   wire [0:0] 				    int_h2c_intr_1_h2c_2;
   wire [0:0] 				    int_h2c_intr_1_h2c_1;
   wire [0:0] 				    int_h2c_intr_1_h2c_0;
   wire [0:0] 				    int_h2c_intr_2_h2c_31;
   wire [0:0] 				    int_h2c_intr_2_h2c_30;
   wire [0:0] 				    int_h2c_intr_2_h2c_29;
   wire [0:0] 				    int_h2c_intr_2_h2c_28;
   wire [0:0] 				    int_h2c_intr_2_h2c_27;
   wire [0:0] 				    int_h2c_intr_2_h2c_26;
   wire [0:0] 				    int_h2c_intr_2_h2c_25;
   wire [0:0] 				    int_h2c_intr_2_h2c_24;
   wire [0:0] 				    int_h2c_intr_2_h2c_23;
   wire [0:0] 				    int_h2c_intr_2_h2c_22;
   wire [0:0] 				    int_h2c_intr_2_h2c_21;
   wire [0:0] 				    int_h2c_intr_2_h2c_20;
   wire [0:0] 				    int_h2c_intr_2_h2c_19;
   wire [0:0] 				    int_h2c_intr_2_h2c_18;
   wire [0:0] 				    int_h2c_intr_2_h2c_17;
   wire [0:0] 				    int_h2c_intr_2_h2c_16;
   wire [0:0] 				    int_h2c_intr_2_h2c_15;
   wire [0:0] 				    int_h2c_intr_2_h2c_14;
   wire [0:0] 				    int_h2c_intr_2_h2c_13;
   wire [0:0] 				    int_h2c_intr_2_h2c_12;
   wire [0:0] 				    int_h2c_intr_2_h2c_11;
   wire [0:0] 				    int_h2c_intr_2_h2c_10;
   wire [0:0] 				    int_h2c_intr_2_h2c_9;
   wire [0:0] 				    int_h2c_intr_2_h2c_8;
   wire [0:0] 				    int_h2c_intr_2_h2c_7;
   wire [0:0] 				    int_h2c_intr_2_h2c_6;
   wire [0:0] 				    int_h2c_intr_2_h2c_5;
   wire [0:0] 				    int_h2c_intr_2_h2c_4;
   wire [0:0] 				    int_h2c_intr_2_h2c_3;
   wire [0:0] 				    int_h2c_intr_2_h2c_2;
   wire [0:0] 				    int_h2c_intr_2_h2c_1;
   wire [0:0] 				    int_h2c_intr_2_h2c_0;
   wire [0:0] 				    int_h2c_intr_3_h2c_31;
   wire [0:0] 				    int_h2c_intr_3_h2c_30;
   wire [0:0] 				    int_h2c_intr_3_h2c_29;
   wire [0:0] 				    int_h2c_intr_3_h2c_28;
   wire [0:0] 				    int_h2c_intr_3_h2c_27;
   wire [0:0] 				    int_h2c_intr_3_h2c_26;
   wire [0:0] 				    int_h2c_intr_3_h2c_25;
   wire [0:0] 				    int_h2c_intr_3_h2c_24;
   wire [0:0] 				    int_h2c_intr_3_h2c_23;
   wire [0:0] 				    int_h2c_intr_3_h2c_22;
   wire [0:0] 				    int_h2c_intr_3_h2c_21;
   wire [0:0] 				    int_h2c_intr_3_h2c_20;
   wire [0:0] 				    int_h2c_intr_3_h2c_19;
   wire [0:0] 				    int_h2c_intr_3_h2c_18;
   wire [0:0] 				    int_h2c_intr_3_h2c_17;
   wire [0:0] 				    int_h2c_intr_3_h2c_16;
   wire [0:0] 				    int_h2c_intr_3_h2c_15;
   wire [0:0] 				    int_h2c_intr_3_h2c_14;
   wire [0:0] 				    int_h2c_intr_3_h2c_13;
   wire [0:0] 				    int_h2c_intr_3_h2c_12;
   wire [0:0] 				    int_h2c_intr_3_h2c_11;
   wire [0:0] 				    int_h2c_intr_3_h2c_10;
   wire [0:0] 				    int_h2c_intr_3_h2c_9;
   wire [0:0] 				    int_h2c_intr_3_h2c_8;
   wire [0:0] 				    int_h2c_intr_3_h2c_7;
   wire [0:0] 				    int_h2c_intr_3_h2c_6;
   wire [0:0] 				    int_h2c_intr_3_h2c_5;
   wire [0:0] 				    int_h2c_intr_3_h2c_4;
   wire [0:0] 				    int_h2c_intr_3_h2c_3;
   wire [0:0] 				    int_h2c_intr_3_h2c_2;
   wire [0:0] 				    int_h2c_intr_3_h2c_1;
   wire [0:0] 				    int_h2c_intr_3_h2c_0;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_31;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_30;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_29;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_28;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_27;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_26;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_25;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_24;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_23;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_22;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_21;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_20;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_19;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_18;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_17;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_16;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_15;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_14;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_13;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_12;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_11;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_10;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_9;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_8;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_7;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_6;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_5;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_4;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_3;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_2;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_1;
   wire [0:0] 				    int_c2h_intr_status_0_c2h_0;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_31;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_30;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_29;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_28;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_27;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_26;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_25;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_24;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_23;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_22;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_21;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_20;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_19;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_18;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_17;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_16;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_15;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_14;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_13;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_12;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_11;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_10;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_9;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_8;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_7;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_6;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_5;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_4;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_3;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_2;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_1;
   wire [0:0] 				    int_intr_c2h_toggle_status_0_t_c2h_0;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_31;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_30;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_29;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_28;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_27;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_26;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_25;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_24;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_23;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_22;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_21;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_20;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_19;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_18;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_17;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_16;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_15;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_14;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_13;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_12;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_11;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_10;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_9;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_8;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_7;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_6;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_5;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_4;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_3;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_2;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_1;
   wire [0:0] 				    int_intr_c2h_toggle_clear_0_clr_t_c2h_0;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_31;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_30;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_29;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_28;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_27;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_26;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_25;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_24;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_23;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_22;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_21;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_20;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_19;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_18;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_17;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_16;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_15;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_14;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_13;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_12;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_11;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_10;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_9;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_8;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_7;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_6;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_5;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_4;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_3;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_2;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_1;
   wire [0:0] 				    int_intr_c2h_toggle_enable_0_en_t_c2h_0;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_31;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_30;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_29;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_28;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_27;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_26;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_25;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_24;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_23;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_22;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_21;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_20;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_19;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_18;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_17;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_16;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_15;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_14;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_13;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_12;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_11;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_10;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_9;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_8;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_7;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_6;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_5;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_4;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_3;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_2;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_1;
   wire [0:0] 				    int_c2h_intr_status_1_c2h_0;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_31;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_30;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_29;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_28;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_27;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_26;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_25;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_24;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_23;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_22;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_21;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_20;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_19;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_18;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_17;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_16;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_15;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_14;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_13;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_12;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_11;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_10;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_9;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_8;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_7;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_6;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_5;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_4;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_3;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_2;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_1;
   wire [0:0] 				    int_intr_c2h_toggle_status_1_t_c2h_0;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_31;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_30;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_29;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_28;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_27;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_26;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_25;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_24;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_23;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_22;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_21;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_20;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_19;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_18;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_17;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_16;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_15;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_14;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_13;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_12;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_11;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_10;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_9;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_8;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_7;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_6;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_5;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_4;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_3;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_2;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_1;
   wire [0:0] 				    int_intr_c2h_toggle_clear_1_clr_t_c2h_0;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_31;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_30;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_29;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_28;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_27;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_26;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_25;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_24;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_23;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_22;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_21;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_20;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_19;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_18;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_17;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_16;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_15;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_14;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_13;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_12;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_11;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_10;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_9;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_8;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_7;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_6;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_5;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_4;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_3;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_2;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_1;
   wire [0:0] 				    int_intr_c2h_toggle_enable_1_en_t_c2h_0;
   wire [0:0] 				    int_c2h_gpio_0_gpio_31;
   wire [0:0] 				    int_c2h_gpio_0_gpio_30;
   wire [0:0] 				    int_c2h_gpio_0_gpio_29;
   wire [0:0] 				    int_c2h_gpio_0_gpio_28;
   wire [0:0] 				    int_c2h_gpio_0_gpio_27;
   wire [0:0] 				    int_c2h_gpio_0_gpio_26;
   wire [0:0] 				    int_c2h_gpio_0_gpio_25;
   wire [0:0] 				    int_c2h_gpio_0_gpio_24;
   wire [0:0] 				    int_c2h_gpio_0_gpio_23;
   wire [0:0] 				    int_c2h_gpio_0_gpio_22;
   wire [0:0] 				    int_c2h_gpio_0_gpio_21;
   wire [0:0] 				    int_c2h_gpio_0_gpio_20;
   wire [0:0] 				    int_c2h_gpio_0_gpio_19;
   wire [0:0] 				    int_c2h_gpio_0_gpio_18;
   wire [0:0] 				    int_c2h_gpio_0_gpio_17;
   wire [0:0] 				    int_c2h_gpio_0_gpio_16;
   wire [0:0] 				    int_c2h_gpio_0_gpio_15;
   wire [0:0] 				    int_c2h_gpio_0_gpio_14;
   wire [0:0] 				    int_c2h_gpio_0_gpio_13;
   wire [0:0] 				    int_c2h_gpio_0_gpio_12;
   wire [0:0] 				    int_c2h_gpio_0_gpio_11;
   wire [0:0] 				    int_c2h_gpio_0_gpio_10;
   wire [0:0] 				    int_c2h_gpio_0_gpio_9;
   wire [0:0] 				    int_c2h_gpio_0_gpio_8;
   wire [0:0] 				    int_c2h_gpio_0_gpio_7;
   wire [0:0] 				    int_c2h_gpio_0_gpio_6;
   wire [0:0] 				    int_c2h_gpio_0_gpio_5;
   wire [0:0] 				    int_c2h_gpio_0_gpio_4;
   wire [0:0] 				    int_c2h_gpio_0_gpio_3;
   wire [0:0] 				    int_c2h_gpio_0_gpio_2;
   wire [0:0] 				    int_c2h_gpio_0_gpio_1;
   wire [0:0] 				    int_c2h_gpio_0_gpio_0;
   wire [0:0] 				    int_c2h_gpio_1_gpio_31;
   wire [0:0] 				    int_c2h_gpio_1_gpio_30;
   wire [0:0] 				    int_c2h_gpio_1_gpio_29;
   wire [0:0] 				    int_c2h_gpio_1_gpio_28;
   wire [0:0] 				    int_c2h_gpio_1_gpio_27;
   wire [0:0] 				    int_c2h_gpio_1_gpio_26;
   wire [0:0] 				    int_c2h_gpio_1_gpio_25;
   wire [0:0] 				    int_c2h_gpio_1_gpio_24;
   wire [0:0] 				    int_c2h_gpio_1_gpio_23;
   wire [0:0] 				    int_c2h_gpio_1_gpio_22;
   wire [0:0] 				    int_c2h_gpio_1_gpio_21;
   wire [0:0] 				    int_c2h_gpio_1_gpio_20;
   wire [0:0] 				    int_c2h_gpio_1_gpio_19;
   wire [0:0] 				    int_c2h_gpio_1_gpio_18;
   wire [0:0] 				    int_c2h_gpio_1_gpio_17;
   wire [0:0] 				    int_c2h_gpio_1_gpio_16;
   wire [0:0] 				    int_c2h_gpio_1_gpio_15;
   wire [0:0] 				    int_c2h_gpio_1_gpio_14;
   wire [0:0] 				    int_c2h_gpio_1_gpio_13;
   wire [0:0] 				    int_c2h_gpio_1_gpio_12;
   wire [0:0] 				    int_c2h_gpio_1_gpio_11;
   wire [0:0] 				    int_c2h_gpio_1_gpio_10;
   wire [0:0] 				    int_c2h_gpio_1_gpio_9;
   wire [0:0] 				    int_c2h_gpio_1_gpio_8;
   wire [0:0] 				    int_c2h_gpio_1_gpio_7;
   wire [0:0] 				    int_c2h_gpio_1_gpio_6;
   wire [0:0] 				    int_c2h_gpio_1_gpio_5;
   wire [0:0] 				    int_c2h_gpio_1_gpio_4;
   wire [0:0] 				    int_c2h_gpio_1_gpio_3;
   wire [0:0] 				    int_c2h_gpio_1_gpio_2;
   wire [0:0] 				    int_c2h_gpio_1_gpio_1;
   wire [0:0] 				    int_c2h_gpio_1_gpio_0;
   wire [0:0] 				    int_c2h_gpio_2_gpio_31;
   wire [0:0] 				    int_c2h_gpio_2_gpio_30;
   wire [0:0] 				    int_c2h_gpio_2_gpio_29;
   wire [0:0] 				    int_c2h_gpio_2_gpio_28;
   wire [0:0] 				    int_c2h_gpio_2_gpio_27;
   wire [0:0] 				    int_c2h_gpio_2_gpio_26;
   wire [0:0] 				    int_c2h_gpio_2_gpio_25;
   wire [0:0] 				    int_c2h_gpio_2_gpio_24;
   wire [0:0] 				    int_c2h_gpio_2_gpio_23;
   wire [0:0] 				    int_c2h_gpio_2_gpio_22;
   wire [0:0] 				    int_c2h_gpio_2_gpio_21;
   wire [0:0] 				    int_c2h_gpio_2_gpio_20;
   wire [0:0] 				    int_c2h_gpio_2_gpio_19;
   wire [0:0] 				    int_c2h_gpio_2_gpio_18;
   wire [0:0] 				    int_c2h_gpio_2_gpio_17;
   wire [0:0] 				    int_c2h_gpio_2_gpio_16;
   wire [0:0] 				    int_c2h_gpio_2_gpio_15;
   wire [0:0] 				    int_c2h_gpio_2_gpio_14;
   wire [0:0] 				    int_c2h_gpio_2_gpio_13;
   wire [0:0] 				    int_c2h_gpio_2_gpio_12;
   wire [0:0] 				    int_c2h_gpio_2_gpio_11;
   wire [0:0] 				    int_c2h_gpio_2_gpio_10;
   wire [0:0] 				    int_c2h_gpio_2_gpio_9;
   wire [0:0] 				    int_c2h_gpio_2_gpio_8;
   wire [0:0] 				    int_c2h_gpio_2_gpio_7;
   wire [0:0] 				    int_c2h_gpio_2_gpio_6;
   wire [0:0] 				    int_c2h_gpio_2_gpio_5;
   wire [0:0] 				    int_c2h_gpio_2_gpio_4;
   wire [0:0] 				    int_c2h_gpio_2_gpio_3;
   wire [0:0] 				    int_c2h_gpio_2_gpio_2;
   wire [0:0] 				    int_c2h_gpio_2_gpio_1;
   wire [0:0] 				    int_c2h_gpio_2_gpio_0;
   wire [0:0] 				    int_c2h_gpio_3_gpio_31;
   wire [0:0] 				    int_c2h_gpio_3_gpio_30;
   wire [0:0] 				    int_c2h_gpio_3_gpio_29;
   wire [0:0] 				    int_c2h_gpio_3_gpio_28;
   wire [0:0] 				    int_c2h_gpio_3_gpio_27;
   wire [0:0] 				    int_c2h_gpio_3_gpio_26;
   wire [0:0] 				    int_c2h_gpio_3_gpio_25;
   wire [0:0] 				    int_c2h_gpio_3_gpio_24;
   wire [0:0] 				    int_c2h_gpio_3_gpio_23;
   wire [0:0] 				    int_c2h_gpio_3_gpio_22;
   wire [0:0] 				    int_c2h_gpio_3_gpio_21;
   wire [0:0] 				    int_c2h_gpio_3_gpio_20;
   wire [0:0] 				    int_c2h_gpio_3_gpio_19;
   wire [0:0] 				    int_c2h_gpio_3_gpio_18;
   wire [0:0] 				    int_c2h_gpio_3_gpio_17;
   wire [0:0] 				    int_c2h_gpio_3_gpio_16;
   wire [0:0] 				    int_c2h_gpio_3_gpio_15;
   wire [0:0] 				    int_c2h_gpio_3_gpio_14;
   wire [0:0] 				    int_c2h_gpio_3_gpio_13;
   wire [0:0] 				    int_c2h_gpio_3_gpio_12;
   wire [0:0] 				    int_c2h_gpio_3_gpio_11;
   wire [0:0] 				    int_c2h_gpio_3_gpio_10;
   wire [0:0] 				    int_c2h_gpio_3_gpio_9;
   wire [0:0] 				    int_c2h_gpio_3_gpio_8;
   wire [0:0] 				    int_c2h_gpio_3_gpio_7;
   wire [0:0] 				    int_c2h_gpio_3_gpio_6;
   wire [0:0] 				    int_c2h_gpio_3_gpio_5;
   wire [0:0] 				    int_c2h_gpio_3_gpio_4;
   wire [0:0] 				    int_c2h_gpio_3_gpio_3;
   wire [0:0] 				    int_c2h_gpio_3_gpio_2;
   wire [0:0] 				    int_c2h_gpio_3_gpio_1;
   wire [0:0] 				    int_c2h_gpio_3_gpio_0;
   wire [0:0] 				    int_c2h_gpio_4_gpio_31;
   wire [0:0] 				    int_c2h_gpio_4_gpio_30;
   wire [0:0] 				    int_c2h_gpio_4_gpio_29;
   wire [0:0] 				    int_c2h_gpio_4_gpio_28;
   wire [0:0] 				    int_c2h_gpio_4_gpio_27;
   wire [0:0] 				    int_c2h_gpio_4_gpio_26;
   wire [0:0] 				    int_c2h_gpio_4_gpio_25;
   wire [0:0] 				    int_c2h_gpio_4_gpio_24;
   wire [0:0] 				    int_c2h_gpio_4_gpio_23;
   wire [0:0] 				    int_c2h_gpio_4_gpio_22;
   wire [0:0] 				    int_c2h_gpio_4_gpio_21;
   wire [0:0] 				    int_c2h_gpio_4_gpio_20;
   wire [0:0] 				    int_c2h_gpio_4_gpio_19;
   wire [0:0] 				    int_c2h_gpio_4_gpio_18;
   wire [0:0] 				    int_c2h_gpio_4_gpio_17;
   wire [0:0] 				    int_c2h_gpio_4_gpio_16;
   wire [0:0] 				    int_c2h_gpio_4_gpio_15;
   wire [0:0] 				    int_c2h_gpio_4_gpio_14;
   wire [0:0] 				    int_c2h_gpio_4_gpio_13;
   wire [0:0] 				    int_c2h_gpio_4_gpio_12;
   wire [0:0] 				    int_c2h_gpio_4_gpio_11;
   wire [0:0] 				    int_c2h_gpio_4_gpio_10;
   wire [0:0] 				    int_c2h_gpio_4_gpio_9;
   wire [0:0] 				    int_c2h_gpio_4_gpio_8;
   wire [0:0] 				    int_c2h_gpio_4_gpio_7;
   wire [0:0] 				    int_c2h_gpio_4_gpio_6;
   wire [0:0] 				    int_c2h_gpio_4_gpio_5;
   wire [0:0] 				    int_c2h_gpio_4_gpio_4;
   wire [0:0] 				    int_c2h_gpio_4_gpio_3;
   wire [0:0] 				    int_c2h_gpio_4_gpio_2;
   wire [0:0] 				    int_c2h_gpio_4_gpio_1;
   wire [0:0] 				    int_c2h_gpio_4_gpio_0;
   wire [0:0] 				    int_c2h_gpio_5_gpio_31;
   wire [0:0] 				    int_c2h_gpio_5_gpio_30;
   wire [0:0] 				    int_c2h_gpio_5_gpio_29;
   wire [0:0] 				    int_c2h_gpio_5_gpio_28;
   wire [0:0] 				    int_c2h_gpio_5_gpio_27;
   wire [0:0] 				    int_c2h_gpio_5_gpio_26;
   wire [0:0] 				    int_c2h_gpio_5_gpio_25;
   wire [0:0] 				    int_c2h_gpio_5_gpio_24;
   wire [0:0] 				    int_c2h_gpio_5_gpio_23;
   wire [0:0] 				    int_c2h_gpio_5_gpio_22;
   wire [0:0] 				    int_c2h_gpio_5_gpio_21;
   wire [0:0] 				    int_c2h_gpio_5_gpio_20;
   wire [0:0] 				    int_c2h_gpio_5_gpio_19;
   wire [0:0] 				    int_c2h_gpio_5_gpio_18;
   wire [0:0] 				    int_c2h_gpio_5_gpio_17;
   wire [0:0] 				    int_c2h_gpio_5_gpio_16;
   wire [0:0] 				    int_c2h_gpio_5_gpio_15;
   wire [0:0] 				    int_c2h_gpio_5_gpio_14;
   wire [0:0] 				    int_c2h_gpio_5_gpio_13;
   wire [0:0] 				    int_c2h_gpio_5_gpio_12;
   wire [0:0] 				    int_c2h_gpio_5_gpio_11;
   wire [0:0] 				    int_c2h_gpio_5_gpio_10;
   wire [0:0] 				    int_c2h_gpio_5_gpio_9;
   wire [0:0] 				    int_c2h_gpio_5_gpio_8;
   wire [0:0] 				    int_c2h_gpio_5_gpio_7;
   wire [0:0] 				    int_c2h_gpio_5_gpio_6;
   wire [0:0] 				    int_c2h_gpio_5_gpio_5;
   wire [0:0] 				    int_c2h_gpio_5_gpio_4;
   wire [0:0] 				    int_c2h_gpio_5_gpio_3;
   wire [0:0] 				    int_c2h_gpio_5_gpio_2;
   wire [0:0] 				    int_c2h_gpio_5_gpio_1;
   wire [0:0] 				    int_c2h_gpio_5_gpio_0;
   wire [0:0] 				    int_c2h_gpio_6_gpio_31;
   wire [0:0] 				    int_c2h_gpio_6_gpio_30;
   wire [0:0] 				    int_c2h_gpio_6_gpio_29;
   wire [0:0] 				    int_c2h_gpio_6_gpio_28;
   wire [0:0] 				    int_c2h_gpio_6_gpio_27;
   wire [0:0] 				    int_c2h_gpio_6_gpio_26;
   wire [0:0] 				    int_c2h_gpio_6_gpio_25;
   wire [0:0] 				    int_c2h_gpio_6_gpio_24;
   wire [0:0] 				    int_c2h_gpio_6_gpio_23;
   wire [0:0] 				    int_c2h_gpio_6_gpio_22;
   wire [0:0] 				    int_c2h_gpio_6_gpio_21;
   wire [0:0] 				    int_c2h_gpio_6_gpio_20;
   wire [0:0] 				    int_c2h_gpio_6_gpio_19;
   wire [0:0] 				    int_c2h_gpio_6_gpio_18;
   wire [0:0] 				    int_c2h_gpio_6_gpio_17;
   wire [0:0] 				    int_c2h_gpio_6_gpio_16;
   wire [0:0] 				    int_c2h_gpio_6_gpio_15;
   wire [0:0] 				    int_c2h_gpio_6_gpio_14;
   wire [0:0] 				    int_c2h_gpio_6_gpio_13;
   wire [0:0] 				    int_c2h_gpio_6_gpio_12;
   wire [0:0] 				    int_c2h_gpio_6_gpio_11;
   wire [0:0] 				    int_c2h_gpio_6_gpio_10;
   wire [0:0] 				    int_c2h_gpio_6_gpio_9;
   wire [0:0] 				    int_c2h_gpio_6_gpio_8;
   wire [0:0] 				    int_c2h_gpio_6_gpio_7;
   wire [0:0] 				    int_c2h_gpio_6_gpio_6;
   wire [0:0] 				    int_c2h_gpio_6_gpio_5;
   wire [0:0] 				    int_c2h_gpio_6_gpio_4;
   wire [0:0] 				    int_c2h_gpio_6_gpio_3;
   wire [0:0] 				    int_c2h_gpio_6_gpio_2;
   wire [0:0] 				    int_c2h_gpio_6_gpio_1;
   wire [0:0] 				    int_c2h_gpio_6_gpio_0;
   wire [0:0] 				    int_c2h_gpio_7_gpio_31;
   wire [0:0] 				    int_c2h_gpio_7_gpio_30;
   wire [0:0] 				    int_c2h_gpio_7_gpio_29;
   wire [0:0] 				    int_c2h_gpio_7_gpio_28;
   wire [0:0] 				    int_c2h_gpio_7_gpio_27;
   wire [0:0] 				    int_c2h_gpio_7_gpio_26;
   wire [0:0] 				    int_c2h_gpio_7_gpio_25;
   wire [0:0] 				    int_c2h_gpio_7_gpio_24;
   wire [0:0] 				    int_c2h_gpio_7_gpio_23;
   wire [0:0] 				    int_c2h_gpio_7_gpio_22;
   wire [0:0] 				    int_c2h_gpio_7_gpio_21;
   wire [0:0] 				    int_c2h_gpio_7_gpio_20;
   wire [0:0] 				    int_c2h_gpio_7_gpio_19;
   wire [0:0] 				    int_c2h_gpio_7_gpio_18;
   wire [0:0] 				    int_c2h_gpio_7_gpio_17;
   wire [0:0] 				    int_c2h_gpio_7_gpio_16;
   wire [0:0] 				    int_c2h_gpio_7_gpio_15;
   wire [0:0] 				    int_c2h_gpio_7_gpio_14;
   wire [0:0] 				    int_c2h_gpio_7_gpio_13;
   wire [0:0] 				    int_c2h_gpio_7_gpio_12;
   wire [0:0] 				    int_c2h_gpio_7_gpio_11;
   wire [0:0] 				    int_c2h_gpio_7_gpio_10;
   wire [0:0] 				    int_c2h_gpio_7_gpio_9;
   wire [0:0] 				    int_c2h_gpio_7_gpio_8;
   wire [0:0] 				    int_c2h_gpio_7_gpio_7;
   wire [0:0] 				    int_c2h_gpio_7_gpio_6;
   wire [0:0] 				    int_c2h_gpio_7_gpio_5;
   wire [0:0] 				    int_c2h_gpio_7_gpio_4;
   wire [0:0] 				    int_c2h_gpio_7_gpio_3;
   wire [0:0] 				    int_c2h_gpio_7_gpio_2;
   wire [0:0] 				    int_c2h_gpio_7_gpio_1;
   wire [0:0] 				    int_c2h_gpio_7_gpio_0;
   wire [0:0] 				    int_c2h_gpio_8_gpio_31;
   wire [0:0] 				    int_c2h_gpio_8_gpio_30;
   wire [0:0] 				    int_c2h_gpio_8_gpio_29;
   wire [0:0] 				    int_c2h_gpio_8_gpio_28;
   wire [0:0] 				    int_c2h_gpio_8_gpio_27;
   wire [0:0] 				    int_c2h_gpio_8_gpio_26;
   wire [0:0] 				    int_c2h_gpio_8_gpio_25;
   wire [0:0] 				    int_c2h_gpio_8_gpio_24;
   wire [0:0] 				    int_c2h_gpio_8_gpio_23;
   wire [0:0] 				    int_c2h_gpio_8_gpio_22;
   wire [0:0] 				    int_c2h_gpio_8_gpio_21;
   wire [0:0] 				    int_c2h_gpio_8_gpio_20;
   wire [0:0] 				    int_c2h_gpio_8_gpio_19;
   wire [0:0] 				    int_c2h_gpio_8_gpio_18;
   wire [0:0] 				    int_c2h_gpio_8_gpio_17;
   wire [0:0] 				    int_c2h_gpio_8_gpio_16;
   wire [0:0] 				    int_c2h_gpio_8_gpio_15;
   wire [0:0] 				    int_c2h_gpio_8_gpio_14;
   wire [0:0] 				    int_c2h_gpio_8_gpio_13;
   wire [0:0] 				    int_c2h_gpio_8_gpio_12;
   wire [0:0] 				    int_c2h_gpio_8_gpio_11;
   wire [0:0] 				    int_c2h_gpio_8_gpio_10;
   wire [0:0] 				    int_c2h_gpio_8_gpio_9;
   wire [0:0] 				    int_c2h_gpio_8_gpio_8;
   wire [0:0] 				    int_c2h_gpio_8_gpio_7;
   wire [0:0] 				    int_c2h_gpio_8_gpio_6;
   wire [0:0] 				    int_c2h_gpio_8_gpio_5;
   wire [0:0] 				    int_c2h_gpio_8_gpio_4;
   wire [0:0] 				    int_c2h_gpio_8_gpio_3;
   wire [0:0] 				    int_c2h_gpio_8_gpio_2;
   wire [0:0] 				    int_c2h_gpio_8_gpio_1;
   wire [0:0] 				    int_c2h_gpio_8_gpio_0;
   wire [0:0] 				    int_c2h_gpio_9_gpio_31;
   wire [0:0] 				    int_c2h_gpio_9_gpio_30;
   wire [0:0] 				    int_c2h_gpio_9_gpio_29;
   wire [0:0] 				    int_c2h_gpio_9_gpio_28;
   wire [0:0] 				    int_c2h_gpio_9_gpio_27;
   wire [0:0] 				    int_c2h_gpio_9_gpio_26;
   wire [0:0] 				    int_c2h_gpio_9_gpio_25;
   wire [0:0] 				    int_c2h_gpio_9_gpio_24;
   wire [0:0] 				    int_c2h_gpio_9_gpio_23;
   wire [0:0] 				    int_c2h_gpio_9_gpio_22;
   wire [0:0] 				    int_c2h_gpio_9_gpio_21;
   wire [0:0] 				    int_c2h_gpio_9_gpio_20;
   wire [0:0] 				    int_c2h_gpio_9_gpio_19;
   wire [0:0] 				    int_c2h_gpio_9_gpio_18;
   wire [0:0] 				    int_c2h_gpio_9_gpio_17;
   wire [0:0] 				    int_c2h_gpio_9_gpio_16;
   wire [0:0] 				    int_c2h_gpio_9_gpio_15;
   wire [0:0] 				    int_c2h_gpio_9_gpio_14;
   wire [0:0] 				    int_c2h_gpio_9_gpio_13;
   wire [0:0] 				    int_c2h_gpio_9_gpio_12;
   wire [0:0] 				    int_c2h_gpio_9_gpio_11;
   wire [0:0] 				    int_c2h_gpio_9_gpio_10;
   wire [0:0] 				    int_c2h_gpio_9_gpio_9;
   wire [0:0] 				    int_c2h_gpio_9_gpio_8;
   wire [0:0] 				    int_c2h_gpio_9_gpio_7;
   wire [0:0] 				    int_c2h_gpio_9_gpio_6;
   wire [0:0] 				    int_c2h_gpio_9_gpio_5;
   wire [0:0] 				    int_c2h_gpio_9_gpio_4;
   wire [0:0] 				    int_c2h_gpio_9_gpio_3;
   wire [0:0] 				    int_c2h_gpio_9_gpio_2;
   wire [0:0] 				    int_c2h_gpio_9_gpio_1;
   wire [0:0] 				    int_c2h_gpio_9_gpio_0;
   wire [0:0] 				    int_c2h_gpio_10_gpio_31;
   wire [0:0] 				    int_c2h_gpio_10_gpio_30;
   wire [0:0] 				    int_c2h_gpio_10_gpio_29;
   wire [0:0] 				    int_c2h_gpio_10_gpio_28;
   wire [0:0] 				    int_c2h_gpio_10_gpio_27;
   wire [0:0] 				    int_c2h_gpio_10_gpio_26;
   wire [0:0] 				    int_c2h_gpio_10_gpio_25;
   wire [0:0] 				    int_c2h_gpio_10_gpio_24;
   wire [0:0] 				    int_c2h_gpio_10_gpio_23;
   wire [0:0] 				    int_c2h_gpio_10_gpio_22;
   wire [0:0] 				    int_c2h_gpio_10_gpio_21;
   wire [0:0] 				    int_c2h_gpio_10_gpio_20;
   wire [0:0] 				    int_c2h_gpio_10_gpio_19;
   wire [0:0] 				    int_c2h_gpio_10_gpio_18;
   wire [0:0] 				    int_c2h_gpio_10_gpio_17;
   wire [0:0] 				    int_c2h_gpio_10_gpio_16;
   wire [0:0] 				    int_c2h_gpio_10_gpio_15;
   wire [0:0] 				    int_c2h_gpio_10_gpio_14;
   wire [0:0] 				    int_c2h_gpio_10_gpio_13;
   wire [0:0] 				    int_c2h_gpio_10_gpio_12;
   wire [0:0] 				    int_c2h_gpio_10_gpio_11;
   wire [0:0] 				    int_c2h_gpio_10_gpio_10;
   wire [0:0] 				    int_c2h_gpio_10_gpio_9;
   wire [0:0] 				    int_c2h_gpio_10_gpio_8;
   wire [0:0] 				    int_c2h_gpio_10_gpio_7;
   wire [0:0] 				    int_c2h_gpio_10_gpio_6;
   wire [0:0] 				    int_c2h_gpio_10_gpio_5;
   wire [0:0] 				    int_c2h_gpio_10_gpio_4;
   wire [0:0] 				    int_c2h_gpio_10_gpio_3;
   wire [0:0] 				    int_c2h_gpio_10_gpio_2;
   wire [0:0] 				    int_c2h_gpio_10_gpio_1;
   wire [0:0] 				    int_c2h_gpio_10_gpio_0;
   wire [0:0] 				    int_c2h_gpio_11_gpio_31;
   wire [0:0] 				    int_c2h_gpio_11_gpio_30;
   wire [0:0] 				    int_c2h_gpio_11_gpio_29;
   wire [0:0] 				    int_c2h_gpio_11_gpio_28;
   wire [0:0] 				    int_c2h_gpio_11_gpio_27;
   wire [0:0] 				    int_c2h_gpio_11_gpio_26;
   wire [0:0] 				    int_c2h_gpio_11_gpio_25;
   wire [0:0] 				    int_c2h_gpio_11_gpio_24;
   wire [0:0] 				    int_c2h_gpio_11_gpio_23;
   wire [0:0] 				    int_c2h_gpio_11_gpio_22;
   wire [0:0] 				    int_c2h_gpio_11_gpio_21;
   wire [0:0] 				    int_c2h_gpio_11_gpio_20;
   wire [0:0] 				    int_c2h_gpio_11_gpio_19;
   wire [0:0] 				    int_c2h_gpio_11_gpio_18;
   wire [0:0] 				    int_c2h_gpio_11_gpio_17;
   wire [0:0] 				    int_c2h_gpio_11_gpio_16;
   wire [0:0] 				    int_c2h_gpio_11_gpio_15;
   wire [0:0] 				    int_c2h_gpio_11_gpio_14;
   wire [0:0] 				    int_c2h_gpio_11_gpio_13;
   wire [0:0] 				    int_c2h_gpio_11_gpio_12;
   wire [0:0] 				    int_c2h_gpio_11_gpio_11;
   wire [0:0] 				    int_c2h_gpio_11_gpio_10;
   wire [0:0] 				    int_c2h_gpio_11_gpio_9;
   wire [0:0] 				    int_c2h_gpio_11_gpio_8;
   wire [0:0] 				    int_c2h_gpio_11_gpio_7;
   wire [0:0] 				    int_c2h_gpio_11_gpio_6;
   wire [0:0] 				    int_c2h_gpio_11_gpio_5;
   wire [0:0] 				    int_c2h_gpio_11_gpio_4;
   wire [0:0] 				    int_c2h_gpio_11_gpio_3;
   wire [0:0] 				    int_c2h_gpio_11_gpio_2;
   wire [0:0] 				    int_c2h_gpio_11_gpio_1;
   wire [0:0] 				    int_c2h_gpio_11_gpio_0;
   wire [0:0] 				    int_c2h_gpio_12_gpio_31;
   wire [0:0] 				    int_c2h_gpio_12_gpio_30;
   wire [0:0] 				    int_c2h_gpio_12_gpio_29;
   wire [0:0] 				    int_c2h_gpio_12_gpio_28;
   wire [0:0] 				    int_c2h_gpio_12_gpio_27;
   wire [0:0] 				    int_c2h_gpio_12_gpio_26;
   wire [0:0] 				    int_c2h_gpio_12_gpio_25;
   wire [0:0] 				    int_c2h_gpio_12_gpio_24;
   wire [0:0] 				    int_c2h_gpio_12_gpio_23;
   wire [0:0] 				    int_c2h_gpio_12_gpio_22;
   wire [0:0] 				    int_c2h_gpio_12_gpio_21;
   wire [0:0] 				    int_c2h_gpio_12_gpio_20;
   wire [0:0] 				    int_c2h_gpio_12_gpio_19;
   wire [0:0] 				    int_c2h_gpio_12_gpio_18;
   wire [0:0] 				    int_c2h_gpio_12_gpio_17;
   wire [0:0] 				    int_c2h_gpio_12_gpio_16;
   wire [0:0] 				    int_c2h_gpio_12_gpio_15;
   wire [0:0] 				    int_c2h_gpio_12_gpio_14;
   wire [0:0] 				    int_c2h_gpio_12_gpio_13;
   wire [0:0] 				    int_c2h_gpio_12_gpio_12;
   wire [0:0] 				    int_c2h_gpio_12_gpio_11;
   wire [0:0] 				    int_c2h_gpio_12_gpio_10;
   wire [0:0] 				    int_c2h_gpio_12_gpio_9;
   wire [0:0] 				    int_c2h_gpio_12_gpio_8;
   wire [0:0] 				    int_c2h_gpio_12_gpio_7;
   wire [0:0] 				    int_c2h_gpio_12_gpio_6;
   wire [0:0] 				    int_c2h_gpio_12_gpio_5;
   wire [0:0] 				    int_c2h_gpio_12_gpio_4;
   wire [0:0] 				    int_c2h_gpio_12_gpio_3;
   wire [0:0] 				    int_c2h_gpio_12_gpio_2;
   wire [0:0] 				    int_c2h_gpio_12_gpio_1;
   wire [0:0] 				    int_c2h_gpio_12_gpio_0;
   wire [0:0] 				    int_c2h_gpio_13_gpio_31;
   wire [0:0] 				    int_c2h_gpio_13_gpio_30;
   wire [0:0] 				    int_c2h_gpio_13_gpio_29;
   wire [0:0] 				    int_c2h_gpio_13_gpio_28;
   wire [0:0] 				    int_c2h_gpio_13_gpio_27;
   wire [0:0] 				    int_c2h_gpio_13_gpio_26;
   wire [0:0] 				    int_c2h_gpio_13_gpio_25;
   wire [0:0] 				    int_c2h_gpio_13_gpio_24;
   wire [0:0] 				    int_c2h_gpio_13_gpio_23;
   wire [0:0] 				    int_c2h_gpio_13_gpio_22;
   wire [0:0] 				    int_c2h_gpio_13_gpio_21;
   wire [0:0] 				    int_c2h_gpio_13_gpio_20;
   wire [0:0] 				    int_c2h_gpio_13_gpio_19;
   wire [0:0] 				    int_c2h_gpio_13_gpio_18;
   wire [0:0] 				    int_c2h_gpio_13_gpio_17;
   wire [0:0] 				    int_c2h_gpio_13_gpio_16;
   wire [0:0] 				    int_c2h_gpio_13_gpio_15;
   wire [0:0] 				    int_c2h_gpio_13_gpio_14;
   wire [0:0] 				    int_c2h_gpio_13_gpio_13;
   wire [0:0] 				    int_c2h_gpio_13_gpio_12;
   wire [0:0] 				    int_c2h_gpio_13_gpio_11;
   wire [0:0] 				    int_c2h_gpio_13_gpio_10;
   wire [0:0] 				    int_c2h_gpio_13_gpio_9;
   wire [0:0] 				    int_c2h_gpio_13_gpio_8;
   wire [0:0] 				    int_c2h_gpio_13_gpio_7;
   wire [0:0] 				    int_c2h_gpio_13_gpio_6;
   wire [0:0] 				    int_c2h_gpio_13_gpio_5;
   wire [0:0] 				    int_c2h_gpio_13_gpio_4;
   wire [0:0] 				    int_c2h_gpio_13_gpio_3;
   wire [0:0] 				    int_c2h_gpio_13_gpio_2;
   wire [0:0] 				    int_c2h_gpio_13_gpio_1;
   wire [0:0] 				    int_c2h_gpio_13_gpio_0;
   wire [0:0] 				    int_c2h_gpio_14_gpio_31;
   wire [0:0] 				    int_c2h_gpio_14_gpio_30;
   wire [0:0] 				    int_c2h_gpio_14_gpio_29;
   wire [0:0] 				    int_c2h_gpio_14_gpio_28;
   wire [0:0] 				    int_c2h_gpio_14_gpio_27;
   wire [0:0] 				    int_c2h_gpio_14_gpio_26;
   wire [0:0] 				    int_c2h_gpio_14_gpio_25;
   wire [0:0] 				    int_c2h_gpio_14_gpio_24;
   wire [0:0] 				    int_c2h_gpio_14_gpio_23;
   wire [0:0] 				    int_c2h_gpio_14_gpio_22;
   wire [0:0] 				    int_c2h_gpio_14_gpio_21;
   wire [0:0] 				    int_c2h_gpio_14_gpio_20;
   wire [0:0] 				    int_c2h_gpio_14_gpio_19;
   wire [0:0] 				    int_c2h_gpio_14_gpio_18;
   wire [0:0] 				    int_c2h_gpio_14_gpio_17;
   wire [0:0] 				    int_c2h_gpio_14_gpio_16;
   wire [0:0] 				    int_c2h_gpio_14_gpio_15;
   wire [0:0] 				    int_c2h_gpio_14_gpio_14;
   wire [0:0] 				    int_c2h_gpio_14_gpio_13;
   wire [0:0] 				    int_c2h_gpio_14_gpio_12;
   wire [0:0] 				    int_c2h_gpio_14_gpio_11;
   wire [0:0] 				    int_c2h_gpio_14_gpio_10;
   wire [0:0] 				    int_c2h_gpio_14_gpio_9;
   wire [0:0] 				    int_c2h_gpio_14_gpio_8;
   wire [0:0] 				    int_c2h_gpio_14_gpio_7;
   wire [0:0] 				    int_c2h_gpio_14_gpio_6;
   wire [0:0] 				    int_c2h_gpio_14_gpio_5;
   wire [0:0] 				    int_c2h_gpio_14_gpio_4;
   wire [0:0] 				    int_c2h_gpio_14_gpio_3;
   wire [0:0] 				    int_c2h_gpio_14_gpio_2;
   wire [0:0] 				    int_c2h_gpio_14_gpio_1;
   wire [0:0] 				    int_c2h_gpio_14_gpio_0;
   wire [0:0] 				    int_c2h_gpio_15_gpio_31;
   wire [0:0] 				    int_c2h_gpio_15_gpio_30;
   wire [0:0] 				    int_c2h_gpio_15_gpio_29;
   wire [0:0] 				    int_c2h_gpio_15_gpio_28;
   wire [0:0] 				    int_c2h_gpio_15_gpio_27;
   wire [0:0] 				    int_c2h_gpio_15_gpio_26;
   wire [0:0] 				    int_c2h_gpio_15_gpio_25;
   wire [0:0] 				    int_c2h_gpio_15_gpio_24;
   wire [0:0] 				    int_c2h_gpio_15_gpio_23;
   wire [0:0] 				    int_c2h_gpio_15_gpio_22;
   wire [0:0] 				    int_c2h_gpio_15_gpio_21;
   wire [0:0] 				    int_c2h_gpio_15_gpio_20;
   wire [0:0] 				    int_c2h_gpio_15_gpio_19;
   wire [0:0] 				    int_c2h_gpio_15_gpio_18;
   wire [0:0] 				    int_c2h_gpio_15_gpio_17;
   wire [0:0] 				    int_c2h_gpio_15_gpio_16;
   wire [0:0] 				    int_c2h_gpio_15_gpio_15;
   wire [0:0] 				    int_c2h_gpio_15_gpio_14;
   wire [0:0] 				    int_c2h_gpio_15_gpio_13;
   wire [0:0] 				    int_c2h_gpio_15_gpio_12;
   wire [0:0] 				    int_c2h_gpio_15_gpio_11;
   wire [0:0] 				    int_c2h_gpio_15_gpio_10;
   wire [0:0] 				    int_c2h_gpio_15_gpio_9;
   wire [0:0] 				    int_c2h_gpio_15_gpio_8;
   wire [0:0] 				    int_c2h_gpio_15_gpio_7;
   wire [0:0] 				    int_c2h_gpio_15_gpio_6;
   wire [0:0] 				    int_c2h_gpio_15_gpio_5;
   wire [0:0] 				    int_c2h_gpio_15_gpio_4;
   wire [0:0] 				    int_c2h_gpio_15_gpio_3;
   wire [0:0] 				    int_c2h_gpio_15_gpio_2;
   wire [0:0] 				    int_c2h_gpio_15_gpio_1;
   wire [0:0] 				    int_c2h_gpio_15_gpio_0;
   wire [0:0] 				    int_h2c_gpio_0_gpio_31;
   wire [0:0] 				    int_h2c_gpio_0_gpio_30;
   wire [0:0] 				    int_h2c_gpio_0_gpio_29;
   wire [0:0] 				    int_h2c_gpio_0_gpio_28;
   wire [0:0] 				    int_h2c_gpio_0_gpio_27;
   wire [0:0] 				    int_h2c_gpio_0_gpio_26;
   wire [0:0] 				    int_h2c_gpio_0_gpio_25;
   wire [0:0] 				    int_h2c_gpio_0_gpio_24;
   wire [0:0] 				    int_h2c_gpio_0_gpio_23;
   wire [0:0] 				    int_h2c_gpio_0_gpio_22;
   wire [0:0] 				    int_h2c_gpio_0_gpio_21;
   wire [0:0] 				    int_h2c_gpio_0_gpio_20;
   wire [0:0] 				    int_h2c_gpio_0_gpio_19;
   wire [0:0] 				    int_h2c_gpio_0_gpio_18;
   wire [0:0] 				    int_h2c_gpio_0_gpio_17;
   wire [0:0] 				    int_h2c_gpio_0_gpio_16;
   wire [0:0] 				    int_h2c_gpio_0_gpio_15;
   wire [0:0] 				    int_h2c_gpio_0_gpio_14;
   wire [0:0] 				    int_h2c_gpio_0_gpio_13;
   wire [0:0] 				    int_h2c_gpio_0_gpio_12;
   wire [0:0] 				    int_h2c_gpio_0_gpio_11;
   wire [0:0] 				    int_h2c_gpio_0_gpio_10;
   wire [0:0] 				    int_h2c_gpio_0_gpio_9;
   wire [0:0] 				    int_h2c_gpio_0_gpio_8;
   wire [0:0] 				    int_h2c_gpio_0_gpio_7;
   wire [0:0] 				    int_h2c_gpio_0_gpio_6;
   wire [0:0] 				    int_h2c_gpio_0_gpio_5;
   wire [0:0] 				    int_h2c_gpio_0_gpio_4;
   wire [0:0] 				    int_h2c_gpio_0_gpio_3;
   wire [0:0] 				    int_h2c_gpio_0_gpio_2;
   wire [0:0] 				    int_h2c_gpio_0_gpio_1;
   wire [0:0] 				    int_h2c_gpio_0_gpio_0;
   wire [0:0] 				    int_h2c_gpio_1_gpio_31;
   wire [0:0] 				    int_h2c_gpio_1_gpio_30;
   wire [0:0] 				    int_h2c_gpio_1_gpio_29;
   wire [0:0] 				    int_h2c_gpio_1_gpio_28;
   wire [0:0] 				    int_h2c_gpio_1_gpio_27;
   wire [0:0] 				    int_h2c_gpio_1_gpio_26;
   wire [0:0] 				    int_h2c_gpio_1_gpio_25;
   wire [0:0] 				    int_h2c_gpio_1_gpio_24;
   wire [0:0] 				    int_h2c_gpio_1_gpio_23;
   wire [0:0] 				    int_h2c_gpio_1_gpio_22;
   wire [0:0] 				    int_h2c_gpio_1_gpio_21;
   wire [0:0] 				    int_h2c_gpio_1_gpio_20;
   wire [0:0] 				    int_h2c_gpio_1_gpio_19;
   wire [0:0] 				    int_h2c_gpio_1_gpio_18;
   wire [0:0] 				    int_h2c_gpio_1_gpio_17;
   wire [0:0] 				    int_h2c_gpio_1_gpio_16;
   wire [0:0] 				    int_h2c_gpio_1_gpio_15;
   wire [0:0] 				    int_h2c_gpio_1_gpio_14;
   wire [0:0] 				    int_h2c_gpio_1_gpio_13;
   wire [0:0] 				    int_h2c_gpio_1_gpio_12;
   wire [0:0] 				    int_h2c_gpio_1_gpio_11;
   wire [0:0] 				    int_h2c_gpio_1_gpio_10;
   wire [0:0] 				    int_h2c_gpio_1_gpio_9;
   wire [0:0] 				    int_h2c_gpio_1_gpio_8;
   wire [0:0] 				    int_h2c_gpio_1_gpio_7;
   wire [0:0] 				    int_h2c_gpio_1_gpio_6;
   wire [0:0] 				    int_h2c_gpio_1_gpio_5;
   wire [0:0] 				    int_h2c_gpio_1_gpio_4;
   wire [0:0] 				    int_h2c_gpio_1_gpio_3;
   wire [0:0] 				    int_h2c_gpio_1_gpio_2;
   wire [0:0] 				    int_h2c_gpio_1_gpio_1;
   wire [0:0] 				    int_h2c_gpio_1_gpio_0;
   wire [0:0] 				    int_h2c_gpio_2_gpio_31;
   wire [0:0] 				    int_h2c_gpio_2_gpio_30;
   wire [0:0] 				    int_h2c_gpio_2_gpio_29;
   wire [0:0] 				    int_h2c_gpio_2_gpio_28;
   wire [0:0] 				    int_h2c_gpio_2_gpio_27;
   wire [0:0] 				    int_h2c_gpio_2_gpio_26;
   wire [0:0] 				    int_h2c_gpio_2_gpio_25;
   wire [0:0] 				    int_h2c_gpio_2_gpio_24;
   wire [0:0] 				    int_h2c_gpio_2_gpio_23;
   wire [0:0] 				    int_h2c_gpio_2_gpio_22;
   wire [0:0] 				    int_h2c_gpio_2_gpio_21;
   wire [0:0] 				    int_h2c_gpio_2_gpio_20;
   wire [0:0] 				    int_h2c_gpio_2_gpio_19;
   wire [0:0] 				    int_h2c_gpio_2_gpio_18;
   wire [0:0] 				    int_h2c_gpio_2_gpio_17;
   wire [0:0] 				    int_h2c_gpio_2_gpio_16;
   wire [0:0] 				    int_h2c_gpio_2_gpio_15;
   wire [0:0] 				    int_h2c_gpio_2_gpio_14;
   wire [0:0] 				    int_h2c_gpio_2_gpio_13;
   wire [0:0] 				    int_h2c_gpio_2_gpio_12;
   wire [0:0] 				    int_h2c_gpio_2_gpio_11;
   wire [0:0] 				    int_h2c_gpio_2_gpio_10;
   wire [0:0] 				    int_h2c_gpio_2_gpio_9;
   wire [0:0] 				    int_h2c_gpio_2_gpio_8;
   wire [0:0] 				    int_h2c_gpio_2_gpio_7;
   wire [0:0] 				    int_h2c_gpio_2_gpio_6;
   wire [0:0] 				    int_h2c_gpio_2_gpio_5;
   wire [0:0] 				    int_h2c_gpio_2_gpio_4;
   wire [0:0] 				    int_h2c_gpio_2_gpio_3;
   wire [0:0] 				    int_h2c_gpio_2_gpio_2;
   wire [0:0] 				    int_h2c_gpio_2_gpio_1;
   wire [0:0] 				    int_h2c_gpio_2_gpio_0;
   wire [0:0] 				    int_h2c_gpio_3_gpio_31;
   wire [0:0] 				    int_h2c_gpio_3_gpio_30;
   wire [0:0] 				    int_h2c_gpio_3_gpio_29;
   wire [0:0] 				    int_h2c_gpio_3_gpio_28;
   wire [0:0] 				    int_h2c_gpio_3_gpio_27;
   wire [0:0] 				    int_h2c_gpio_3_gpio_26;
   wire [0:0] 				    int_h2c_gpio_3_gpio_25;
   wire [0:0] 				    int_h2c_gpio_3_gpio_24;
   wire [0:0] 				    int_h2c_gpio_3_gpio_23;
   wire [0:0] 				    int_h2c_gpio_3_gpio_22;
   wire [0:0] 				    int_h2c_gpio_3_gpio_21;
   wire [0:0] 				    int_h2c_gpio_3_gpio_20;
   wire [0:0] 				    int_h2c_gpio_3_gpio_19;
   wire [0:0] 				    int_h2c_gpio_3_gpio_18;
   wire [0:0] 				    int_h2c_gpio_3_gpio_17;
   wire [0:0] 				    int_h2c_gpio_3_gpio_16;
   wire [0:0] 				    int_h2c_gpio_3_gpio_15;
   wire [0:0] 				    int_h2c_gpio_3_gpio_14;
   wire [0:0] 				    int_h2c_gpio_3_gpio_13;
   wire [0:0] 				    int_h2c_gpio_3_gpio_12;
   wire [0:0] 				    int_h2c_gpio_3_gpio_11;
   wire [0:0] 				    int_h2c_gpio_3_gpio_10;
   wire [0:0] 				    int_h2c_gpio_3_gpio_9;
   wire [0:0] 				    int_h2c_gpio_3_gpio_8;
   wire [0:0] 				    int_h2c_gpio_3_gpio_7;
   wire [0:0] 				    int_h2c_gpio_3_gpio_6;
   wire [0:0] 				    int_h2c_gpio_3_gpio_5;
   wire [0:0] 				    int_h2c_gpio_3_gpio_4;
   wire [0:0] 				    int_h2c_gpio_3_gpio_3;
   wire [0:0] 				    int_h2c_gpio_3_gpio_2;
   wire [0:0] 				    int_h2c_gpio_3_gpio_1;
   wire [0:0] 				    int_h2c_gpio_3_gpio_0;
   wire [0:0] 				    int_h2c_gpio_4_gpio_31;
   wire [0:0] 				    int_h2c_gpio_4_gpio_30;
   wire [0:0] 				    int_h2c_gpio_4_gpio_29;
   wire [0:0] 				    int_h2c_gpio_4_gpio_28;
   wire [0:0] 				    int_h2c_gpio_4_gpio_27;
   wire [0:0] 				    int_h2c_gpio_4_gpio_26;
   wire [0:0] 				    int_h2c_gpio_4_gpio_25;
   wire [0:0] 				    int_h2c_gpio_4_gpio_24;
   wire [0:0] 				    int_h2c_gpio_4_gpio_23;
   wire [0:0] 				    int_h2c_gpio_4_gpio_22;
   wire [0:0] 				    int_h2c_gpio_4_gpio_21;
   wire [0:0] 				    int_h2c_gpio_4_gpio_20;
   wire [0:0] 				    int_h2c_gpio_4_gpio_19;
   wire [0:0] 				    int_h2c_gpio_4_gpio_18;
   wire [0:0] 				    int_h2c_gpio_4_gpio_17;
   wire [0:0] 				    int_h2c_gpio_4_gpio_16;
   wire [0:0] 				    int_h2c_gpio_4_gpio_15;
   wire [0:0] 				    int_h2c_gpio_4_gpio_14;
   wire [0:0] 				    int_h2c_gpio_4_gpio_13;
   wire [0:0] 				    int_h2c_gpio_4_gpio_12;
   wire [0:0] 				    int_h2c_gpio_4_gpio_11;
   wire [0:0] 				    int_h2c_gpio_4_gpio_10;
   wire [0:0] 				    int_h2c_gpio_4_gpio_9;
   wire [0:0] 				    int_h2c_gpio_4_gpio_8;
   wire [0:0] 				    int_h2c_gpio_4_gpio_7;
   wire [0:0] 				    int_h2c_gpio_4_gpio_6;
   wire [0:0] 				    int_h2c_gpio_4_gpio_5;
   wire [0:0] 				    int_h2c_gpio_4_gpio_4;
   wire [0:0] 				    int_h2c_gpio_4_gpio_3;
   wire [0:0] 				    int_h2c_gpio_4_gpio_2;
   wire [0:0] 				    int_h2c_gpio_4_gpio_1;
   wire [0:0] 				    int_h2c_gpio_4_gpio_0;
   wire [0:0] 				    int_h2c_gpio_5_gpio_31;
   wire [0:0] 				    int_h2c_gpio_5_gpio_30;
   wire [0:0] 				    int_h2c_gpio_5_gpio_29;
   wire [0:0] 				    int_h2c_gpio_5_gpio_28;
   wire [0:0] 				    int_h2c_gpio_5_gpio_27;
   wire [0:0] 				    int_h2c_gpio_5_gpio_26;
   wire [0:0] 				    int_h2c_gpio_5_gpio_25;
   wire [0:0] 				    int_h2c_gpio_5_gpio_24;
   wire [0:0] 				    int_h2c_gpio_5_gpio_23;
   wire [0:0] 				    int_h2c_gpio_5_gpio_22;
   wire [0:0] 				    int_h2c_gpio_5_gpio_21;
   wire [0:0] 				    int_h2c_gpio_5_gpio_20;
   wire [0:0] 				    int_h2c_gpio_5_gpio_19;
   wire [0:0] 				    int_h2c_gpio_5_gpio_18;
   wire [0:0] 				    int_h2c_gpio_5_gpio_17;
   wire [0:0] 				    int_h2c_gpio_5_gpio_16;
   wire [0:0] 				    int_h2c_gpio_5_gpio_15;
   wire [0:0] 				    int_h2c_gpio_5_gpio_14;
   wire [0:0] 				    int_h2c_gpio_5_gpio_13;
   wire [0:0] 				    int_h2c_gpio_5_gpio_12;
   wire [0:0] 				    int_h2c_gpio_5_gpio_11;
   wire [0:0] 				    int_h2c_gpio_5_gpio_10;
   wire [0:0] 				    int_h2c_gpio_5_gpio_9;
   wire [0:0] 				    int_h2c_gpio_5_gpio_8;
   wire [0:0] 				    int_h2c_gpio_5_gpio_7;
   wire [0:0] 				    int_h2c_gpio_5_gpio_6;
   wire [0:0] 				    int_h2c_gpio_5_gpio_5;
   wire [0:0] 				    int_h2c_gpio_5_gpio_4;
   wire [0:0] 				    int_h2c_gpio_5_gpio_3;
   wire [0:0] 				    int_h2c_gpio_5_gpio_2;
   wire [0:0] 				    int_h2c_gpio_5_gpio_1;
   wire [0:0] 				    int_h2c_gpio_5_gpio_0;
   wire [0:0] 				    int_h2c_gpio_6_gpio_31;
   wire [0:0] 				    int_h2c_gpio_6_gpio_30;
   wire [0:0] 				    int_h2c_gpio_6_gpio_29;
   wire [0:0] 				    int_h2c_gpio_6_gpio_28;
   wire [0:0] 				    int_h2c_gpio_6_gpio_27;
   wire [0:0] 				    int_h2c_gpio_6_gpio_26;
   wire [0:0] 				    int_h2c_gpio_6_gpio_25;
   wire [0:0] 				    int_h2c_gpio_6_gpio_24;
   wire [0:0] 				    int_h2c_gpio_6_gpio_23;
   wire [0:0] 				    int_h2c_gpio_6_gpio_22;
   wire [0:0] 				    int_h2c_gpio_6_gpio_21;
   wire [0:0] 				    int_h2c_gpio_6_gpio_20;
   wire [0:0] 				    int_h2c_gpio_6_gpio_19;
   wire [0:0] 				    int_h2c_gpio_6_gpio_18;
   wire [0:0] 				    int_h2c_gpio_6_gpio_17;
   wire [0:0] 				    int_h2c_gpio_6_gpio_16;
   wire [0:0] 				    int_h2c_gpio_6_gpio_15;
   wire [0:0] 				    int_h2c_gpio_6_gpio_14;
   wire [0:0] 				    int_h2c_gpio_6_gpio_13;
   wire [0:0] 				    int_h2c_gpio_6_gpio_12;
   wire [0:0] 				    int_h2c_gpio_6_gpio_11;
   wire [0:0] 				    int_h2c_gpio_6_gpio_10;
   wire [0:0] 				    int_h2c_gpio_6_gpio_9;
   wire [0:0] 				    int_h2c_gpio_6_gpio_8;
   wire [0:0] 				    int_h2c_gpio_6_gpio_7;
   wire [0:0] 				    int_h2c_gpio_6_gpio_6;
   wire [0:0] 				    int_h2c_gpio_6_gpio_5;
   wire [0:0] 				    int_h2c_gpio_6_gpio_4;
   wire [0:0] 				    int_h2c_gpio_6_gpio_3;
   wire [0:0] 				    int_h2c_gpio_6_gpio_2;
   wire [0:0] 				    int_h2c_gpio_6_gpio_1;
   wire [0:0] 				    int_h2c_gpio_6_gpio_0;
   wire [0:0] 				    int_h2c_gpio_7_gpio_31;
   wire [0:0] 				    int_h2c_gpio_7_gpio_30;
   wire [0:0] 				    int_h2c_gpio_7_gpio_29;
   wire [0:0] 				    int_h2c_gpio_7_gpio_28;
   wire [0:0] 				    int_h2c_gpio_7_gpio_27;
   wire [0:0] 				    int_h2c_gpio_7_gpio_26;
   wire [0:0] 				    int_h2c_gpio_7_gpio_25;
   wire [0:0] 				    int_h2c_gpio_7_gpio_24;
   wire [0:0] 				    int_h2c_gpio_7_gpio_23;
   wire [0:0] 				    int_h2c_gpio_7_gpio_22;
   wire [0:0] 				    int_h2c_gpio_7_gpio_21;
   wire [0:0] 				    int_h2c_gpio_7_gpio_20;
   wire [0:0] 				    int_h2c_gpio_7_gpio_19;
   wire [0:0] 				    int_h2c_gpio_7_gpio_18;
   wire [0:0] 				    int_h2c_gpio_7_gpio_17;
   wire [0:0] 				    int_h2c_gpio_7_gpio_16;
   wire [0:0] 				    int_h2c_gpio_7_gpio_15;
   wire [0:0] 				    int_h2c_gpio_7_gpio_14;
   wire [0:0] 				    int_h2c_gpio_7_gpio_13;
   wire [0:0] 				    int_h2c_gpio_7_gpio_12;
   wire [0:0] 				    int_h2c_gpio_7_gpio_11;
   wire [0:0] 				    int_h2c_gpio_7_gpio_10;
   wire [0:0] 				    int_h2c_gpio_7_gpio_9;
   wire [0:0] 				    int_h2c_gpio_7_gpio_8;
   wire [0:0] 				    int_h2c_gpio_7_gpio_7;
   wire [0:0] 				    int_h2c_gpio_7_gpio_6;
   wire [0:0] 				    int_h2c_gpio_7_gpio_5;
   wire [0:0] 				    int_h2c_gpio_7_gpio_4;
   wire [0:0] 				    int_h2c_gpio_7_gpio_3;
   wire [0:0] 				    int_h2c_gpio_7_gpio_2;
   wire [0:0] 				    int_h2c_gpio_7_gpio_1;
   wire [0:0] 				    int_h2c_gpio_7_gpio_0;
   wire [0:0] 				    int_h2c_gpio_8_gpio_31;
   wire [0:0] 				    int_h2c_gpio_8_gpio_30;
   wire [0:0] 				    int_h2c_gpio_8_gpio_29;
   wire [0:0] 				    int_h2c_gpio_8_gpio_28;
   wire [0:0] 				    int_h2c_gpio_8_gpio_27;
   wire [0:0] 				    int_h2c_gpio_8_gpio_26;
   wire [0:0] 				    int_h2c_gpio_8_gpio_25;
   wire [0:0] 				    int_h2c_gpio_8_gpio_24;
   wire [0:0] 				    int_h2c_gpio_8_gpio_23;
   wire [0:0] 				    int_h2c_gpio_8_gpio_22;
   wire [0:0] 				    int_h2c_gpio_8_gpio_21;
   wire [0:0] 				    int_h2c_gpio_8_gpio_20;
   wire [0:0] 				    int_h2c_gpio_8_gpio_19;
   wire [0:0] 				    int_h2c_gpio_8_gpio_18;
   wire [0:0] 				    int_h2c_gpio_8_gpio_17;
   wire [0:0] 				    int_h2c_gpio_8_gpio_16;
   wire [0:0] 				    int_h2c_gpio_8_gpio_15;
   wire [0:0] 				    int_h2c_gpio_8_gpio_14;
   wire [0:0] 				    int_h2c_gpio_8_gpio_13;
   wire [0:0] 				    int_h2c_gpio_8_gpio_12;
   wire [0:0] 				    int_h2c_gpio_8_gpio_11;
   wire [0:0] 				    int_h2c_gpio_8_gpio_10;
   wire [0:0] 				    int_h2c_gpio_8_gpio_9;
   wire [0:0] 				    int_h2c_gpio_8_gpio_8;
   wire [0:0] 				    int_h2c_gpio_8_gpio_7;
   wire [0:0] 				    int_h2c_gpio_8_gpio_6;
   wire [0:0] 				    int_h2c_gpio_8_gpio_5;
   wire [0:0] 				    int_h2c_gpio_8_gpio_4;
   wire [0:0] 				    int_h2c_gpio_8_gpio_3;
   wire [0:0] 				    int_h2c_gpio_8_gpio_2;
   wire [0:0] 				    int_h2c_gpio_8_gpio_1;
   wire [0:0] 				    int_h2c_gpio_8_gpio_0;
   wire [0:0] 				    int_h2c_gpio_9_gpio_31;
   wire [0:0] 				    int_h2c_gpio_9_gpio_30;
   wire [0:0] 				    int_h2c_gpio_9_gpio_29;
   wire [0:0] 				    int_h2c_gpio_9_gpio_28;
   wire [0:0] 				    int_h2c_gpio_9_gpio_27;
   wire [0:0] 				    int_h2c_gpio_9_gpio_26;
   wire [0:0] 				    int_h2c_gpio_9_gpio_25;
   wire [0:0] 				    int_h2c_gpio_9_gpio_24;
   wire [0:0] 				    int_h2c_gpio_9_gpio_23;
   wire [0:0] 				    int_h2c_gpio_9_gpio_22;
   wire [0:0] 				    int_h2c_gpio_9_gpio_21;
   wire [0:0] 				    int_h2c_gpio_9_gpio_20;
   wire [0:0] 				    int_h2c_gpio_9_gpio_19;
   wire [0:0] 				    int_h2c_gpio_9_gpio_18;
   wire [0:0] 				    int_h2c_gpio_9_gpio_17;
   wire [0:0] 				    int_h2c_gpio_9_gpio_16;
   wire [0:0] 				    int_h2c_gpio_9_gpio_15;
   wire [0:0] 				    int_h2c_gpio_9_gpio_14;
   wire [0:0] 				    int_h2c_gpio_9_gpio_13;
   wire [0:0] 				    int_h2c_gpio_9_gpio_12;
   wire [0:0] 				    int_h2c_gpio_9_gpio_11;
   wire [0:0] 				    int_h2c_gpio_9_gpio_10;
   wire [0:0] 				    int_h2c_gpio_9_gpio_9;
   wire [0:0] 				    int_h2c_gpio_9_gpio_8;
   wire [0:0] 				    int_h2c_gpio_9_gpio_7;
   wire [0:0] 				    int_h2c_gpio_9_gpio_6;
   wire [0:0] 				    int_h2c_gpio_9_gpio_5;
   wire [0:0] 				    int_h2c_gpio_9_gpio_4;
   wire [0:0] 				    int_h2c_gpio_9_gpio_3;
   wire [0:0] 				    int_h2c_gpio_9_gpio_2;
   wire [0:0] 				    int_h2c_gpio_9_gpio_1;
   wire [0:0] 				    int_h2c_gpio_9_gpio_0;
   wire [0:0] 				    int_h2c_gpio_10_gpio_31;
   wire [0:0] 				    int_h2c_gpio_10_gpio_30;
   wire [0:0] 				    int_h2c_gpio_10_gpio_29;
   wire [0:0] 				    int_h2c_gpio_10_gpio_28;
   wire [0:0] 				    int_h2c_gpio_10_gpio_27;
   wire [0:0] 				    int_h2c_gpio_10_gpio_26;
   wire [0:0] 				    int_h2c_gpio_10_gpio_25;
   wire [0:0] 				    int_h2c_gpio_10_gpio_24;
   wire [0:0] 				    int_h2c_gpio_10_gpio_23;
   wire [0:0] 				    int_h2c_gpio_10_gpio_22;
   wire [0:0] 				    int_h2c_gpio_10_gpio_21;
   wire [0:0] 				    int_h2c_gpio_10_gpio_20;
   wire [0:0] 				    int_h2c_gpio_10_gpio_19;
   wire [0:0] 				    int_h2c_gpio_10_gpio_18;
   wire [0:0] 				    int_h2c_gpio_10_gpio_17;
   wire [0:0] 				    int_h2c_gpio_10_gpio_16;
   wire [0:0] 				    int_h2c_gpio_10_gpio_15;
   wire [0:0] 				    int_h2c_gpio_10_gpio_14;
   wire [0:0] 				    int_h2c_gpio_10_gpio_13;
   wire [0:0] 				    int_h2c_gpio_10_gpio_12;
   wire [0:0] 				    int_h2c_gpio_10_gpio_11;
   wire [0:0] 				    int_h2c_gpio_10_gpio_10;
   wire [0:0] 				    int_h2c_gpio_10_gpio_9;
   wire [0:0] 				    int_h2c_gpio_10_gpio_8;
   wire [0:0] 				    int_h2c_gpio_10_gpio_7;
   wire [0:0] 				    int_h2c_gpio_10_gpio_6;
   wire [0:0] 				    int_h2c_gpio_10_gpio_5;
   wire [0:0] 				    int_h2c_gpio_10_gpio_4;
   wire [0:0] 				    int_h2c_gpio_10_gpio_3;
   wire [0:0] 				    int_h2c_gpio_10_gpio_2;
   wire [0:0] 				    int_h2c_gpio_10_gpio_1;
   wire [0:0] 				    int_h2c_gpio_10_gpio_0;
   wire [0:0] 				    int_h2c_gpio_11_gpio_31;
   wire [0:0] 				    int_h2c_gpio_11_gpio_30;
   wire [0:0] 				    int_h2c_gpio_11_gpio_29;
   wire [0:0] 				    int_h2c_gpio_11_gpio_28;
   wire [0:0] 				    int_h2c_gpio_11_gpio_27;
   wire [0:0] 				    int_h2c_gpio_11_gpio_26;
   wire [0:0] 				    int_h2c_gpio_11_gpio_25;
   wire [0:0] 				    int_h2c_gpio_11_gpio_24;
   wire [0:0] 				    int_h2c_gpio_11_gpio_23;
   wire [0:0] 				    int_h2c_gpio_11_gpio_22;
   wire [0:0] 				    int_h2c_gpio_11_gpio_21;
   wire [0:0] 				    int_h2c_gpio_11_gpio_20;
   wire [0:0] 				    int_h2c_gpio_11_gpio_19;
   wire [0:0] 				    int_h2c_gpio_11_gpio_18;
   wire [0:0] 				    int_h2c_gpio_11_gpio_17;
   wire [0:0] 				    int_h2c_gpio_11_gpio_16;
   wire [0:0] 				    int_h2c_gpio_11_gpio_15;
   wire [0:0] 				    int_h2c_gpio_11_gpio_14;
   wire [0:0] 				    int_h2c_gpio_11_gpio_13;
   wire [0:0] 				    int_h2c_gpio_11_gpio_12;
   wire [0:0] 				    int_h2c_gpio_11_gpio_11;
   wire [0:0] 				    int_h2c_gpio_11_gpio_10;
   wire [0:0] 				    int_h2c_gpio_11_gpio_9;
   wire [0:0] 				    int_h2c_gpio_11_gpio_8;
   wire [0:0] 				    int_h2c_gpio_11_gpio_7;
   wire [0:0] 				    int_h2c_gpio_11_gpio_6;
   wire [0:0] 				    int_h2c_gpio_11_gpio_5;
   wire [0:0] 				    int_h2c_gpio_11_gpio_4;
   wire [0:0] 				    int_h2c_gpio_11_gpio_3;
   wire [0:0] 				    int_h2c_gpio_11_gpio_2;
   wire [0:0] 				    int_h2c_gpio_11_gpio_1;
   wire [0:0] 				    int_h2c_gpio_11_gpio_0;
   wire [0:0] 				    int_h2c_gpio_12_gpio_31;
   wire [0:0] 				    int_h2c_gpio_12_gpio_30;
   wire [0:0] 				    int_h2c_gpio_12_gpio_29;
   wire [0:0] 				    int_h2c_gpio_12_gpio_28;
   wire [0:0] 				    int_h2c_gpio_12_gpio_27;
   wire [0:0] 				    int_h2c_gpio_12_gpio_26;
   wire [0:0] 				    int_h2c_gpio_12_gpio_25;
   wire [0:0] 				    int_h2c_gpio_12_gpio_24;
   wire [0:0] 				    int_h2c_gpio_12_gpio_23;
   wire [0:0] 				    int_h2c_gpio_12_gpio_22;
   wire [0:0] 				    int_h2c_gpio_12_gpio_21;
   wire [0:0] 				    int_h2c_gpio_12_gpio_20;
   wire [0:0] 				    int_h2c_gpio_12_gpio_19;
   wire [0:0] 				    int_h2c_gpio_12_gpio_18;
   wire [0:0] 				    int_h2c_gpio_12_gpio_17;
   wire [0:0] 				    int_h2c_gpio_12_gpio_16;
   wire [0:0] 				    int_h2c_gpio_12_gpio_15;
   wire [0:0] 				    int_h2c_gpio_12_gpio_14;
   wire [0:0] 				    int_h2c_gpio_12_gpio_13;
   wire [0:0] 				    int_h2c_gpio_12_gpio_12;
   wire [0:0] 				    int_h2c_gpio_12_gpio_11;
   wire [0:0] 				    int_h2c_gpio_12_gpio_10;
   wire [0:0] 				    int_h2c_gpio_12_gpio_9;
   wire [0:0] 				    int_h2c_gpio_12_gpio_8;
   wire [0:0] 				    int_h2c_gpio_12_gpio_7;
   wire [0:0] 				    int_h2c_gpio_12_gpio_6;
   wire [0:0] 				    int_h2c_gpio_12_gpio_5;
   wire [0:0] 				    int_h2c_gpio_12_gpio_4;
   wire [0:0] 				    int_h2c_gpio_12_gpio_3;
   wire [0:0] 				    int_h2c_gpio_12_gpio_2;
   wire [0:0] 				    int_h2c_gpio_12_gpio_1;
   wire [0:0] 				    int_h2c_gpio_12_gpio_0;
   wire [0:0] 				    int_h2c_gpio_13_gpio_31;
   wire [0:0] 				    int_h2c_gpio_13_gpio_30;
   wire [0:0] 				    int_h2c_gpio_13_gpio_29;
   wire [0:0] 				    int_h2c_gpio_13_gpio_28;
   wire [0:0] 				    int_h2c_gpio_13_gpio_27;
   wire [0:0] 				    int_h2c_gpio_13_gpio_26;
   wire [0:0] 				    int_h2c_gpio_13_gpio_25;
   wire [0:0] 				    int_h2c_gpio_13_gpio_24;
   wire [0:0] 				    int_h2c_gpio_13_gpio_23;
   wire [0:0] 				    int_h2c_gpio_13_gpio_22;
   wire [0:0] 				    int_h2c_gpio_13_gpio_21;
   wire [0:0] 				    int_h2c_gpio_13_gpio_20;
   wire [0:0] 				    int_h2c_gpio_13_gpio_19;
   wire [0:0] 				    int_h2c_gpio_13_gpio_18;
   wire [0:0] 				    int_h2c_gpio_13_gpio_17;
   wire [0:0] 				    int_h2c_gpio_13_gpio_16;
   wire [0:0] 				    int_h2c_gpio_13_gpio_15;
   wire [0:0] 				    int_h2c_gpio_13_gpio_14;
   wire [0:0] 				    int_h2c_gpio_13_gpio_13;
   wire [0:0] 				    int_h2c_gpio_13_gpio_12;
   wire [0:0] 				    int_h2c_gpio_13_gpio_11;
   wire [0:0] 				    int_h2c_gpio_13_gpio_10;
   wire [0:0] 				    int_h2c_gpio_13_gpio_9;
   wire [0:0] 				    int_h2c_gpio_13_gpio_8;
   wire [0:0] 				    int_h2c_gpio_13_gpio_7;
   wire [0:0] 				    int_h2c_gpio_13_gpio_6;
   wire [0:0] 				    int_h2c_gpio_13_gpio_5;
   wire [0:0] 				    int_h2c_gpio_13_gpio_4;
   wire [0:0] 				    int_h2c_gpio_13_gpio_3;
   wire [0:0] 				    int_h2c_gpio_13_gpio_2;
   wire [0:0] 				    int_h2c_gpio_13_gpio_1;
   wire [0:0] 				    int_h2c_gpio_13_gpio_0;
   wire [0:0] 				    int_h2c_gpio_14_gpio_31;
   wire [0:0] 				    int_h2c_gpio_14_gpio_30;
   wire [0:0] 				    int_h2c_gpio_14_gpio_29;
   wire [0:0] 				    int_h2c_gpio_14_gpio_28;
   wire [0:0] 				    int_h2c_gpio_14_gpio_27;
   wire [0:0] 				    int_h2c_gpio_14_gpio_26;
   wire [0:0] 				    int_h2c_gpio_14_gpio_25;
   wire [0:0] 				    int_h2c_gpio_14_gpio_24;
   wire [0:0] 				    int_h2c_gpio_14_gpio_23;
   wire [0:0] 				    int_h2c_gpio_14_gpio_22;
   wire [0:0] 				    int_h2c_gpio_14_gpio_21;
   wire [0:0] 				    int_h2c_gpio_14_gpio_20;
   wire [0:0] 				    int_h2c_gpio_14_gpio_19;
   wire [0:0] 				    int_h2c_gpio_14_gpio_18;
   wire [0:0] 				    int_h2c_gpio_14_gpio_17;
   wire [0:0] 				    int_h2c_gpio_14_gpio_16;
   wire [0:0] 				    int_h2c_gpio_14_gpio_15;
   wire [0:0] 				    int_h2c_gpio_14_gpio_14;
   wire [0:0] 				    int_h2c_gpio_14_gpio_13;
   wire [0:0] 				    int_h2c_gpio_14_gpio_12;
   wire [0:0] 				    int_h2c_gpio_14_gpio_11;
   wire [0:0] 				    int_h2c_gpio_14_gpio_10;
   wire [0:0] 				    int_h2c_gpio_14_gpio_9;
   wire [0:0] 				    int_h2c_gpio_14_gpio_8;
   wire [0:0] 				    int_h2c_gpio_14_gpio_7;
   wire [0:0] 				    int_h2c_gpio_14_gpio_6;
   wire [0:0] 				    int_h2c_gpio_14_gpio_5;
   wire [0:0] 				    int_h2c_gpio_14_gpio_4;
   wire [0:0] 				    int_h2c_gpio_14_gpio_3;
   wire [0:0] 				    int_h2c_gpio_14_gpio_2;
   wire [0:0] 				    int_h2c_gpio_14_gpio_1;
   wire [0:0] 				    int_h2c_gpio_14_gpio_0;
   wire [0:0] 				    int_h2c_gpio_15_gpio_31;
   wire [0:0] 				    int_h2c_gpio_15_gpio_30;
   wire [0:0] 				    int_h2c_gpio_15_gpio_29;
   wire [0:0] 				    int_h2c_gpio_15_gpio_28;
   wire [0:0] 				    int_h2c_gpio_15_gpio_27;
   wire [0:0] 				    int_h2c_gpio_15_gpio_26;
   wire [0:0] 				    int_h2c_gpio_15_gpio_25;
   wire [0:0] 				    int_h2c_gpio_15_gpio_24;
   wire [0:0] 				    int_h2c_gpio_15_gpio_23;
   wire [0:0] 				    int_h2c_gpio_15_gpio_22;
   wire [0:0] 				    int_h2c_gpio_15_gpio_21;
   wire [0:0] 				    int_h2c_gpio_15_gpio_20;
   wire [0:0] 				    int_h2c_gpio_15_gpio_19;
   wire [0:0] 				    int_h2c_gpio_15_gpio_18;
   wire [0:0] 				    int_h2c_gpio_15_gpio_17;
   wire [0:0] 				    int_h2c_gpio_15_gpio_16;
   wire [0:0] 				    int_h2c_gpio_15_gpio_15;
   wire [0:0] 				    int_h2c_gpio_15_gpio_14;
   wire [0:0] 				    int_h2c_gpio_15_gpio_13;
   wire [0:0] 				    int_h2c_gpio_15_gpio_12;
   wire [0:0] 				    int_h2c_gpio_15_gpio_11;
   wire [0:0] 				    int_h2c_gpio_15_gpio_10;
   wire [0:0] 				    int_h2c_gpio_15_gpio_9;
   wire [0:0] 				    int_h2c_gpio_15_gpio_8;
   wire [0:0] 				    int_h2c_gpio_15_gpio_7;
   wire [0:0] 				    int_h2c_gpio_15_gpio_6;
   wire [0:0] 				    int_h2c_gpio_15_gpio_5;
   wire [0:0] 				    int_h2c_gpio_15_gpio_4;
   wire [0:0] 				    int_h2c_gpio_15_gpio_3;
   wire [0:0] 				    int_h2c_gpio_15_gpio_2;
   wire [0:0] 				    int_h2c_gpio_15_gpio_1;
   wire [0:0] 				    int_h2c_gpio_15_gpio_0;
   wire [31:0] 				    int_rd_req_desc_0_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_0_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_0_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_0_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_0_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_0_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_0_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_0_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_0_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_0_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_0_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_0_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_0_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_0_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_0_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_0_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_0_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_0_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_0_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_0_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_0_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_0_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_0_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_0_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_0_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_0_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_0_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_0_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_0_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_0_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_0_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_0_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_0_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_0_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_0_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_0_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_0_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_0_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_0_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_0_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_0_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_0_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_0_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_0_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_0_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_0_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_0_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_0_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_0_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_0_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_0_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_0_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_0_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_0_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_0_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_0_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_0_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_0_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_0_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_0_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_0_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_0_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_0_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_0_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_0_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_0_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_0_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_0_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_0_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_0_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_0_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_0_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_0_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_0_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_0_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_0_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_0_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_0_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_0_resp_resp;
   wire [31:0] 				    int_rd_req_desc_1_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_1_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_1_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_1_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_1_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_1_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_1_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_1_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_1_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_1_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_1_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_1_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_1_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_1_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_1_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_1_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_1_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_1_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_1_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_1_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_1_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_1_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_1_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_1_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_1_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_1_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_1_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_1_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_1_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_1_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_1_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_1_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_1_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_1_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_1_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_1_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_1_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_1_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_1_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_1_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_1_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_1_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_1_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_1_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_1_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_1_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_1_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_1_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_1_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_1_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_1_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_1_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_1_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_1_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_1_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_1_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_1_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_1_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_1_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_1_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_1_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_1_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_1_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_1_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_1_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_1_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_1_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_1_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_1_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_1_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_1_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_1_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_1_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_1_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_1_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_1_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_1_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_1_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_1_resp_resp;
   wire [31:0] 				    int_rd_req_desc_2_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_2_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_2_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_2_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_2_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_2_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_2_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_2_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_2_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_2_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_2_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_2_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_2_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_2_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_2_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_2_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_2_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_2_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_2_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_2_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_2_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_2_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_2_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_2_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_2_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_2_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_2_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_2_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_2_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_2_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_2_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_2_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_2_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_2_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_2_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_2_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_2_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_2_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_2_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_2_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_2_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_2_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_2_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_2_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_2_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_2_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_2_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_2_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_2_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_2_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_2_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_2_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_2_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_2_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_2_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_2_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_2_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_2_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_2_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_2_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_2_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_2_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_2_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_2_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_2_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_2_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_2_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_2_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_2_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_2_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_2_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_2_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_2_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_2_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_2_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_2_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_2_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_2_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_2_resp_resp;
   wire [31:0] 				    int_rd_req_desc_3_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_3_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_3_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_3_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_3_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_3_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_3_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_3_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_3_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_3_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_3_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_3_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_3_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_3_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_3_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_3_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_3_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_3_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_3_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_3_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_3_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_3_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_3_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_3_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_3_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_3_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_3_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_3_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_3_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_3_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_3_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_3_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_3_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_3_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_3_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_3_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_3_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_3_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_3_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_3_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_3_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_3_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_3_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_3_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_3_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_3_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_3_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_3_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_3_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_3_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_3_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_3_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_3_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_3_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_3_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_3_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_3_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_3_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_3_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_3_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_3_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_3_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_3_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_3_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_3_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_3_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_3_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_3_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_3_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_3_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_3_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_3_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_3_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_3_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_3_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_3_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_3_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_3_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_3_resp_resp;
   wire [31:0] 				    int_rd_req_desc_4_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_4_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_4_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_4_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_4_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_4_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_4_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_4_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_4_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_4_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_4_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_4_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_4_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_4_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_4_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_4_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_4_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_4_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_4_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_4_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_4_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_4_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_4_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_4_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_4_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_4_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_4_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_4_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_4_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_4_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_4_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_4_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_4_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_4_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_4_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_4_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_4_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_4_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_4_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_4_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_4_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_4_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_4_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_4_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_4_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_4_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_4_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_4_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_4_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_4_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_4_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_4_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_4_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_4_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_4_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_4_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_4_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_4_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_4_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_4_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_4_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_4_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_4_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_4_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_4_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_4_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_4_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_4_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_4_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_4_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_4_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_4_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_4_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_4_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_4_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_4_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_4_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_4_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_4_resp_resp;
   wire [31:0] 				    int_rd_req_desc_5_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_5_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_5_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_5_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_5_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_5_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_5_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_5_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_5_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_5_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_5_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_5_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_5_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_5_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_5_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_5_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_5_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_5_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_5_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_5_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_5_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_5_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_5_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_5_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_5_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_5_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_5_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_5_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_5_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_5_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_5_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_5_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_5_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_5_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_5_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_5_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_5_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_5_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_5_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_5_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_5_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_5_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_5_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_5_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_5_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_5_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_5_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_5_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_5_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_5_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_5_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_5_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_5_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_5_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_5_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_5_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_5_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_5_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_5_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_5_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_5_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_5_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_5_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_5_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_5_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_5_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_5_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_5_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_5_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_5_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_5_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_5_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_5_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_5_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_5_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_5_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_5_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_5_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_5_resp_resp;
   wire [31:0] 				    int_rd_req_desc_6_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_6_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_6_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_6_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_6_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_6_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_6_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_6_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_6_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_6_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_6_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_6_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_6_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_6_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_6_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_6_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_6_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_6_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_6_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_6_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_6_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_6_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_6_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_6_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_6_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_6_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_6_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_6_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_6_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_6_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_6_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_6_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_6_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_6_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_6_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_6_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_6_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_6_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_6_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_6_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_6_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_6_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_6_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_6_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_6_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_6_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_6_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_6_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_6_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_6_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_6_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_6_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_6_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_6_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_6_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_6_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_6_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_6_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_6_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_6_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_6_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_6_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_6_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_6_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_6_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_6_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_6_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_6_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_6_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_6_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_6_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_6_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_6_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_6_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_6_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_6_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_6_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_6_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_6_resp_resp;
   wire [31:0] 				    int_rd_req_desc_7_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_7_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_7_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_7_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_7_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_7_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_7_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_7_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_7_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_7_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_7_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_7_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_7_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_7_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_7_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_7_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_7_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_7_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_7_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_7_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_7_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_7_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_7_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_7_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_7_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_7_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_7_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_7_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_7_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_7_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_7_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_7_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_7_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_7_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_7_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_7_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_7_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_7_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_7_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_7_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_7_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_7_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_7_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_7_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_7_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_7_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_7_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_7_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_7_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_7_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_7_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_7_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_7_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_7_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_7_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_7_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_7_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_7_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_7_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_7_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_7_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_7_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_7_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_7_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_7_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_7_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_7_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_7_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_7_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_7_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_7_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_7_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_7_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_7_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_7_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_7_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_7_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_7_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_7_resp_resp;
   wire [31:0] 				    int_rd_req_desc_8_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_8_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_8_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_8_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_8_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_8_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_8_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_8_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_8_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_8_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_8_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_8_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_8_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_8_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_8_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_8_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_8_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_8_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_8_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_8_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_8_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_8_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_8_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_8_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_8_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_8_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_8_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_8_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_8_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_8_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_8_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_8_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_8_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_8_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_8_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_8_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_8_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_8_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_8_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_8_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_8_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_8_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_8_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_8_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_8_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_8_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_8_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_8_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_8_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_8_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_8_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_8_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_8_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_8_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_8_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_8_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_8_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_8_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_8_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_8_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_8_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_8_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_8_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_8_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_8_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_8_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_8_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_8_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_8_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_8_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_8_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_8_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_8_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_8_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_8_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_8_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_8_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_8_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_8_resp_resp;
   wire [31:0] 				    int_rd_req_desc_9_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_9_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_9_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_9_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_9_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_9_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_9_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_9_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_9_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_9_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_9_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_9_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_9_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_9_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_9_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_9_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_9_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_9_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_9_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_9_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_9_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_9_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_9_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_9_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_9_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_9_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_9_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_9_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_9_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_9_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_9_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_9_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_9_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_9_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_9_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_9_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_9_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_9_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_9_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_9_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_9_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_9_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_9_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_9_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_9_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_9_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_9_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_9_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_9_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_9_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_9_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_9_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_9_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_9_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_9_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_9_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_9_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_9_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_9_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_9_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_9_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_9_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_9_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_9_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_9_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_9_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_9_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_9_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_9_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_9_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_9_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_9_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_9_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_9_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_9_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_9_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_9_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_9_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_9_resp_resp;
   wire [31:0] 				    int_rd_req_desc_a_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_a_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_a_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_a_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_a_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_a_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_a_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_a_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_a_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_a_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_a_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_a_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_a_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_a_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_a_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_a_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_a_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_a_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_a_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_a_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_a_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_a_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_a_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_a_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_a_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_a_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_a_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_a_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_a_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_a_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_a_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_a_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_a_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_a_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_a_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_a_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_a_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_a_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_a_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_a_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_a_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_a_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_a_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_a_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_a_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_a_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_a_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_a_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_a_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_a_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_a_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_a_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_a_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_a_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_a_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_a_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_a_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_a_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_a_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_a_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_a_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_a_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_a_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_a_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_a_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_a_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_a_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_a_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_a_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_a_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_a_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_a_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_a_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_a_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_a_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_a_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_a_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_a_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_a_resp_resp;
   wire [31:0] 				    int_rd_req_desc_b_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_b_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_b_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_b_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_b_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_b_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_b_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_b_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_b_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_b_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_b_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_b_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_b_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_b_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_b_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_b_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_b_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_b_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_b_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_b_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_b_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_b_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_b_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_b_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_b_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_b_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_b_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_b_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_b_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_b_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_b_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_b_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_b_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_b_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_b_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_b_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_b_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_b_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_b_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_b_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_b_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_b_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_b_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_b_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_b_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_b_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_b_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_b_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_b_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_b_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_b_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_b_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_b_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_b_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_b_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_b_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_b_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_b_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_b_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_b_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_b_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_b_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_b_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_b_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_b_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_b_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_b_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_b_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_b_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_b_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_b_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_b_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_b_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_b_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_b_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_b_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_b_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_b_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_b_resp_resp;
   wire [31:0] 				    int_rd_req_desc_c_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_c_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_c_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_c_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_c_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_c_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_c_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_c_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_c_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_c_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_c_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_c_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_c_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_c_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_c_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_c_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_c_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_c_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_c_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_c_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_c_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_c_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_c_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_c_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_c_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_c_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_c_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_c_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_c_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_c_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_c_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_c_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_c_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_c_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_c_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_c_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_c_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_c_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_c_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_c_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_c_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_c_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_c_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_c_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_c_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_c_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_c_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_c_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_c_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_c_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_c_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_c_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_c_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_c_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_c_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_c_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_c_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_c_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_c_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_c_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_c_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_c_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_c_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_c_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_c_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_c_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_c_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_c_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_c_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_c_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_c_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_c_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_c_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_c_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_c_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_c_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_c_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_c_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_c_resp_resp;
   wire [31:0] 				    int_rd_req_desc_d_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_d_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_d_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_d_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_d_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_d_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_d_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_d_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_d_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_d_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_d_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_d_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_d_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_d_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_d_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_d_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_d_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_d_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_d_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_d_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_d_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_d_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_d_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_d_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_d_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_d_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_d_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_d_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_d_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_d_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_d_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_d_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_d_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_d_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_d_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_d_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_d_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_d_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_d_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_d_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_d_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_d_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_d_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_d_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_d_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_d_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_d_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_d_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_d_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_d_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_d_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_d_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_d_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_d_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_d_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_d_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_d_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_d_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_d_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_d_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_d_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_d_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_d_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_d_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_d_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_d_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_d_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_d_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_d_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_d_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_d_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_d_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_d_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_d_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_d_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_d_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_d_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_d_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_d_resp_resp;
   wire [31:0] 				    int_rd_req_desc_e_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_e_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_e_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_e_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_e_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_e_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_e_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_e_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_e_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_e_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_e_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_e_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_e_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_e_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_e_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_e_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_e_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_e_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_e_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_e_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_e_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_e_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_e_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_e_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_e_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_e_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_e_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_e_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_e_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_e_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_e_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_e_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_e_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_e_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_e_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_e_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_e_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_e_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_e_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_e_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_e_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_e_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_e_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_e_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_e_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_e_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_e_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_e_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_e_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_e_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_e_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_e_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_e_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_e_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_e_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_e_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_e_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_e_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_e_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_e_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_e_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_e_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_e_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_e_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_e_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_e_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_e_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_e_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_e_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_e_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_e_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_e_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_e_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_e_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_e_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_e_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_e_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_e_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_e_resp_resp;
   wire [31:0] 				    int_rd_req_desc_f_size_txn_size;
   wire [2:0] 				    int_rd_req_desc_f_axsize_axsize;
   wire [3:0] 				    int_rd_req_desc_f_attr_axsnoop;
   wire [1:0] 				    int_rd_req_desc_f_attr_axdomain;
   wire [1:0] 				    int_rd_req_desc_f_attr_axbar;
   wire [3:0] 				    int_rd_req_desc_f_attr_axregion;
   wire [3:0] 				    int_rd_req_desc_f_attr_axqos;
   wire [2:0] 				    int_rd_req_desc_f_attr_axprot;
   wire [3:0] 				    int_rd_req_desc_f_attr_axcache;
   wire [0:0] 				    int_rd_req_desc_f_attr_axlock;
   wire [1:0] 				    int_rd_req_desc_f_attr_axburst;
   wire [31:0] 				    int_rd_req_desc_f_axaddr_0_addr;
   wire [31:0] 				    int_rd_req_desc_f_axaddr_1_addr;
   wire [31:0] 				    int_rd_req_desc_f_axaddr_2_addr;
   wire [31:0] 				    int_rd_req_desc_f_axaddr_3_addr;
   wire [31:0] 				    int_rd_req_desc_f_axid_0_axid;
   wire [31:0] 				    int_rd_req_desc_f_axid_1_axid;
   wire [31:0] 				    int_rd_req_desc_f_axid_2_axid;
   wire [31:0] 				    int_rd_req_desc_f_axid_3_axid;
   wire [31:0] 				    int_rd_req_desc_f_axuser_0_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_1_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_2_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_3_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_4_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_5_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_6_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_7_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_8_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_9_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_10_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_11_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_12_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_13_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_14_axuser;
   wire [31:0] 				    int_rd_req_desc_f_axuser_15_axuser;
   wire [13:0] 				    int_rd_resp_desc_f_data_offset_addr;
   wire [31:0] 				    int_rd_resp_desc_f_data_size_size;
   wire [31:0] 				    int_rd_resp_desc_f_data_host_addr_0_addr;
   wire [31:0] 				    int_rd_resp_desc_f_data_host_addr_1_addr;
   wire [31:0] 				    int_rd_resp_desc_f_data_host_addr_2_addr;
   wire [31:0] 				    int_rd_resp_desc_f_data_host_addr_3_addr;
   wire [4:0] 				    int_rd_resp_desc_f_resp_resp;
   wire [31:0] 				    int_rd_resp_desc_f_xid_0_xid;
   wire [31:0] 				    int_rd_resp_desc_f_xid_1_xid;
   wire [31:0] 				    int_rd_resp_desc_f_xid_2_xid;
   wire [31:0] 				    int_rd_resp_desc_f_xid_3_xid;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_0_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_1_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_2_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_3_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_4_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_5_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_6_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_7_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_8_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_9_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_10_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_11_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_12_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_13_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_14_xuser;
   wire [31:0] 				    int_rd_resp_desc_f_xuser_15_xuser;
   wire [0:0] 				    int_wr_req_desc_f_txn_type_wr_strb;
   wire [31:0] 				    int_wr_req_desc_f_size_txn_size;
   wire [13:0] 				    int_wr_req_desc_f_data_offset_addr;
   wire [31:0] 				    int_wr_req_desc_f_data_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_f_data_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_f_data_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_f_data_host_addr_3_addr;
   wire [31:0] 				    int_wr_req_desc_f_wstrb_host_addr_0_addr;
   wire [31:0] 				    int_wr_req_desc_f_wstrb_host_addr_1_addr;
   wire [31:0] 				    int_wr_req_desc_f_wstrb_host_addr_2_addr;
   wire [31:0] 				    int_wr_req_desc_f_wstrb_host_addr_3_addr;
   wire [2:0] 				    int_wr_req_desc_f_axsize_axsize;
   wire [3:0] 				    int_wr_req_desc_f_attr_axsnoop;
   wire [1:0] 				    int_wr_req_desc_f_attr_axdomain;
   wire [1:0] 				    int_wr_req_desc_f_attr_axbar;
   wire [0:0] 				    int_wr_req_desc_f_attr_awunique;
   wire [3:0] 				    int_wr_req_desc_f_attr_axregion;
   wire [3:0] 				    int_wr_req_desc_f_attr_axqos;
   wire [2:0] 				    int_wr_req_desc_f_attr_axprot;
   wire [3:0] 				    int_wr_req_desc_f_attr_axcache;
   wire [0:0] 				    int_wr_req_desc_f_attr_axlock;
   wire [1:0] 				    int_wr_req_desc_f_attr_axburst;
   wire [31:0] 				    int_wr_req_desc_f_axaddr_0_addr;
   wire [31:0] 				    int_wr_req_desc_f_axaddr_1_addr;
   wire [31:0] 				    int_wr_req_desc_f_axaddr_2_addr;
   wire [31:0] 				    int_wr_req_desc_f_axaddr_3_addr;
   wire [31:0] 				    int_wr_req_desc_f_axid_0_axid;
   wire [31:0] 				    int_wr_req_desc_f_axid_1_axid;
   wire [31:0] 				    int_wr_req_desc_f_axid_2_axid;
   wire [31:0] 				    int_wr_req_desc_f_axid_3_axid;
   wire [31:0] 				    int_wr_req_desc_f_axuser_0_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_1_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_2_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_3_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_4_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_5_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_6_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_7_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_8_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_9_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_10_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_11_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_12_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_13_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_14_axuser;
   wire [31:0] 				    int_wr_req_desc_f_axuser_15_axuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_0_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_1_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_2_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_3_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_4_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_5_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_6_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_7_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_8_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_9_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_10_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_11_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_12_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_13_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_14_wuser;
   wire [31:0] 				    int_wr_req_desc_f_wuser_15_wuser;
   wire [4:0] 				    int_wr_resp_desc_f_resp_resp;
   wire [31:0] 				    int_wr_resp_desc_f_xid_0_xid;
   wire [31:0] 				    int_wr_resp_desc_f_xid_1_xid;
   wire [31:0] 				    int_wr_resp_desc_f_xid_2_xid;
   wire [31:0] 				    int_wr_resp_desc_f_xid_3_xid;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_0_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_1_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_2_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_3_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_4_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_5_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_6_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_7_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_8_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_9_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_10_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_11_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_12_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_13_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_14_xuser;
   wire [31:0] 				    int_wr_resp_desc_f_xuser_15_xuser;
   wire [3:0] 				    int_sn_req_desc_f_attr_acsnoop;
   wire [2:0] 				    int_sn_req_desc_f_attr_acprot;
   wire [31:0] 				    int_sn_req_desc_f_acaddr_0_addr;
   wire [31:0] 				    int_sn_req_desc_f_acaddr_1_addr;
   wire [31:0] 				    int_sn_req_desc_f_acaddr_2_addr;
   wire [31:0] 				    int_sn_req_desc_f_acaddr_3_addr;
   wire [4:0] 				    int_sn_resp_desc_f_resp_resp;


   //Derive fields from registers of RB

   assign bridge_identification_last_bridge_f = bridge_identification_reg[0];
   assign version_major_ver_f = version_reg[15:8];
   assign version_minor_ver_f = version_reg[7:0];
   assign bridge_type_type_f = bridge_type_reg[7:0];
   assign bridge_config_extend_wstrb_f = bridge_config_reg[12];
   assign bridge_config_id_width_f = bridge_config_reg[11:4];
   assign bridge_config_data_width_f = bridge_config_reg[2:0];
   assign bridge_rd_user_config_ruser_width_f = bridge_rd_user_config_reg[19:10];
   assign bridge_rd_user_config_aruser_width_f = bridge_rd_user_config_reg[9:0];
   assign bridge_wr_user_config_buser_width_f = bridge_wr_user_config_reg[29:20];
   assign bridge_wr_user_config_wuser_width_f = bridge_wr_user_config_reg[19:10];
   assign bridge_wr_user_config_awuser_width_f = bridge_wr_user_config_reg[9:0];
   assign rd_max_desc_resp_max_desc_f = rd_max_desc_reg[15:8];
   assign rd_max_desc_req_max_desc_f = rd_max_desc_reg[7:0];
   assign wr_max_desc_resp_max_desc_f = wr_max_desc_reg[15:8];
   assign wr_max_desc_req_max_desc_f = wr_max_desc_reg[7:0];
   assign sn_max_desc_data_max_desc_f = sn_max_desc_reg[23:16];
   assign sn_max_desc_resp_max_desc_f = sn_max_desc_reg[15:8];
   assign sn_max_desc_req_max_desc_f = sn_max_desc_reg[7:0];
   assign reset_dut_srst_3_f = reset_reg[4];
   assign reset_dut_srst_2_f = reset_reg[3];
   assign reset_dut_srst_1_f = reset_reg[2];
   assign reset_dut_srst_0_f = reset_reg[1];
   assign reset_srst_f = reset_reg[0];
   assign mode_select_mode_0_1_f = mode_select_reg[0];
   assign intr_status_sn_data_fifo_nonempty_f = intr_status_reg[10];
   assign intr_status_sn_resp_fifo_nonempty_f = intr_status_reg[9];
   assign intr_status_sn_req_comp_f = intr_status_reg[8];
   assign intr_status_wr_resp_comp_f = intr_status_reg[7];
   assign intr_status_wr_req_fifo_nonempty_f = intr_status_reg[6];
   assign intr_status_rd_resp_comp_f = intr_status_reg[5];
   assign intr_status_rd_req_fifo_nonempty_f = intr_status_reg[4];
   assign intr_status_c2h_f = intr_status_reg[2];
   assign intr_status_error_f = intr_status_reg[1];
   assign intr_error_status_err_1_f = intr_error_status_reg[1];
   assign intr_error_status_err_0_f = intr_error_status_reg[0];
   assign intr_error_clear_clr_err_2_f = intr_error_clear_reg[2];
   assign intr_error_clear_clr_err_1_f = intr_error_clear_reg[1];
   assign intr_error_clear_clr_err_0_f = intr_error_clear_reg[0];
   assign intr_error_enable_en_err_2_f = intr_error_enable_reg[2];
   assign intr_error_enable_en_err_1_f = intr_error_enable_reg[1];
   assign intr_error_enable_en_err_0_f = intr_error_enable_reg[0];
   assign rd_req_free_desc_desc_f = rd_req_free_desc_reg[15:0];
   assign rd_req_fifo_pop_desc_valid_f = rd_req_fifo_pop_desc_reg[31];
   assign rd_req_fifo_pop_desc_desc_index_f = rd_req_fifo_pop_desc_reg[3:0];
   assign rd_req_fifo_fill_level_fill_f = rd_req_fifo_fill_level_reg[4:0];
   assign rd_resp_fifo_push_desc_valid_f = rd_resp_fifo_push_desc_reg[31];
   assign rd_resp_fifo_push_desc_desc_index_f = rd_resp_fifo_push_desc_reg[3:0];
   assign rd_resp_fifo_free_level_free_f = rd_resp_fifo_free_level_reg[4:0];
   assign rd_resp_intr_comp_status_comp_f = rd_resp_intr_comp_status_reg[15:0];
   assign rd_resp_intr_comp_clear_clr_comp_f = rd_resp_intr_comp_clear_reg[15:0];
   assign rd_resp_intr_comp_enable_en_comp_f = rd_resp_intr_comp_enable_reg[15:0];
   assign wr_req_free_desc_desc_f = wr_req_free_desc_reg[15:0];
   assign wr_req_fifo_pop_desc_valid_f = wr_req_fifo_pop_desc_reg[31];
   assign wr_req_fifo_pop_desc_desc_index_f = wr_req_fifo_pop_desc_reg[3:0];
   assign wr_req_fifo_fill_level_fill_f = wr_req_fifo_fill_level_reg[4:0];
   assign wr_resp_fifo_push_desc_valid_f = wr_resp_fifo_push_desc_reg[31];
   assign wr_resp_fifo_push_desc_desc_index_f = wr_resp_fifo_push_desc_reg[3:0];
   assign wr_resp_fifo_free_level_free_f = wr_resp_fifo_free_level_reg[4:0];
   assign wr_resp_intr_comp_status_comp_f = wr_resp_intr_comp_status_reg[15:0];
   assign wr_resp_intr_comp_clear_clr_comp_f = wr_resp_intr_comp_clear_reg[15:0];
   assign wr_resp_intr_comp_enable_en_comp_f = wr_resp_intr_comp_enable_reg[15:0];
   assign sn_req_fifo_push_desc_valid_f = sn_req_fifo_push_desc_reg[31];
   assign sn_req_fifo_push_desc_desc_index_f = sn_req_fifo_push_desc_reg[3:0];
   assign sn_req_fifo_free_level_free_f = sn_req_fifo_free_level_reg[4:0];
   assign sn_req_intr_comp_status_comp_f = sn_req_intr_comp_status_reg[15:0];
   assign sn_req_intr_comp_clear_clr_comp_f = sn_req_intr_comp_clear_reg[15:0];
   assign sn_req_intr_comp_enable_en_comp_f = sn_req_intr_comp_enable_reg[15:0];
   assign sn_resp_free_desc_desc_f = sn_resp_free_desc_reg[15:0];
   assign sn_resp_fifo_pop_desc_valid_f = sn_resp_fifo_pop_desc_reg[31];
   assign sn_resp_fifo_pop_desc_desc_index_f = sn_resp_fifo_pop_desc_reg[3:0];
   assign sn_resp_fifo_fill_level_fill_f = sn_resp_fifo_fill_level_reg[4:0];
   assign sn_data_free_desc_desc_f = sn_data_free_desc_reg[15:0];
   assign sn_data_fifo_pop_desc_valid_f = sn_data_fifo_pop_desc_reg[31];
   assign sn_data_fifo_pop_desc_desc_index_f = sn_data_fifo_pop_desc_reg[3:0];
   assign sn_data_fifo_fill_level_fill_f = sn_data_fifo_fill_level_reg[4:0];
   assign intr_fifo_enable_en_sn_data_fifo_nonempty_f = intr_fifo_enable_reg[3];
   assign intr_fifo_enable_en_sn_resp_fifo_nonempty_f = intr_fifo_enable_reg[2];
   assign intr_fifo_enable_en_wr_req_fifo_nonempty_f = intr_fifo_enable_reg[1];
   assign intr_fifo_enable_en_rd_req_fifo_nonempty_f = intr_fifo_enable_reg[0];
   assign h2c_intr_0_h2c_31_f = h2c_intr_0_reg[31];
   assign h2c_intr_0_h2c_30_f = h2c_intr_0_reg[30];
   assign h2c_intr_0_h2c_29_f = h2c_intr_0_reg[29];
   assign h2c_intr_0_h2c_28_f = h2c_intr_0_reg[28];
   assign h2c_intr_0_h2c_27_f = h2c_intr_0_reg[27];
   assign h2c_intr_0_h2c_26_f = h2c_intr_0_reg[26];
   assign h2c_intr_0_h2c_25_f = h2c_intr_0_reg[25];
   assign h2c_intr_0_h2c_24_f = h2c_intr_0_reg[24];
   assign h2c_intr_0_h2c_23_f = h2c_intr_0_reg[23];
   assign h2c_intr_0_h2c_22_f = h2c_intr_0_reg[22];
   assign h2c_intr_0_h2c_21_f = h2c_intr_0_reg[21];
   assign h2c_intr_0_h2c_20_f = h2c_intr_0_reg[20];
   assign h2c_intr_0_h2c_19_f = h2c_intr_0_reg[19];
   assign h2c_intr_0_h2c_18_f = h2c_intr_0_reg[18];
   assign h2c_intr_0_h2c_17_f = h2c_intr_0_reg[17];
   assign h2c_intr_0_h2c_16_f = h2c_intr_0_reg[16];
   assign h2c_intr_0_h2c_15_f = h2c_intr_0_reg[15];
   assign h2c_intr_0_h2c_14_f = h2c_intr_0_reg[14];
   assign h2c_intr_0_h2c_13_f = h2c_intr_0_reg[13];
   assign h2c_intr_0_h2c_12_f = h2c_intr_0_reg[12];
   assign h2c_intr_0_h2c_11_f = h2c_intr_0_reg[11];
   assign h2c_intr_0_h2c_10_f = h2c_intr_0_reg[10];
   assign h2c_intr_0_h2c_9_f = h2c_intr_0_reg[9];
   assign h2c_intr_0_h2c_8_f = h2c_intr_0_reg[8];
   assign h2c_intr_0_h2c_7_f = h2c_intr_0_reg[7];
   assign h2c_intr_0_h2c_6_f = h2c_intr_0_reg[6];
   assign h2c_intr_0_h2c_5_f = h2c_intr_0_reg[5];
   assign h2c_intr_0_h2c_4_f = h2c_intr_0_reg[4];
   assign h2c_intr_0_h2c_3_f = h2c_intr_0_reg[3];
   assign h2c_intr_0_h2c_2_f = h2c_intr_0_reg[2];
   assign h2c_intr_0_h2c_1_f = h2c_intr_0_reg[1];
   assign h2c_intr_0_h2c_0_f = h2c_intr_0_reg[0];
   assign h2c_intr_1_h2c_31_f = h2c_intr_1_reg[31];
   assign h2c_intr_1_h2c_30_f = h2c_intr_1_reg[30];
   assign h2c_intr_1_h2c_29_f = h2c_intr_1_reg[29];
   assign h2c_intr_1_h2c_28_f = h2c_intr_1_reg[28];
   assign h2c_intr_1_h2c_27_f = h2c_intr_1_reg[27];
   assign h2c_intr_1_h2c_26_f = h2c_intr_1_reg[26];
   assign h2c_intr_1_h2c_25_f = h2c_intr_1_reg[25];
   assign h2c_intr_1_h2c_24_f = h2c_intr_1_reg[24];
   assign h2c_intr_1_h2c_23_f = h2c_intr_1_reg[23];
   assign h2c_intr_1_h2c_22_f = h2c_intr_1_reg[22];
   assign h2c_intr_1_h2c_21_f = h2c_intr_1_reg[21];
   assign h2c_intr_1_h2c_20_f = h2c_intr_1_reg[20];
   assign h2c_intr_1_h2c_19_f = h2c_intr_1_reg[19];
   assign h2c_intr_1_h2c_18_f = h2c_intr_1_reg[18];
   assign h2c_intr_1_h2c_17_f = h2c_intr_1_reg[17];
   assign h2c_intr_1_h2c_16_f = h2c_intr_1_reg[16];
   assign h2c_intr_1_h2c_15_f = h2c_intr_1_reg[15];
   assign h2c_intr_1_h2c_14_f = h2c_intr_1_reg[14];
   assign h2c_intr_1_h2c_13_f = h2c_intr_1_reg[13];
   assign h2c_intr_1_h2c_12_f = h2c_intr_1_reg[12];
   assign h2c_intr_1_h2c_11_f = h2c_intr_1_reg[11];
   assign h2c_intr_1_h2c_10_f = h2c_intr_1_reg[10];
   assign h2c_intr_1_h2c_9_f = h2c_intr_1_reg[9];
   assign h2c_intr_1_h2c_8_f = h2c_intr_1_reg[8];
   assign h2c_intr_1_h2c_7_f = h2c_intr_1_reg[7];
   assign h2c_intr_1_h2c_6_f = h2c_intr_1_reg[6];
   assign h2c_intr_1_h2c_5_f = h2c_intr_1_reg[5];
   assign h2c_intr_1_h2c_4_f = h2c_intr_1_reg[4];
   assign h2c_intr_1_h2c_3_f = h2c_intr_1_reg[3];
   assign h2c_intr_1_h2c_2_f = h2c_intr_1_reg[2];
   assign h2c_intr_1_h2c_1_f = h2c_intr_1_reg[1];
   assign h2c_intr_1_h2c_0_f = h2c_intr_1_reg[0];
   assign h2c_intr_2_h2c_31_f = h2c_intr_2_reg[31];
   assign h2c_intr_2_h2c_30_f = h2c_intr_2_reg[30];
   assign h2c_intr_2_h2c_29_f = h2c_intr_2_reg[29];
   assign h2c_intr_2_h2c_28_f = h2c_intr_2_reg[28];
   assign h2c_intr_2_h2c_27_f = h2c_intr_2_reg[27];
   assign h2c_intr_2_h2c_26_f = h2c_intr_2_reg[26];
   assign h2c_intr_2_h2c_25_f = h2c_intr_2_reg[25];
   assign h2c_intr_2_h2c_24_f = h2c_intr_2_reg[24];
   assign h2c_intr_2_h2c_23_f = h2c_intr_2_reg[23];
   assign h2c_intr_2_h2c_22_f = h2c_intr_2_reg[22];
   assign h2c_intr_2_h2c_21_f = h2c_intr_2_reg[21];
   assign h2c_intr_2_h2c_20_f = h2c_intr_2_reg[20];
   assign h2c_intr_2_h2c_19_f = h2c_intr_2_reg[19];
   assign h2c_intr_2_h2c_18_f = h2c_intr_2_reg[18];
   assign h2c_intr_2_h2c_17_f = h2c_intr_2_reg[17];
   assign h2c_intr_2_h2c_16_f = h2c_intr_2_reg[16];
   assign h2c_intr_2_h2c_15_f = h2c_intr_2_reg[15];
   assign h2c_intr_2_h2c_14_f = h2c_intr_2_reg[14];
   assign h2c_intr_2_h2c_13_f = h2c_intr_2_reg[13];
   assign h2c_intr_2_h2c_12_f = h2c_intr_2_reg[12];
   assign h2c_intr_2_h2c_11_f = h2c_intr_2_reg[11];
   assign h2c_intr_2_h2c_10_f = h2c_intr_2_reg[10];
   assign h2c_intr_2_h2c_9_f = h2c_intr_2_reg[9];
   assign h2c_intr_2_h2c_8_f = h2c_intr_2_reg[8];
   assign h2c_intr_2_h2c_7_f = h2c_intr_2_reg[7];
   assign h2c_intr_2_h2c_6_f = h2c_intr_2_reg[6];
   assign h2c_intr_2_h2c_5_f = h2c_intr_2_reg[5];
   assign h2c_intr_2_h2c_4_f = h2c_intr_2_reg[4];
   assign h2c_intr_2_h2c_3_f = h2c_intr_2_reg[3];
   assign h2c_intr_2_h2c_2_f = h2c_intr_2_reg[2];
   assign h2c_intr_2_h2c_1_f = h2c_intr_2_reg[1];
   assign h2c_intr_2_h2c_0_f = h2c_intr_2_reg[0];
   assign h2c_intr_3_h2c_31_f = h2c_intr_3_reg[31];
   assign h2c_intr_3_h2c_30_f = h2c_intr_3_reg[30];
   assign h2c_intr_3_h2c_29_f = h2c_intr_3_reg[29];
   assign h2c_intr_3_h2c_28_f = h2c_intr_3_reg[28];
   assign h2c_intr_3_h2c_27_f = h2c_intr_3_reg[27];
   assign h2c_intr_3_h2c_26_f = h2c_intr_3_reg[26];
   assign h2c_intr_3_h2c_25_f = h2c_intr_3_reg[25];
   assign h2c_intr_3_h2c_24_f = h2c_intr_3_reg[24];
   assign h2c_intr_3_h2c_23_f = h2c_intr_3_reg[23];
   assign h2c_intr_3_h2c_22_f = h2c_intr_3_reg[22];
   assign h2c_intr_3_h2c_21_f = h2c_intr_3_reg[21];
   assign h2c_intr_3_h2c_20_f = h2c_intr_3_reg[20];
   assign h2c_intr_3_h2c_19_f = h2c_intr_3_reg[19];
   assign h2c_intr_3_h2c_18_f = h2c_intr_3_reg[18];
   assign h2c_intr_3_h2c_17_f = h2c_intr_3_reg[17];
   assign h2c_intr_3_h2c_16_f = h2c_intr_3_reg[16];
   assign h2c_intr_3_h2c_15_f = h2c_intr_3_reg[15];
   assign h2c_intr_3_h2c_14_f = h2c_intr_3_reg[14];
   assign h2c_intr_3_h2c_13_f = h2c_intr_3_reg[13];
   assign h2c_intr_3_h2c_12_f = h2c_intr_3_reg[12];
   assign h2c_intr_3_h2c_11_f = h2c_intr_3_reg[11];
   assign h2c_intr_3_h2c_10_f = h2c_intr_3_reg[10];
   assign h2c_intr_3_h2c_9_f = h2c_intr_3_reg[9];
   assign h2c_intr_3_h2c_8_f = h2c_intr_3_reg[8];
   assign h2c_intr_3_h2c_7_f = h2c_intr_3_reg[7];
   assign h2c_intr_3_h2c_6_f = h2c_intr_3_reg[6];
   assign h2c_intr_3_h2c_5_f = h2c_intr_3_reg[5];
   assign h2c_intr_3_h2c_4_f = h2c_intr_3_reg[4];
   assign h2c_intr_3_h2c_3_f = h2c_intr_3_reg[3];
   assign h2c_intr_3_h2c_2_f = h2c_intr_3_reg[2];
   assign h2c_intr_3_h2c_1_f = h2c_intr_3_reg[1];
   assign h2c_intr_3_h2c_0_f = h2c_intr_3_reg[0];
   assign c2h_intr_status_0_c2h_31_f = c2h_intr_status_0_reg[31];
   assign c2h_intr_status_0_c2h_30_f = c2h_intr_status_0_reg[30];
   assign c2h_intr_status_0_c2h_29_f = c2h_intr_status_0_reg[29];
   assign c2h_intr_status_0_c2h_28_f = c2h_intr_status_0_reg[28];
   assign c2h_intr_status_0_c2h_27_f = c2h_intr_status_0_reg[27];
   assign c2h_intr_status_0_c2h_26_f = c2h_intr_status_0_reg[26];
   assign c2h_intr_status_0_c2h_25_f = c2h_intr_status_0_reg[25];
   assign c2h_intr_status_0_c2h_24_f = c2h_intr_status_0_reg[24];
   assign c2h_intr_status_0_c2h_23_f = c2h_intr_status_0_reg[23];
   assign c2h_intr_status_0_c2h_22_f = c2h_intr_status_0_reg[22];
   assign c2h_intr_status_0_c2h_21_f = c2h_intr_status_0_reg[21];
   assign c2h_intr_status_0_c2h_20_f = c2h_intr_status_0_reg[20];
   assign c2h_intr_status_0_c2h_19_f = c2h_intr_status_0_reg[19];
   assign c2h_intr_status_0_c2h_18_f = c2h_intr_status_0_reg[18];
   assign c2h_intr_status_0_c2h_17_f = c2h_intr_status_0_reg[17];
   assign c2h_intr_status_0_c2h_16_f = c2h_intr_status_0_reg[16];
   assign c2h_intr_status_0_c2h_15_f = c2h_intr_status_0_reg[15];
   assign c2h_intr_status_0_c2h_14_f = c2h_intr_status_0_reg[14];
   assign c2h_intr_status_0_c2h_13_f = c2h_intr_status_0_reg[13];
   assign c2h_intr_status_0_c2h_12_f = c2h_intr_status_0_reg[12];
   assign c2h_intr_status_0_c2h_11_f = c2h_intr_status_0_reg[11];
   assign c2h_intr_status_0_c2h_10_f = c2h_intr_status_0_reg[10];
   assign c2h_intr_status_0_c2h_9_f = c2h_intr_status_0_reg[9];
   assign c2h_intr_status_0_c2h_8_f = c2h_intr_status_0_reg[8];
   assign c2h_intr_status_0_c2h_7_f = c2h_intr_status_0_reg[7];
   assign c2h_intr_status_0_c2h_6_f = c2h_intr_status_0_reg[6];
   assign c2h_intr_status_0_c2h_5_f = c2h_intr_status_0_reg[5];
   assign c2h_intr_status_0_c2h_4_f = c2h_intr_status_0_reg[4];
   assign c2h_intr_status_0_c2h_3_f = c2h_intr_status_0_reg[3];
   assign c2h_intr_status_0_c2h_2_f = c2h_intr_status_0_reg[2];
   assign c2h_intr_status_0_c2h_1_f = c2h_intr_status_0_reg[1];
   assign c2h_intr_status_0_c2h_0_f = c2h_intr_status_0_reg[0];
   assign intr_c2h_toggle_status_0_t_c2h_31_f = intr_c2h_toggle_status_0_reg[31];
   assign intr_c2h_toggle_status_0_t_c2h_30_f = intr_c2h_toggle_status_0_reg[30];
   assign intr_c2h_toggle_status_0_t_c2h_29_f = intr_c2h_toggle_status_0_reg[29];
   assign intr_c2h_toggle_status_0_t_c2h_28_f = intr_c2h_toggle_status_0_reg[28];
   assign intr_c2h_toggle_status_0_t_c2h_27_f = intr_c2h_toggle_status_0_reg[27];
   assign intr_c2h_toggle_status_0_t_c2h_26_f = intr_c2h_toggle_status_0_reg[26];
   assign intr_c2h_toggle_status_0_t_c2h_25_f = intr_c2h_toggle_status_0_reg[25];
   assign intr_c2h_toggle_status_0_t_c2h_24_f = intr_c2h_toggle_status_0_reg[24];
   assign intr_c2h_toggle_status_0_t_c2h_23_f = intr_c2h_toggle_status_0_reg[23];
   assign intr_c2h_toggle_status_0_t_c2h_22_f = intr_c2h_toggle_status_0_reg[22];
   assign intr_c2h_toggle_status_0_t_c2h_21_f = intr_c2h_toggle_status_0_reg[21];
   assign intr_c2h_toggle_status_0_t_c2h_20_f = intr_c2h_toggle_status_0_reg[20];
   assign intr_c2h_toggle_status_0_t_c2h_19_f = intr_c2h_toggle_status_0_reg[19];
   assign intr_c2h_toggle_status_0_t_c2h_18_f = intr_c2h_toggle_status_0_reg[18];
   assign intr_c2h_toggle_status_0_t_c2h_17_f = intr_c2h_toggle_status_0_reg[17];
   assign intr_c2h_toggle_status_0_t_c2h_16_f = intr_c2h_toggle_status_0_reg[16];
   assign intr_c2h_toggle_status_0_t_c2h_15_f = intr_c2h_toggle_status_0_reg[15];
   assign intr_c2h_toggle_status_0_t_c2h_14_f = intr_c2h_toggle_status_0_reg[14];
   assign intr_c2h_toggle_status_0_t_c2h_13_f = intr_c2h_toggle_status_0_reg[13];
   assign intr_c2h_toggle_status_0_t_c2h_12_f = intr_c2h_toggle_status_0_reg[12];
   assign intr_c2h_toggle_status_0_t_c2h_11_f = intr_c2h_toggle_status_0_reg[11];
   assign intr_c2h_toggle_status_0_t_c2h_10_f = intr_c2h_toggle_status_0_reg[10];
   assign intr_c2h_toggle_status_0_t_c2h_9_f = intr_c2h_toggle_status_0_reg[9];
   assign intr_c2h_toggle_status_0_t_c2h_8_f = intr_c2h_toggle_status_0_reg[8];
   assign intr_c2h_toggle_status_0_t_c2h_7_f = intr_c2h_toggle_status_0_reg[7];
   assign intr_c2h_toggle_status_0_t_c2h_6_f = intr_c2h_toggle_status_0_reg[6];
   assign intr_c2h_toggle_status_0_t_c2h_5_f = intr_c2h_toggle_status_0_reg[5];
   assign intr_c2h_toggle_status_0_t_c2h_4_f = intr_c2h_toggle_status_0_reg[4];
   assign intr_c2h_toggle_status_0_t_c2h_3_f = intr_c2h_toggle_status_0_reg[3];
   assign intr_c2h_toggle_status_0_t_c2h_2_f = intr_c2h_toggle_status_0_reg[2];
   assign intr_c2h_toggle_status_0_t_c2h_1_f = intr_c2h_toggle_status_0_reg[1];
   assign intr_c2h_toggle_status_0_t_c2h_0_f = intr_c2h_toggle_status_0_reg[0];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_31_f = intr_c2h_toggle_clear_0_reg[31];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_30_f = intr_c2h_toggle_clear_0_reg[30];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_29_f = intr_c2h_toggle_clear_0_reg[29];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_28_f = intr_c2h_toggle_clear_0_reg[28];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_27_f = intr_c2h_toggle_clear_0_reg[27];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_26_f = intr_c2h_toggle_clear_0_reg[26];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_25_f = intr_c2h_toggle_clear_0_reg[25];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_24_f = intr_c2h_toggle_clear_0_reg[24];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_23_f = intr_c2h_toggle_clear_0_reg[23];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_22_f = intr_c2h_toggle_clear_0_reg[22];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_21_f = intr_c2h_toggle_clear_0_reg[21];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_20_f = intr_c2h_toggle_clear_0_reg[20];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_19_f = intr_c2h_toggle_clear_0_reg[19];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_18_f = intr_c2h_toggle_clear_0_reg[18];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_17_f = intr_c2h_toggle_clear_0_reg[17];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_16_f = intr_c2h_toggle_clear_0_reg[16];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_15_f = intr_c2h_toggle_clear_0_reg[15];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_14_f = intr_c2h_toggle_clear_0_reg[14];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_13_f = intr_c2h_toggle_clear_0_reg[13];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_12_f = intr_c2h_toggle_clear_0_reg[12];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_11_f = intr_c2h_toggle_clear_0_reg[11];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_10_f = intr_c2h_toggle_clear_0_reg[10];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_9_f = intr_c2h_toggle_clear_0_reg[9];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_8_f = intr_c2h_toggle_clear_0_reg[8];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_7_f = intr_c2h_toggle_clear_0_reg[7];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_6_f = intr_c2h_toggle_clear_0_reg[6];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_5_f = intr_c2h_toggle_clear_0_reg[5];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_4_f = intr_c2h_toggle_clear_0_reg[4];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_3_f = intr_c2h_toggle_clear_0_reg[3];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_2_f = intr_c2h_toggle_clear_0_reg[2];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_1_f = intr_c2h_toggle_clear_0_reg[1];
   assign intr_c2h_toggle_clear_0_clr_t_c2h_0_f = intr_c2h_toggle_clear_0_reg[0];
   assign intr_c2h_toggle_enable_0_en_t_c2h_31_f = intr_c2h_toggle_enable_0_reg[31];
   assign intr_c2h_toggle_enable_0_en_t_c2h_30_f = intr_c2h_toggle_enable_0_reg[30];
   assign intr_c2h_toggle_enable_0_en_t_c2h_29_f = intr_c2h_toggle_enable_0_reg[29];
   assign intr_c2h_toggle_enable_0_en_t_c2h_28_f = intr_c2h_toggle_enable_0_reg[28];
   assign intr_c2h_toggle_enable_0_en_t_c2h_27_f = intr_c2h_toggle_enable_0_reg[27];
   assign intr_c2h_toggle_enable_0_en_t_c2h_26_f = intr_c2h_toggle_enable_0_reg[26];
   assign intr_c2h_toggle_enable_0_en_t_c2h_25_f = intr_c2h_toggle_enable_0_reg[25];
   assign intr_c2h_toggle_enable_0_en_t_c2h_24_f = intr_c2h_toggle_enable_0_reg[24];
   assign intr_c2h_toggle_enable_0_en_t_c2h_23_f = intr_c2h_toggle_enable_0_reg[23];
   assign intr_c2h_toggle_enable_0_en_t_c2h_22_f = intr_c2h_toggle_enable_0_reg[22];
   assign intr_c2h_toggle_enable_0_en_t_c2h_21_f = intr_c2h_toggle_enable_0_reg[21];
   assign intr_c2h_toggle_enable_0_en_t_c2h_20_f = intr_c2h_toggle_enable_0_reg[20];
   assign intr_c2h_toggle_enable_0_en_t_c2h_19_f = intr_c2h_toggle_enable_0_reg[19];
   assign intr_c2h_toggle_enable_0_en_t_c2h_18_f = intr_c2h_toggle_enable_0_reg[18];
   assign intr_c2h_toggle_enable_0_en_t_c2h_17_f = intr_c2h_toggle_enable_0_reg[17];
   assign intr_c2h_toggle_enable_0_en_t_c2h_16_f = intr_c2h_toggle_enable_0_reg[16];
   assign intr_c2h_toggle_enable_0_en_t_c2h_15_f = intr_c2h_toggle_enable_0_reg[15];
   assign intr_c2h_toggle_enable_0_en_t_c2h_14_f = intr_c2h_toggle_enable_0_reg[14];
   assign intr_c2h_toggle_enable_0_en_t_c2h_13_f = intr_c2h_toggle_enable_0_reg[13];
   assign intr_c2h_toggle_enable_0_en_t_c2h_12_f = intr_c2h_toggle_enable_0_reg[12];
   assign intr_c2h_toggle_enable_0_en_t_c2h_11_f = intr_c2h_toggle_enable_0_reg[11];
   assign intr_c2h_toggle_enable_0_en_t_c2h_10_f = intr_c2h_toggle_enable_0_reg[10];
   assign intr_c2h_toggle_enable_0_en_t_c2h_9_f = intr_c2h_toggle_enable_0_reg[9];
   assign intr_c2h_toggle_enable_0_en_t_c2h_8_f = intr_c2h_toggle_enable_0_reg[8];
   assign intr_c2h_toggle_enable_0_en_t_c2h_7_f = intr_c2h_toggle_enable_0_reg[7];
   assign intr_c2h_toggle_enable_0_en_t_c2h_6_f = intr_c2h_toggle_enable_0_reg[6];
   assign intr_c2h_toggle_enable_0_en_t_c2h_5_f = intr_c2h_toggle_enable_0_reg[5];
   assign intr_c2h_toggle_enable_0_en_t_c2h_4_f = intr_c2h_toggle_enable_0_reg[4];
   assign intr_c2h_toggle_enable_0_en_t_c2h_3_f = intr_c2h_toggle_enable_0_reg[3];
   assign intr_c2h_toggle_enable_0_en_t_c2h_2_f = intr_c2h_toggle_enable_0_reg[2];
   assign intr_c2h_toggle_enable_0_en_t_c2h_1_f = intr_c2h_toggle_enable_0_reg[1];
   assign intr_c2h_toggle_enable_0_en_t_c2h_0_f = intr_c2h_toggle_enable_0_reg[0];
   assign c2h_intr_status_1_c2h_31_f = c2h_intr_status_1_reg[31];
   assign c2h_intr_status_1_c2h_30_f = c2h_intr_status_1_reg[30];
   assign c2h_intr_status_1_c2h_29_f = c2h_intr_status_1_reg[29];
   assign c2h_intr_status_1_c2h_28_f = c2h_intr_status_1_reg[28];
   assign c2h_intr_status_1_c2h_27_f = c2h_intr_status_1_reg[27];
   assign c2h_intr_status_1_c2h_26_f = c2h_intr_status_1_reg[26];
   assign c2h_intr_status_1_c2h_25_f = c2h_intr_status_1_reg[25];
   assign c2h_intr_status_1_c2h_24_f = c2h_intr_status_1_reg[24];
   assign c2h_intr_status_1_c2h_23_f = c2h_intr_status_1_reg[23];
   assign c2h_intr_status_1_c2h_22_f = c2h_intr_status_1_reg[22];
   assign c2h_intr_status_1_c2h_21_f = c2h_intr_status_1_reg[21];
   assign c2h_intr_status_1_c2h_20_f = c2h_intr_status_1_reg[20];
   assign c2h_intr_status_1_c2h_19_f = c2h_intr_status_1_reg[19];
   assign c2h_intr_status_1_c2h_18_f = c2h_intr_status_1_reg[18];
   assign c2h_intr_status_1_c2h_17_f = c2h_intr_status_1_reg[17];
   assign c2h_intr_status_1_c2h_16_f = c2h_intr_status_1_reg[16];
   assign c2h_intr_status_1_c2h_15_f = c2h_intr_status_1_reg[15];
   assign c2h_intr_status_1_c2h_14_f = c2h_intr_status_1_reg[14];
   assign c2h_intr_status_1_c2h_13_f = c2h_intr_status_1_reg[13];
   assign c2h_intr_status_1_c2h_12_f = c2h_intr_status_1_reg[12];
   assign c2h_intr_status_1_c2h_11_f = c2h_intr_status_1_reg[11];
   assign c2h_intr_status_1_c2h_10_f = c2h_intr_status_1_reg[10];
   assign c2h_intr_status_1_c2h_9_f = c2h_intr_status_1_reg[9];
   assign c2h_intr_status_1_c2h_8_f = c2h_intr_status_1_reg[8];
   assign c2h_intr_status_1_c2h_7_f = c2h_intr_status_1_reg[7];
   assign c2h_intr_status_1_c2h_6_f = c2h_intr_status_1_reg[6];
   assign c2h_intr_status_1_c2h_5_f = c2h_intr_status_1_reg[5];
   assign c2h_intr_status_1_c2h_4_f = c2h_intr_status_1_reg[4];
   assign c2h_intr_status_1_c2h_3_f = c2h_intr_status_1_reg[3];
   assign c2h_intr_status_1_c2h_2_f = c2h_intr_status_1_reg[2];
   assign c2h_intr_status_1_c2h_1_f = c2h_intr_status_1_reg[1];
   assign c2h_intr_status_1_c2h_0_f = c2h_intr_status_1_reg[0];
   assign intr_c2h_toggle_status_1_t_c2h_31_f = intr_c2h_toggle_status_1_reg[31];
   assign intr_c2h_toggle_status_1_t_c2h_30_f = intr_c2h_toggle_status_1_reg[30];
   assign intr_c2h_toggle_status_1_t_c2h_29_f = intr_c2h_toggle_status_1_reg[29];
   assign intr_c2h_toggle_status_1_t_c2h_28_f = intr_c2h_toggle_status_1_reg[28];
   assign intr_c2h_toggle_status_1_t_c2h_27_f = intr_c2h_toggle_status_1_reg[27];
   assign intr_c2h_toggle_status_1_t_c2h_26_f = intr_c2h_toggle_status_1_reg[26];
   assign intr_c2h_toggle_status_1_t_c2h_25_f = intr_c2h_toggle_status_1_reg[25];
   assign intr_c2h_toggle_status_1_t_c2h_24_f = intr_c2h_toggle_status_1_reg[24];
   assign intr_c2h_toggle_status_1_t_c2h_23_f = intr_c2h_toggle_status_1_reg[23];
   assign intr_c2h_toggle_status_1_t_c2h_22_f = intr_c2h_toggle_status_1_reg[22];
   assign intr_c2h_toggle_status_1_t_c2h_21_f = intr_c2h_toggle_status_1_reg[21];
   assign intr_c2h_toggle_status_1_t_c2h_20_f = intr_c2h_toggle_status_1_reg[20];
   assign intr_c2h_toggle_status_1_t_c2h_19_f = intr_c2h_toggle_status_1_reg[19];
   assign intr_c2h_toggle_status_1_t_c2h_18_f = intr_c2h_toggle_status_1_reg[18];
   assign intr_c2h_toggle_status_1_t_c2h_17_f = intr_c2h_toggle_status_1_reg[17];
   assign intr_c2h_toggle_status_1_t_c2h_16_f = intr_c2h_toggle_status_1_reg[16];
   assign intr_c2h_toggle_status_1_t_c2h_15_f = intr_c2h_toggle_status_1_reg[15];
   assign intr_c2h_toggle_status_1_t_c2h_14_f = intr_c2h_toggle_status_1_reg[14];
   assign intr_c2h_toggle_status_1_t_c2h_13_f = intr_c2h_toggle_status_1_reg[13];
   assign intr_c2h_toggle_status_1_t_c2h_12_f = intr_c2h_toggle_status_1_reg[12];
   assign intr_c2h_toggle_status_1_t_c2h_11_f = intr_c2h_toggle_status_1_reg[11];
   assign intr_c2h_toggle_status_1_t_c2h_10_f = intr_c2h_toggle_status_1_reg[10];
   assign intr_c2h_toggle_status_1_t_c2h_9_f = intr_c2h_toggle_status_1_reg[9];
   assign intr_c2h_toggle_status_1_t_c2h_8_f = intr_c2h_toggle_status_1_reg[8];
   assign intr_c2h_toggle_status_1_t_c2h_7_f = intr_c2h_toggle_status_1_reg[7];
   assign intr_c2h_toggle_status_1_t_c2h_6_f = intr_c2h_toggle_status_1_reg[6];
   assign intr_c2h_toggle_status_1_t_c2h_5_f = intr_c2h_toggle_status_1_reg[5];
   assign intr_c2h_toggle_status_1_t_c2h_4_f = intr_c2h_toggle_status_1_reg[4];
   assign intr_c2h_toggle_status_1_t_c2h_3_f = intr_c2h_toggle_status_1_reg[3];
   assign intr_c2h_toggle_status_1_t_c2h_2_f = intr_c2h_toggle_status_1_reg[2];
   assign intr_c2h_toggle_status_1_t_c2h_1_f = intr_c2h_toggle_status_1_reg[1];
   assign intr_c2h_toggle_status_1_t_c2h_0_f = intr_c2h_toggle_status_1_reg[0];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_31_f = intr_c2h_toggle_clear_1_reg[31];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_30_f = intr_c2h_toggle_clear_1_reg[30];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_29_f = intr_c2h_toggle_clear_1_reg[29];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_28_f = intr_c2h_toggle_clear_1_reg[28];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_27_f = intr_c2h_toggle_clear_1_reg[27];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_26_f = intr_c2h_toggle_clear_1_reg[26];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_25_f = intr_c2h_toggle_clear_1_reg[25];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_24_f = intr_c2h_toggle_clear_1_reg[24];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_23_f = intr_c2h_toggle_clear_1_reg[23];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_22_f = intr_c2h_toggle_clear_1_reg[22];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_21_f = intr_c2h_toggle_clear_1_reg[21];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_20_f = intr_c2h_toggle_clear_1_reg[20];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_19_f = intr_c2h_toggle_clear_1_reg[19];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_18_f = intr_c2h_toggle_clear_1_reg[18];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_17_f = intr_c2h_toggle_clear_1_reg[17];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_16_f = intr_c2h_toggle_clear_1_reg[16];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_15_f = intr_c2h_toggle_clear_1_reg[15];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_14_f = intr_c2h_toggle_clear_1_reg[14];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_13_f = intr_c2h_toggle_clear_1_reg[13];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_12_f = intr_c2h_toggle_clear_1_reg[12];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_11_f = intr_c2h_toggle_clear_1_reg[11];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_10_f = intr_c2h_toggle_clear_1_reg[10];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_9_f = intr_c2h_toggle_clear_1_reg[9];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_8_f = intr_c2h_toggle_clear_1_reg[8];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_7_f = intr_c2h_toggle_clear_1_reg[7];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_6_f = intr_c2h_toggle_clear_1_reg[6];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_5_f = intr_c2h_toggle_clear_1_reg[5];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_4_f = intr_c2h_toggle_clear_1_reg[4];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_3_f = intr_c2h_toggle_clear_1_reg[3];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_2_f = intr_c2h_toggle_clear_1_reg[2];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_1_f = intr_c2h_toggle_clear_1_reg[1];
   assign intr_c2h_toggle_clear_1_clr_t_c2h_0_f = intr_c2h_toggle_clear_1_reg[0];
   assign intr_c2h_toggle_enable_1_en_t_c2h_31_f = intr_c2h_toggle_enable_1_reg[31];
   assign intr_c2h_toggle_enable_1_en_t_c2h_30_f = intr_c2h_toggle_enable_1_reg[30];
   assign intr_c2h_toggle_enable_1_en_t_c2h_29_f = intr_c2h_toggle_enable_1_reg[29];
   assign intr_c2h_toggle_enable_1_en_t_c2h_28_f = intr_c2h_toggle_enable_1_reg[28];
   assign intr_c2h_toggle_enable_1_en_t_c2h_27_f = intr_c2h_toggle_enable_1_reg[27];
   assign intr_c2h_toggle_enable_1_en_t_c2h_26_f = intr_c2h_toggle_enable_1_reg[26];
   assign intr_c2h_toggle_enable_1_en_t_c2h_25_f = intr_c2h_toggle_enable_1_reg[25];
   assign intr_c2h_toggle_enable_1_en_t_c2h_24_f = intr_c2h_toggle_enable_1_reg[24];
   assign intr_c2h_toggle_enable_1_en_t_c2h_23_f = intr_c2h_toggle_enable_1_reg[23];
   assign intr_c2h_toggle_enable_1_en_t_c2h_22_f = intr_c2h_toggle_enable_1_reg[22];
   assign intr_c2h_toggle_enable_1_en_t_c2h_21_f = intr_c2h_toggle_enable_1_reg[21];
   assign intr_c2h_toggle_enable_1_en_t_c2h_20_f = intr_c2h_toggle_enable_1_reg[20];
   assign intr_c2h_toggle_enable_1_en_t_c2h_19_f = intr_c2h_toggle_enable_1_reg[19];
   assign intr_c2h_toggle_enable_1_en_t_c2h_18_f = intr_c2h_toggle_enable_1_reg[18];
   assign intr_c2h_toggle_enable_1_en_t_c2h_17_f = intr_c2h_toggle_enable_1_reg[17];
   assign intr_c2h_toggle_enable_1_en_t_c2h_16_f = intr_c2h_toggle_enable_1_reg[16];
   assign intr_c2h_toggle_enable_1_en_t_c2h_15_f = intr_c2h_toggle_enable_1_reg[15];
   assign intr_c2h_toggle_enable_1_en_t_c2h_14_f = intr_c2h_toggle_enable_1_reg[14];
   assign intr_c2h_toggle_enable_1_en_t_c2h_13_f = intr_c2h_toggle_enable_1_reg[13];
   assign intr_c2h_toggle_enable_1_en_t_c2h_12_f = intr_c2h_toggle_enable_1_reg[12];
   assign intr_c2h_toggle_enable_1_en_t_c2h_11_f = intr_c2h_toggle_enable_1_reg[11];
   assign intr_c2h_toggle_enable_1_en_t_c2h_10_f = intr_c2h_toggle_enable_1_reg[10];
   assign intr_c2h_toggle_enable_1_en_t_c2h_9_f = intr_c2h_toggle_enable_1_reg[9];
   assign intr_c2h_toggle_enable_1_en_t_c2h_8_f = intr_c2h_toggle_enable_1_reg[8];
   assign intr_c2h_toggle_enable_1_en_t_c2h_7_f = intr_c2h_toggle_enable_1_reg[7];
   assign intr_c2h_toggle_enable_1_en_t_c2h_6_f = intr_c2h_toggle_enable_1_reg[6];
   assign intr_c2h_toggle_enable_1_en_t_c2h_5_f = intr_c2h_toggle_enable_1_reg[5];
   assign intr_c2h_toggle_enable_1_en_t_c2h_4_f = intr_c2h_toggle_enable_1_reg[4];
   assign intr_c2h_toggle_enable_1_en_t_c2h_3_f = intr_c2h_toggle_enable_1_reg[3];
   assign intr_c2h_toggle_enable_1_en_t_c2h_2_f = intr_c2h_toggle_enable_1_reg[2];
   assign intr_c2h_toggle_enable_1_en_t_c2h_1_f = intr_c2h_toggle_enable_1_reg[1];
   assign intr_c2h_toggle_enable_1_en_t_c2h_0_f = intr_c2h_toggle_enable_1_reg[0];
   assign c2h_gpio_0_gpio_31_f = c2h_gpio_0_reg[31];
   assign c2h_gpio_0_gpio_30_f = c2h_gpio_0_reg[30];
   assign c2h_gpio_0_gpio_29_f = c2h_gpio_0_reg[29];
   assign c2h_gpio_0_gpio_28_f = c2h_gpio_0_reg[28];
   assign c2h_gpio_0_gpio_27_f = c2h_gpio_0_reg[27];
   assign c2h_gpio_0_gpio_26_f = c2h_gpio_0_reg[26];
   assign c2h_gpio_0_gpio_25_f = c2h_gpio_0_reg[25];
   assign c2h_gpio_0_gpio_24_f = c2h_gpio_0_reg[24];
   assign c2h_gpio_0_gpio_23_f = c2h_gpio_0_reg[23];
   assign c2h_gpio_0_gpio_22_f = c2h_gpio_0_reg[22];
   assign c2h_gpio_0_gpio_21_f = c2h_gpio_0_reg[21];
   assign c2h_gpio_0_gpio_20_f = c2h_gpio_0_reg[20];
   assign c2h_gpio_0_gpio_19_f = c2h_gpio_0_reg[19];
   assign c2h_gpio_0_gpio_18_f = c2h_gpio_0_reg[18];
   assign c2h_gpio_0_gpio_17_f = c2h_gpio_0_reg[17];
   assign c2h_gpio_0_gpio_16_f = c2h_gpio_0_reg[16];
   assign c2h_gpio_0_gpio_15_f = c2h_gpio_0_reg[15];
   assign c2h_gpio_0_gpio_14_f = c2h_gpio_0_reg[14];
   assign c2h_gpio_0_gpio_13_f = c2h_gpio_0_reg[13];
   assign c2h_gpio_0_gpio_12_f = c2h_gpio_0_reg[12];
   assign c2h_gpio_0_gpio_11_f = c2h_gpio_0_reg[11];
   assign c2h_gpio_0_gpio_10_f = c2h_gpio_0_reg[10];
   assign c2h_gpio_0_gpio_9_f = c2h_gpio_0_reg[9];
   assign c2h_gpio_0_gpio_8_f = c2h_gpio_0_reg[8];
   assign c2h_gpio_0_gpio_7_f = c2h_gpio_0_reg[7];
   assign c2h_gpio_0_gpio_6_f = c2h_gpio_0_reg[6];
   assign c2h_gpio_0_gpio_5_f = c2h_gpio_0_reg[5];
   assign c2h_gpio_0_gpio_4_f = c2h_gpio_0_reg[4];
   assign c2h_gpio_0_gpio_3_f = c2h_gpio_0_reg[3];
   assign c2h_gpio_0_gpio_2_f = c2h_gpio_0_reg[2];
   assign c2h_gpio_0_gpio_1_f = c2h_gpio_0_reg[1];
   assign c2h_gpio_0_gpio_0_f = c2h_gpio_0_reg[0];
   assign c2h_gpio_1_gpio_31_f = c2h_gpio_1_reg[31];
   assign c2h_gpio_1_gpio_30_f = c2h_gpio_1_reg[30];
   assign c2h_gpio_1_gpio_29_f = c2h_gpio_1_reg[29];
   assign c2h_gpio_1_gpio_28_f = c2h_gpio_1_reg[28];
   assign c2h_gpio_1_gpio_27_f = c2h_gpio_1_reg[27];
   assign c2h_gpio_1_gpio_26_f = c2h_gpio_1_reg[26];
   assign c2h_gpio_1_gpio_25_f = c2h_gpio_1_reg[25];
   assign c2h_gpio_1_gpio_24_f = c2h_gpio_1_reg[24];
   assign c2h_gpio_1_gpio_23_f = c2h_gpio_1_reg[23];
   assign c2h_gpio_1_gpio_22_f = c2h_gpio_1_reg[22];
   assign c2h_gpio_1_gpio_21_f = c2h_gpio_1_reg[21];
   assign c2h_gpio_1_gpio_20_f = c2h_gpio_1_reg[20];
   assign c2h_gpio_1_gpio_19_f = c2h_gpio_1_reg[19];
   assign c2h_gpio_1_gpio_18_f = c2h_gpio_1_reg[18];
   assign c2h_gpio_1_gpio_17_f = c2h_gpio_1_reg[17];
   assign c2h_gpio_1_gpio_16_f = c2h_gpio_1_reg[16];
   assign c2h_gpio_1_gpio_15_f = c2h_gpio_1_reg[15];
   assign c2h_gpio_1_gpio_14_f = c2h_gpio_1_reg[14];
   assign c2h_gpio_1_gpio_13_f = c2h_gpio_1_reg[13];
   assign c2h_gpio_1_gpio_12_f = c2h_gpio_1_reg[12];
   assign c2h_gpio_1_gpio_11_f = c2h_gpio_1_reg[11];
   assign c2h_gpio_1_gpio_10_f = c2h_gpio_1_reg[10];
   assign c2h_gpio_1_gpio_9_f = c2h_gpio_1_reg[9];
   assign c2h_gpio_1_gpio_8_f = c2h_gpio_1_reg[8];
   assign c2h_gpio_1_gpio_7_f = c2h_gpio_1_reg[7];
   assign c2h_gpio_1_gpio_6_f = c2h_gpio_1_reg[6];
   assign c2h_gpio_1_gpio_5_f = c2h_gpio_1_reg[5];
   assign c2h_gpio_1_gpio_4_f = c2h_gpio_1_reg[4];
   assign c2h_gpio_1_gpio_3_f = c2h_gpio_1_reg[3];
   assign c2h_gpio_1_gpio_2_f = c2h_gpio_1_reg[2];
   assign c2h_gpio_1_gpio_1_f = c2h_gpio_1_reg[1];
   assign c2h_gpio_1_gpio_0_f = c2h_gpio_1_reg[0];
   assign c2h_gpio_2_gpio_31_f = c2h_gpio_2_reg[31];
   assign c2h_gpio_2_gpio_30_f = c2h_gpio_2_reg[30];
   assign c2h_gpio_2_gpio_29_f = c2h_gpio_2_reg[29];
   assign c2h_gpio_2_gpio_28_f = c2h_gpio_2_reg[28];
   assign c2h_gpio_2_gpio_27_f = c2h_gpio_2_reg[27];
   assign c2h_gpio_2_gpio_26_f = c2h_gpio_2_reg[26];
   assign c2h_gpio_2_gpio_25_f = c2h_gpio_2_reg[25];
   assign c2h_gpio_2_gpio_24_f = c2h_gpio_2_reg[24];
   assign c2h_gpio_2_gpio_23_f = c2h_gpio_2_reg[23];
   assign c2h_gpio_2_gpio_22_f = c2h_gpio_2_reg[22];
   assign c2h_gpio_2_gpio_21_f = c2h_gpio_2_reg[21];
   assign c2h_gpio_2_gpio_20_f = c2h_gpio_2_reg[20];
   assign c2h_gpio_2_gpio_19_f = c2h_gpio_2_reg[19];
   assign c2h_gpio_2_gpio_18_f = c2h_gpio_2_reg[18];
   assign c2h_gpio_2_gpio_17_f = c2h_gpio_2_reg[17];
   assign c2h_gpio_2_gpio_16_f = c2h_gpio_2_reg[16];
   assign c2h_gpio_2_gpio_15_f = c2h_gpio_2_reg[15];
   assign c2h_gpio_2_gpio_14_f = c2h_gpio_2_reg[14];
   assign c2h_gpio_2_gpio_13_f = c2h_gpio_2_reg[13];
   assign c2h_gpio_2_gpio_12_f = c2h_gpio_2_reg[12];
   assign c2h_gpio_2_gpio_11_f = c2h_gpio_2_reg[11];
   assign c2h_gpio_2_gpio_10_f = c2h_gpio_2_reg[10];
   assign c2h_gpio_2_gpio_9_f = c2h_gpio_2_reg[9];
   assign c2h_gpio_2_gpio_8_f = c2h_gpio_2_reg[8];
   assign c2h_gpio_2_gpio_7_f = c2h_gpio_2_reg[7];
   assign c2h_gpio_2_gpio_6_f = c2h_gpio_2_reg[6];
   assign c2h_gpio_2_gpio_5_f = c2h_gpio_2_reg[5];
   assign c2h_gpio_2_gpio_4_f = c2h_gpio_2_reg[4];
   assign c2h_gpio_2_gpio_3_f = c2h_gpio_2_reg[3];
   assign c2h_gpio_2_gpio_2_f = c2h_gpio_2_reg[2];
   assign c2h_gpio_2_gpio_1_f = c2h_gpio_2_reg[1];
   assign c2h_gpio_2_gpio_0_f = c2h_gpio_2_reg[0];
   assign c2h_gpio_3_gpio_31_f = c2h_gpio_3_reg[31];
   assign c2h_gpio_3_gpio_30_f = c2h_gpio_3_reg[30];
   assign c2h_gpio_3_gpio_29_f = c2h_gpio_3_reg[29];
   assign c2h_gpio_3_gpio_28_f = c2h_gpio_3_reg[28];
   assign c2h_gpio_3_gpio_27_f = c2h_gpio_3_reg[27];
   assign c2h_gpio_3_gpio_26_f = c2h_gpio_3_reg[26];
   assign c2h_gpio_3_gpio_25_f = c2h_gpio_3_reg[25];
   assign c2h_gpio_3_gpio_24_f = c2h_gpio_3_reg[24];
   assign c2h_gpio_3_gpio_23_f = c2h_gpio_3_reg[23];
   assign c2h_gpio_3_gpio_22_f = c2h_gpio_3_reg[22];
   assign c2h_gpio_3_gpio_21_f = c2h_gpio_3_reg[21];
   assign c2h_gpio_3_gpio_20_f = c2h_gpio_3_reg[20];
   assign c2h_gpio_3_gpio_19_f = c2h_gpio_3_reg[19];
   assign c2h_gpio_3_gpio_18_f = c2h_gpio_3_reg[18];
   assign c2h_gpio_3_gpio_17_f = c2h_gpio_3_reg[17];
   assign c2h_gpio_3_gpio_16_f = c2h_gpio_3_reg[16];
   assign c2h_gpio_3_gpio_15_f = c2h_gpio_3_reg[15];
   assign c2h_gpio_3_gpio_14_f = c2h_gpio_3_reg[14];
   assign c2h_gpio_3_gpio_13_f = c2h_gpio_3_reg[13];
   assign c2h_gpio_3_gpio_12_f = c2h_gpio_3_reg[12];
   assign c2h_gpio_3_gpio_11_f = c2h_gpio_3_reg[11];
   assign c2h_gpio_3_gpio_10_f = c2h_gpio_3_reg[10];
   assign c2h_gpio_3_gpio_9_f = c2h_gpio_3_reg[9];
   assign c2h_gpio_3_gpio_8_f = c2h_gpio_3_reg[8];
   assign c2h_gpio_3_gpio_7_f = c2h_gpio_3_reg[7];
   assign c2h_gpio_3_gpio_6_f = c2h_gpio_3_reg[6];
   assign c2h_gpio_3_gpio_5_f = c2h_gpio_3_reg[5];
   assign c2h_gpio_3_gpio_4_f = c2h_gpio_3_reg[4];
   assign c2h_gpio_3_gpio_3_f = c2h_gpio_3_reg[3];
   assign c2h_gpio_3_gpio_2_f = c2h_gpio_3_reg[2];
   assign c2h_gpio_3_gpio_1_f = c2h_gpio_3_reg[1];
   assign c2h_gpio_3_gpio_0_f = c2h_gpio_3_reg[0];
   assign c2h_gpio_4_gpio_31_f = c2h_gpio_4_reg[31];
   assign c2h_gpio_4_gpio_30_f = c2h_gpio_4_reg[30];
   assign c2h_gpio_4_gpio_29_f = c2h_gpio_4_reg[29];
   assign c2h_gpio_4_gpio_28_f = c2h_gpio_4_reg[28];
   assign c2h_gpio_4_gpio_27_f = c2h_gpio_4_reg[27];
   assign c2h_gpio_4_gpio_26_f = c2h_gpio_4_reg[26];
   assign c2h_gpio_4_gpio_25_f = c2h_gpio_4_reg[25];
   assign c2h_gpio_4_gpio_24_f = c2h_gpio_4_reg[24];
   assign c2h_gpio_4_gpio_23_f = c2h_gpio_4_reg[23];
   assign c2h_gpio_4_gpio_22_f = c2h_gpio_4_reg[22];
   assign c2h_gpio_4_gpio_21_f = c2h_gpio_4_reg[21];
   assign c2h_gpio_4_gpio_20_f = c2h_gpio_4_reg[20];
   assign c2h_gpio_4_gpio_19_f = c2h_gpio_4_reg[19];
   assign c2h_gpio_4_gpio_18_f = c2h_gpio_4_reg[18];
   assign c2h_gpio_4_gpio_17_f = c2h_gpio_4_reg[17];
   assign c2h_gpio_4_gpio_16_f = c2h_gpio_4_reg[16];
   assign c2h_gpio_4_gpio_15_f = c2h_gpio_4_reg[15];
   assign c2h_gpio_4_gpio_14_f = c2h_gpio_4_reg[14];
   assign c2h_gpio_4_gpio_13_f = c2h_gpio_4_reg[13];
   assign c2h_gpio_4_gpio_12_f = c2h_gpio_4_reg[12];
   assign c2h_gpio_4_gpio_11_f = c2h_gpio_4_reg[11];
   assign c2h_gpio_4_gpio_10_f = c2h_gpio_4_reg[10];
   assign c2h_gpio_4_gpio_9_f = c2h_gpio_4_reg[9];
   assign c2h_gpio_4_gpio_8_f = c2h_gpio_4_reg[8];
   assign c2h_gpio_4_gpio_7_f = c2h_gpio_4_reg[7];
   assign c2h_gpio_4_gpio_6_f = c2h_gpio_4_reg[6];
   assign c2h_gpio_4_gpio_5_f = c2h_gpio_4_reg[5];
   assign c2h_gpio_4_gpio_4_f = c2h_gpio_4_reg[4];
   assign c2h_gpio_4_gpio_3_f = c2h_gpio_4_reg[3];
   assign c2h_gpio_4_gpio_2_f = c2h_gpio_4_reg[2];
   assign c2h_gpio_4_gpio_1_f = c2h_gpio_4_reg[1];
   assign c2h_gpio_4_gpio_0_f = c2h_gpio_4_reg[0];
   assign c2h_gpio_5_gpio_31_f = c2h_gpio_5_reg[31];
   assign c2h_gpio_5_gpio_30_f = c2h_gpio_5_reg[30];
   assign c2h_gpio_5_gpio_29_f = c2h_gpio_5_reg[29];
   assign c2h_gpio_5_gpio_28_f = c2h_gpio_5_reg[28];
   assign c2h_gpio_5_gpio_27_f = c2h_gpio_5_reg[27];
   assign c2h_gpio_5_gpio_26_f = c2h_gpio_5_reg[26];
   assign c2h_gpio_5_gpio_25_f = c2h_gpio_5_reg[25];
   assign c2h_gpio_5_gpio_24_f = c2h_gpio_5_reg[24];
   assign c2h_gpio_5_gpio_23_f = c2h_gpio_5_reg[23];
   assign c2h_gpio_5_gpio_22_f = c2h_gpio_5_reg[22];
   assign c2h_gpio_5_gpio_21_f = c2h_gpio_5_reg[21];
   assign c2h_gpio_5_gpio_20_f = c2h_gpio_5_reg[20];
   assign c2h_gpio_5_gpio_19_f = c2h_gpio_5_reg[19];
   assign c2h_gpio_5_gpio_18_f = c2h_gpio_5_reg[18];
   assign c2h_gpio_5_gpio_17_f = c2h_gpio_5_reg[17];
   assign c2h_gpio_5_gpio_16_f = c2h_gpio_5_reg[16];
   assign c2h_gpio_5_gpio_15_f = c2h_gpio_5_reg[15];
   assign c2h_gpio_5_gpio_14_f = c2h_gpio_5_reg[14];
   assign c2h_gpio_5_gpio_13_f = c2h_gpio_5_reg[13];
   assign c2h_gpio_5_gpio_12_f = c2h_gpio_5_reg[12];
   assign c2h_gpio_5_gpio_11_f = c2h_gpio_5_reg[11];
   assign c2h_gpio_5_gpio_10_f = c2h_gpio_5_reg[10];
   assign c2h_gpio_5_gpio_9_f = c2h_gpio_5_reg[9];
   assign c2h_gpio_5_gpio_8_f = c2h_gpio_5_reg[8];
   assign c2h_gpio_5_gpio_7_f = c2h_gpio_5_reg[7];
   assign c2h_gpio_5_gpio_6_f = c2h_gpio_5_reg[6];
   assign c2h_gpio_5_gpio_5_f = c2h_gpio_5_reg[5];
   assign c2h_gpio_5_gpio_4_f = c2h_gpio_5_reg[4];
   assign c2h_gpio_5_gpio_3_f = c2h_gpio_5_reg[3];
   assign c2h_gpio_5_gpio_2_f = c2h_gpio_5_reg[2];
   assign c2h_gpio_5_gpio_1_f = c2h_gpio_5_reg[1];
   assign c2h_gpio_5_gpio_0_f = c2h_gpio_5_reg[0];
   assign c2h_gpio_6_gpio_31_f = c2h_gpio_6_reg[31];
   assign c2h_gpio_6_gpio_30_f = c2h_gpio_6_reg[30];
   assign c2h_gpio_6_gpio_29_f = c2h_gpio_6_reg[29];
   assign c2h_gpio_6_gpio_28_f = c2h_gpio_6_reg[28];
   assign c2h_gpio_6_gpio_27_f = c2h_gpio_6_reg[27];
   assign c2h_gpio_6_gpio_26_f = c2h_gpio_6_reg[26];
   assign c2h_gpio_6_gpio_25_f = c2h_gpio_6_reg[25];
   assign c2h_gpio_6_gpio_24_f = c2h_gpio_6_reg[24];
   assign c2h_gpio_6_gpio_23_f = c2h_gpio_6_reg[23];
   assign c2h_gpio_6_gpio_22_f = c2h_gpio_6_reg[22];
   assign c2h_gpio_6_gpio_21_f = c2h_gpio_6_reg[21];
   assign c2h_gpio_6_gpio_20_f = c2h_gpio_6_reg[20];
   assign c2h_gpio_6_gpio_19_f = c2h_gpio_6_reg[19];
   assign c2h_gpio_6_gpio_18_f = c2h_gpio_6_reg[18];
   assign c2h_gpio_6_gpio_17_f = c2h_gpio_6_reg[17];
   assign c2h_gpio_6_gpio_16_f = c2h_gpio_6_reg[16];
   assign c2h_gpio_6_gpio_15_f = c2h_gpio_6_reg[15];
   assign c2h_gpio_6_gpio_14_f = c2h_gpio_6_reg[14];
   assign c2h_gpio_6_gpio_13_f = c2h_gpio_6_reg[13];
   assign c2h_gpio_6_gpio_12_f = c2h_gpio_6_reg[12];
   assign c2h_gpio_6_gpio_11_f = c2h_gpio_6_reg[11];
   assign c2h_gpio_6_gpio_10_f = c2h_gpio_6_reg[10];
   assign c2h_gpio_6_gpio_9_f = c2h_gpio_6_reg[9];
   assign c2h_gpio_6_gpio_8_f = c2h_gpio_6_reg[8];
   assign c2h_gpio_6_gpio_7_f = c2h_gpio_6_reg[7];
   assign c2h_gpio_6_gpio_6_f = c2h_gpio_6_reg[6];
   assign c2h_gpio_6_gpio_5_f = c2h_gpio_6_reg[5];
   assign c2h_gpio_6_gpio_4_f = c2h_gpio_6_reg[4];
   assign c2h_gpio_6_gpio_3_f = c2h_gpio_6_reg[3];
   assign c2h_gpio_6_gpio_2_f = c2h_gpio_6_reg[2];
   assign c2h_gpio_6_gpio_1_f = c2h_gpio_6_reg[1];
   assign c2h_gpio_6_gpio_0_f = c2h_gpio_6_reg[0];
   assign c2h_gpio_7_gpio_31_f = c2h_gpio_7_reg[31];
   assign c2h_gpio_7_gpio_30_f = c2h_gpio_7_reg[30];
   assign c2h_gpio_7_gpio_29_f = c2h_gpio_7_reg[29];
   assign c2h_gpio_7_gpio_28_f = c2h_gpio_7_reg[28];
   assign c2h_gpio_7_gpio_27_f = c2h_gpio_7_reg[27];
   assign c2h_gpio_7_gpio_26_f = c2h_gpio_7_reg[26];
   assign c2h_gpio_7_gpio_25_f = c2h_gpio_7_reg[25];
   assign c2h_gpio_7_gpio_24_f = c2h_gpio_7_reg[24];
   assign c2h_gpio_7_gpio_23_f = c2h_gpio_7_reg[23];
   assign c2h_gpio_7_gpio_22_f = c2h_gpio_7_reg[22];
   assign c2h_gpio_7_gpio_21_f = c2h_gpio_7_reg[21];
   assign c2h_gpio_7_gpio_20_f = c2h_gpio_7_reg[20];
   assign c2h_gpio_7_gpio_19_f = c2h_gpio_7_reg[19];
   assign c2h_gpio_7_gpio_18_f = c2h_gpio_7_reg[18];
   assign c2h_gpio_7_gpio_17_f = c2h_gpio_7_reg[17];
   assign c2h_gpio_7_gpio_16_f = c2h_gpio_7_reg[16];
   assign c2h_gpio_7_gpio_15_f = c2h_gpio_7_reg[15];
   assign c2h_gpio_7_gpio_14_f = c2h_gpio_7_reg[14];
   assign c2h_gpio_7_gpio_13_f = c2h_gpio_7_reg[13];
   assign c2h_gpio_7_gpio_12_f = c2h_gpio_7_reg[12];
   assign c2h_gpio_7_gpio_11_f = c2h_gpio_7_reg[11];
   assign c2h_gpio_7_gpio_10_f = c2h_gpio_7_reg[10];
   assign c2h_gpio_7_gpio_9_f = c2h_gpio_7_reg[9];
   assign c2h_gpio_7_gpio_8_f = c2h_gpio_7_reg[8];
   assign c2h_gpio_7_gpio_7_f = c2h_gpio_7_reg[7];
   assign c2h_gpio_7_gpio_6_f = c2h_gpio_7_reg[6];
   assign c2h_gpio_7_gpio_5_f = c2h_gpio_7_reg[5];
   assign c2h_gpio_7_gpio_4_f = c2h_gpio_7_reg[4];
   assign c2h_gpio_7_gpio_3_f = c2h_gpio_7_reg[3];
   assign c2h_gpio_7_gpio_2_f = c2h_gpio_7_reg[2];
   assign c2h_gpio_7_gpio_1_f = c2h_gpio_7_reg[1];
   assign c2h_gpio_7_gpio_0_f = c2h_gpio_7_reg[0];
   assign c2h_gpio_8_gpio_31_f = c2h_gpio_8_reg[31];
   assign c2h_gpio_8_gpio_30_f = c2h_gpio_8_reg[30];
   assign c2h_gpio_8_gpio_29_f = c2h_gpio_8_reg[29];
   assign c2h_gpio_8_gpio_28_f = c2h_gpio_8_reg[28];
   assign c2h_gpio_8_gpio_27_f = c2h_gpio_8_reg[27];
   assign c2h_gpio_8_gpio_26_f = c2h_gpio_8_reg[26];
   assign c2h_gpio_8_gpio_25_f = c2h_gpio_8_reg[25];
   assign c2h_gpio_8_gpio_24_f = c2h_gpio_8_reg[24];
   assign c2h_gpio_8_gpio_23_f = c2h_gpio_8_reg[23];
   assign c2h_gpio_8_gpio_22_f = c2h_gpio_8_reg[22];
   assign c2h_gpio_8_gpio_21_f = c2h_gpio_8_reg[21];
   assign c2h_gpio_8_gpio_20_f = c2h_gpio_8_reg[20];
   assign c2h_gpio_8_gpio_19_f = c2h_gpio_8_reg[19];
   assign c2h_gpio_8_gpio_18_f = c2h_gpio_8_reg[18];
   assign c2h_gpio_8_gpio_17_f = c2h_gpio_8_reg[17];
   assign c2h_gpio_8_gpio_16_f = c2h_gpio_8_reg[16];
   assign c2h_gpio_8_gpio_15_f = c2h_gpio_8_reg[15];
   assign c2h_gpio_8_gpio_14_f = c2h_gpio_8_reg[14];
   assign c2h_gpio_8_gpio_13_f = c2h_gpio_8_reg[13];
   assign c2h_gpio_8_gpio_12_f = c2h_gpio_8_reg[12];
   assign c2h_gpio_8_gpio_11_f = c2h_gpio_8_reg[11];
   assign c2h_gpio_8_gpio_10_f = c2h_gpio_8_reg[10];
   assign c2h_gpio_8_gpio_9_f = c2h_gpio_8_reg[9];
   assign c2h_gpio_8_gpio_8_f = c2h_gpio_8_reg[8];
   assign c2h_gpio_8_gpio_7_f = c2h_gpio_8_reg[7];
   assign c2h_gpio_8_gpio_6_f = c2h_gpio_8_reg[6];
   assign c2h_gpio_8_gpio_5_f = c2h_gpio_8_reg[5];
   assign c2h_gpio_8_gpio_4_f = c2h_gpio_8_reg[4];
   assign c2h_gpio_8_gpio_3_f = c2h_gpio_8_reg[3];
   assign c2h_gpio_8_gpio_2_f = c2h_gpio_8_reg[2];
   assign c2h_gpio_8_gpio_1_f = c2h_gpio_8_reg[1];
   assign c2h_gpio_8_gpio_0_f = c2h_gpio_8_reg[0];
   assign c2h_gpio_9_gpio_31_f = c2h_gpio_9_reg[31];
   assign c2h_gpio_9_gpio_30_f = c2h_gpio_9_reg[30];
   assign c2h_gpio_9_gpio_29_f = c2h_gpio_9_reg[29];
   assign c2h_gpio_9_gpio_28_f = c2h_gpio_9_reg[28];
   assign c2h_gpio_9_gpio_27_f = c2h_gpio_9_reg[27];
   assign c2h_gpio_9_gpio_26_f = c2h_gpio_9_reg[26];
   assign c2h_gpio_9_gpio_25_f = c2h_gpio_9_reg[25];
   assign c2h_gpio_9_gpio_24_f = c2h_gpio_9_reg[24];
   assign c2h_gpio_9_gpio_23_f = c2h_gpio_9_reg[23];
   assign c2h_gpio_9_gpio_22_f = c2h_gpio_9_reg[22];
   assign c2h_gpio_9_gpio_21_f = c2h_gpio_9_reg[21];
   assign c2h_gpio_9_gpio_20_f = c2h_gpio_9_reg[20];
   assign c2h_gpio_9_gpio_19_f = c2h_gpio_9_reg[19];
   assign c2h_gpio_9_gpio_18_f = c2h_gpio_9_reg[18];
   assign c2h_gpio_9_gpio_17_f = c2h_gpio_9_reg[17];
   assign c2h_gpio_9_gpio_16_f = c2h_gpio_9_reg[16];
   assign c2h_gpio_9_gpio_15_f = c2h_gpio_9_reg[15];
   assign c2h_gpio_9_gpio_14_f = c2h_gpio_9_reg[14];
   assign c2h_gpio_9_gpio_13_f = c2h_gpio_9_reg[13];
   assign c2h_gpio_9_gpio_12_f = c2h_gpio_9_reg[12];
   assign c2h_gpio_9_gpio_11_f = c2h_gpio_9_reg[11];
   assign c2h_gpio_9_gpio_10_f = c2h_gpio_9_reg[10];
   assign c2h_gpio_9_gpio_9_f = c2h_gpio_9_reg[9];
   assign c2h_gpio_9_gpio_8_f = c2h_gpio_9_reg[8];
   assign c2h_gpio_9_gpio_7_f = c2h_gpio_9_reg[7];
   assign c2h_gpio_9_gpio_6_f = c2h_gpio_9_reg[6];
   assign c2h_gpio_9_gpio_5_f = c2h_gpio_9_reg[5];
   assign c2h_gpio_9_gpio_4_f = c2h_gpio_9_reg[4];
   assign c2h_gpio_9_gpio_3_f = c2h_gpio_9_reg[3];
   assign c2h_gpio_9_gpio_2_f = c2h_gpio_9_reg[2];
   assign c2h_gpio_9_gpio_1_f = c2h_gpio_9_reg[1];
   assign c2h_gpio_9_gpio_0_f = c2h_gpio_9_reg[0];
   assign c2h_gpio_10_gpio_31_f = c2h_gpio_10_reg[31];
   assign c2h_gpio_10_gpio_30_f = c2h_gpio_10_reg[30];
   assign c2h_gpio_10_gpio_29_f = c2h_gpio_10_reg[29];
   assign c2h_gpio_10_gpio_28_f = c2h_gpio_10_reg[28];
   assign c2h_gpio_10_gpio_27_f = c2h_gpio_10_reg[27];
   assign c2h_gpio_10_gpio_26_f = c2h_gpio_10_reg[26];
   assign c2h_gpio_10_gpio_25_f = c2h_gpio_10_reg[25];
   assign c2h_gpio_10_gpio_24_f = c2h_gpio_10_reg[24];
   assign c2h_gpio_10_gpio_23_f = c2h_gpio_10_reg[23];
   assign c2h_gpio_10_gpio_22_f = c2h_gpio_10_reg[22];
   assign c2h_gpio_10_gpio_21_f = c2h_gpio_10_reg[21];
   assign c2h_gpio_10_gpio_20_f = c2h_gpio_10_reg[20];
   assign c2h_gpio_10_gpio_19_f = c2h_gpio_10_reg[19];
   assign c2h_gpio_10_gpio_18_f = c2h_gpio_10_reg[18];
   assign c2h_gpio_10_gpio_17_f = c2h_gpio_10_reg[17];
   assign c2h_gpio_10_gpio_16_f = c2h_gpio_10_reg[16];
   assign c2h_gpio_10_gpio_15_f = c2h_gpio_10_reg[15];
   assign c2h_gpio_10_gpio_14_f = c2h_gpio_10_reg[14];
   assign c2h_gpio_10_gpio_13_f = c2h_gpio_10_reg[13];
   assign c2h_gpio_10_gpio_12_f = c2h_gpio_10_reg[12];
   assign c2h_gpio_10_gpio_11_f = c2h_gpio_10_reg[11];
   assign c2h_gpio_10_gpio_10_f = c2h_gpio_10_reg[10];
   assign c2h_gpio_10_gpio_9_f = c2h_gpio_10_reg[9];
   assign c2h_gpio_10_gpio_8_f = c2h_gpio_10_reg[8];
   assign c2h_gpio_10_gpio_7_f = c2h_gpio_10_reg[7];
   assign c2h_gpio_10_gpio_6_f = c2h_gpio_10_reg[6];
   assign c2h_gpio_10_gpio_5_f = c2h_gpio_10_reg[5];
   assign c2h_gpio_10_gpio_4_f = c2h_gpio_10_reg[4];
   assign c2h_gpio_10_gpio_3_f = c2h_gpio_10_reg[3];
   assign c2h_gpio_10_gpio_2_f = c2h_gpio_10_reg[2];
   assign c2h_gpio_10_gpio_1_f = c2h_gpio_10_reg[1];
   assign c2h_gpio_10_gpio_0_f = c2h_gpio_10_reg[0];
   assign c2h_gpio_11_gpio_31_f = c2h_gpio_11_reg[31];
   assign c2h_gpio_11_gpio_30_f = c2h_gpio_11_reg[30];
   assign c2h_gpio_11_gpio_29_f = c2h_gpio_11_reg[29];
   assign c2h_gpio_11_gpio_28_f = c2h_gpio_11_reg[28];
   assign c2h_gpio_11_gpio_27_f = c2h_gpio_11_reg[27];
   assign c2h_gpio_11_gpio_26_f = c2h_gpio_11_reg[26];
   assign c2h_gpio_11_gpio_25_f = c2h_gpio_11_reg[25];
   assign c2h_gpio_11_gpio_24_f = c2h_gpio_11_reg[24];
   assign c2h_gpio_11_gpio_23_f = c2h_gpio_11_reg[23];
   assign c2h_gpio_11_gpio_22_f = c2h_gpio_11_reg[22];
   assign c2h_gpio_11_gpio_21_f = c2h_gpio_11_reg[21];
   assign c2h_gpio_11_gpio_20_f = c2h_gpio_11_reg[20];
   assign c2h_gpio_11_gpio_19_f = c2h_gpio_11_reg[19];
   assign c2h_gpio_11_gpio_18_f = c2h_gpio_11_reg[18];
   assign c2h_gpio_11_gpio_17_f = c2h_gpio_11_reg[17];
   assign c2h_gpio_11_gpio_16_f = c2h_gpio_11_reg[16];
   assign c2h_gpio_11_gpio_15_f = c2h_gpio_11_reg[15];
   assign c2h_gpio_11_gpio_14_f = c2h_gpio_11_reg[14];
   assign c2h_gpio_11_gpio_13_f = c2h_gpio_11_reg[13];
   assign c2h_gpio_11_gpio_12_f = c2h_gpio_11_reg[12];
   assign c2h_gpio_11_gpio_11_f = c2h_gpio_11_reg[11];
   assign c2h_gpio_11_gpio_10_f = c2h_gpio_11_reg[10];
   assign c2h_gpio_11_gpio_9_f = c2h_gpio_11_reg[9];
   assign c2h_gpio_11_gpio_8_f = c2h_gpio_11_reg[8];
   assign c2h_gpio_11_gpio_7_f = c2h_gpio_11_reg[7];
   assign c2h_gpio_11_gpio_6_f = c2h_gpio_11_reg[6];
   assign c2h_gpio_11_gpio_5_f = c2h_gpio_11_reg[5];
   assign c2h_gpio_11_gpio_4_f = c2h_gpio_11_reg[4];
   assign c2h_gpio_11_gpio_3_f = c2h_gpio_11_reg[3];
   assign c2h_gpio_11_gpio_2_f = c2h_gpio_11_reg[2];
   assign c2h_gpio_11_gpio_1_f = c2h_gpio_11_reg[1];
   assign c2h_gpio_11_gpio_0_f = c2h_gpio_11_reg[0];
   assign c2h_gpio_12_gpio_31_f = c2h_gpio_12_reg[31];
   assign c2h_gpio_12_gpio_30_f = c2h_gpio_12_reg[30];
   assign c2h_gpio_12_gpio_29_f = c2h_gpio_12_reg[29];
   assign c2h_gpio_12_gpio_28_f = c2h_gpio_12_reg[28];
   assign c2h_gpio_12_gpio_27_f = c2h_gpio_12_reg[27];
   assign c2h_gpio_12_gpio_26_f = c2h_gpio_12_reg[26];
   assign c2h_gpio_12_gpio_25_f = c2h_gpio_12_reg[25];
   assign c2h_gpio_12_gpio_24_f = c2h_gpio_12_reg[24];
   assign c2h_gpio_12_gpio_23_f = c2h_gpio_12_reg[23];
   assign c2h_gpio_12_gpio_22_f = c2h_gpio_12_reg[22];
   assign c2h_gpio_12_gpio_21_f = c2h_gpio_12_reg[21];
   assign c2h_gpio_12_gpio_20_f = c2h_gpio_12_reg[20];
   assign c2h_gpio_12_gpio_19_f = c2h_gpio_12_reg[19];
   assign c2h_gpio_12_gpio_18_f = c2h_gpio_12_reg[18];
   assign c2h_gpio_12_gpio_17_f = c2h_gpio_12_reg[17];
   assign c2h_gpio_12_gpio_16_f = c2h_gpio_12_reg[16];
   assign c2h_gpio_12_gpio_15_f = c2h_gpio_12_reg[15];
   assign c2h_gpio_12_gpio_14_f = c2h_gpio_12_reg[14];
   assign c2h_gpio_12_gpio_13_f = c2h_gpio_12_reg[13];
   assign c2h_gpio_12_gpio_12_f = c2h_gpio_12_reg[12];
   assign c2h_gpio_12_gpio_11_f = c2h_gpio_12_reg[11];
   assign c2h_gpio_12_gpio_10_f = c2h_gpio_12_reg[10];
   assign c2h_gpio_12_gpio_9_f = c2h_gpio_12_reg[9];
   assign c2h_gpio_12_gpio_8_f = c2h_gpio_12_reg[8];
   assign c2h_gpio_12_gpio_7_f = c2h_gpio_12_reg[7];
   assign c2h_gpio_12_gpio_6_f = c2h_gpio_12_reg[6];
   assign c2h_gpio_12_gpio_5_f = c2h_gpio_12_reg[5];
   assign c2h_gpio_12_gpio_4_f = c2h_gpio_12_reg[4];
   assign c2h_gpio_12_gpio_3_f = c2h_gpio_12_reg[3];
   assign c2h_gpio_12_gpio_2_f = c2h_gpio_12_reg[2];
   assign c2h_gpio_12_gpio_1_f = c2h_gpio_12_reg[1];
   assign c2h_gpio_12_gpio_0_f = c2h_gpio_12_reg[0];
   assign c2h_gpio_13_gpio_31_f = c2h_gpio_13_reg[31];
   assign c2h_gpio_13_gpio_30_f = c2h_gpio_13_reg[30];
   assign c2h_gpio_13_gpio_29_f = c2h_gpio_13_reg[29];
   assign c2h_gpio_13_gpio_28_f = c2h_gpio_13_reg[28];
   assign c2h_gpio_13_gpio_27_f = c2h_gpio_13_reg[27];
   assign c2h_gpio_13_gpio_26_f = c2h_gpio_13_reg[26];
   assign c2h_gpio_13_gpio_25_f = c2h_gpio_13_reg[25];
   assign c2h_gpio_13_gpio_24_f = c2h_gpio_13_reg[24];
   assign c2h_gpio_13_gpio_23_f = c2h_gpio_13_reg[23];
   assign c2h_gpio_13_gpio_22_f = c2h_gpio_13_reg[22];
   assign c2h_gpio_13_gpio_21_f = c2h_gpio_13_reg[21];
   assign c2h_gpio_13_gpio_20_f = c2h_gpio_13_reg[20];
   assign c2h_gpio_13_gpio_19_f = c2h_gpio_13_reg[19];
   assign c2h_gpio_13_gpio_18_f = c2h_gpio_13_reg[18];
   assign c2h_gpio_13_gpio_17_f = c2h_gpio_13_reg[17];
   assign c2h_gpio_13_gpio_16_f = c2h_gpio_13_reg[16];
   assign c2h_gpio_13_gpio_15_f = c2h_gpio_13_reg[15];
   assign c2h_gpio_13_gpio_14_f = c2h_gpio_13_reg[14];
   assign c2h_gpio_13_gpio_13_f = c2h_gpio_13_reg[13];
   assign c2h_gpio_13_gpio_12_f = c2h_gpio_13_reg[12];
   assign c2h_gpio_13_gpio_11_f = c2h_gpio_13_reg[11];
   assign c2h_gpio_13_gpio_10_f = c2h_gpio_13_reg[10];
   assign c2h_gpio_13_gpio_9_f = c2h_gpio_13_reg[9];
   assign c2h_gpio_13_gpio_8_f = c2h_gpio_13_reg[8];
   assign c2h_gpio_13_gpio_7_f = c2h_gpio_13_reg[7];
   assign c2h_gpio_13_gpio_6_f = c2h_gpio_13_reg[6];
   assign c2h_gpio_13_gpio_5_f = c2h_gpio_13_reg[5];
   assign c2h_gpio_13_gpio_4_f = c2h_gpio_13_reg[4];
   assign c2h_gpio_13_gpio_3_f = c2h_gpio_13_reg[3];
   assign c2h_gpio_13_gpio_2_f = c2h_gpio_13_reg[2];
   assign c2h_gpio_13_gpio_1_f = c2h_gpio_13_reg[1];
   assign c2h_gpio_13_gpio_0_f = c2h_gpio_13_reg[0];
   assign c2h_gpio_14_gpio_31_f = c2h_gpio_14_reg[31];
   assign c2h_gpio_14_gpio_30_f = c2h_gpio_14_reg[30];
   assign c2h_gpio_14_gpio_29_f = c2h_gpio_14_reg[29];
   assign c2h_gpio_14_gpio_28_f = c2h_gpio_14_reg[28];
   assign c2h_gpio_14_gpio_27_f = c2h_gpio_14_reg[27];
   assign c2h_gpio_14_gpio_26_f = c2h_gpio_14_reg[26];
   assign c2h_gpio_14_gpio_25_f = c2h_gpio_14_reg[25];
   assign c2h_gpio_14_gpio_24_f = c2h_gpio_14_reg[24];
   assign c2h_gpio_14_gpio_23_f = c2h_gpio_14_reg[23];
   assign c2h_gpio_14_gpio_22_f = c2h_gpio_14_reg[22];
   assign c2h_gpio_14_gpio_21_f = c2h_gpio_14_reg[21];
   assign c2h_gpio_14_gpio_20_f = c2h_gpio_14_reg[20];
   assign c2h_gpio_14_gpio_19_f = c2h_gpio_14_reg[19];
   assign c2h_gpio_14_gpio_18_f = c2h_gpio_14_reg[18];
   assign c2h_gpio_14_gpio_17_f = c2h_gpio_14_reg[17];
   assign c2h_gpio_14_gpio_16_f = c2h_gpio_14_reg[16];
   assign c2h_gpio_14_gpio_15_f = c2h_gpio_14_reg[15];
   assign c2h_gpio_14_gpio_14_f = c2h_gpio_14_reg[14];
   assign c2h_gpio_14_gpio_13_f = c2h_gpio_14_reg[13];
   assign c2h_gpio_14_gpio_12_f = c2h_gpio_14_reg[12];
   assign c2h_gpio_14_gpio_11_f = c2h_gpio_14_reg[11];
   assign c2h_gpio_14_gpio_10_f = c2h_gpio_14_reg[10];
   assign c2h_gpio_14_gpio_9_f = c2h_gpio_14_reg[9];
   assign c2h_gpio_14_gpio_8_f = c2h_gpio_14_reg[8];
   assign c2h_gpio_14_gpio_7_f = c2h_gpio_14_reg[7];
   assign c2h_gpio_14_gpio_6_f = c2h_gpio_14_reg[6];
   assign c2h_gpio_14_gpio_5_f = c2h_gpio_14_reg[5];
   assign c2h_gpio_14_gpio_4_f = c2h_gpio_14_reg[4];
   assign c2h_gpio_14_gpio_3_f = c2h_gpio_14_reg[3];
   assign c2h_gpio_14_gpio_2_f = c2h_gpio_14_reg[2];
   assign c2h_gpio_14_gpio_1_f = c2h_gpio_14_reg[1];
   assign c2h_gpio_14_gpio_0_f = c2h_gpio_14_reg[0];
   assign c2h_gpio_15_gpio_31_f = c2h_gpio_15_reg[31];
   assign c2h_gpio_15_gpio_30_f = c2h_gpio_15_reg[30];
   assign c2h_gpio_15_gpio_29_f = c2h_gpio_15_reg[29];
   assign c2h_gpio_15_gpio_28_f = c2h_gpio_15_reg[28];
   assign c2h_gpio_15_gpio_27_f = c2h_gpio_15_reg[27];
   assign c2h_gpio_15_gpio_26_f = c2h_gpio_15_reg[26];
   assign c2h_gpio_15_gpio_25_f = c2h_gpio_15_reg[25];
   assign c2h_gpio_15_gpio_24_f = c2h_gpio_15_reg[24];
   assign c2h_gpio_15_gpio_23_f = c2h_gpio_15_reg[23];
   assign c2h_gpio_15_gpio_22_f = c2h_gpio_15_reg[22];
   assign c2h_gpio_15_gpio_21_f = c2h_gpio_15_reg[21];
   assign c2h_gpio_15_gpio_20_f = c2h_gpio_15_reg[20];
   assign c2h_gpio_15_gpio_19_f = c2h_gpio_15_reg[19];
   assign c2h_gpio_15_gpio_18_f = c2h_gpio_15_reg[18];
   assign c2h_gpio_15_gpio_17_f = c2h_gpio_15_reg[17];
   assign c2h_gpio_15_gpio_16_f = c2h_gpio_15_reg[16];
   assign c2h_gpio_15_gpio_15_f = c2h_gpio_15_reg[15];
   assign c2h_gpio_15_gpio_14_f = c2h_gpio_15_reg[14];
   assign c2h_gpio_15_gpio_13_f = c2h_gpio_15_reg[13];
   assign c2h_gpio_15_gpio_12_f = c2h_gpio_15_reg[12];
   assign c2h_gpio_15_gpio_11_f = c2h_gpio_15_reg[11];
   assign c2h_gpio_15_gpio_10_f = c2h_gpio_15_reg[10];
   assign c2h_gpio_15_gpio_9_f = c2h_gpio_15_reg[9];
   assign c2h_gpio_15_gpio_8_f = c2h_gpio_15_reg[8];
   assign c2h_gpio_15_gpio_7_f = c2h_gpio_15_reg[7];
   assign c2h_gpio_15_gpio_6_f = c2h_gpio_15_reg[6];
   assign c2h_gpio_15_gpio_5_f = c2h_gpio_15_reg[5];
   assign c2h_gpio_15_gpio_4_f = c2h_gpio_15_reg[4];
   assign c2h_gpio_15_gpio_3_f = c2h_gpio_15_reg[3];
   assign c2h_gpio_15_gpio_2_f = c2h_gpio_15_reg[2];
   assign c2h_gpio_15_gpio_1_f = c2h_gpio_15_reg[1];
   assign c2h_gpio_15_gpio_0_f = c2h_gpio_15_reg[0];
   assign h2c_gpio_0_gpio_31_f = h2c_gpio_0_reg[31];
   assign h2c_gpio_0_gpio_30_f = h2c_gpio_0_reg[30];
   assign h2c_gpio_0_gpio_29_f = h2c_gpio_0_reg[29];
   assign h2c_gpio_0_gpio_28_f = h2c_gpio_0_reg[28];
   assign h2c_gpio_0_gpio_27_f = h2c_gpio_0_reg[27];
   assign h2c_gpio_0_gpio_26_f = h2c_gpio_0_reg[26];
   assign h2c_gpio_0_gpio_25_f = h2c_gpio_0_reg[25];
   assign h2c_gpio_0_gpio_24_f = h2c_gpio_0_reg[24];
   assign h2c_gpio_0_gpio_23_f = h2c_gpio_0_reg[23];
   assign h2c_gpio_0_gpio_22_f = h2c_gpio_0_reg[22];
   assign h2c_gpio_0_gpio_21_f = h2c_gpio_0_reg[21];
   assign h2c_gpio_0_gpio_20_f = h2c_gpio_0_reg[20];
   assign h2c_gpio_0_gpio_19_f = h2c_gpio_0_reg[19];
   assign h2c_gpio_0_gpio_18_f = h2c_gpio_0_reg[18];
   assign h2c_gpio_0_gpio_17_f = h2c_gpio_0_reg[17];
   assign h2c_gpio_0_gpio_16_f = h2c_gpio_0_reg[16];
   assign h2c_gpio_0_gpio_15_f = h2c_gpio_0_reg[15];
   assign h2c_gpio_0_gpio_14_f = h2c_gpio_0_reg[14];
   assign h2c_gpio_0_gpio_13_f = h2c_gpio_0_reg[13];
   assign h2c_gpio_0_gpio_12_f = h2c_gpio_0_reg[12];
   assign h2c_gpio_0_gpio_11_f = h2c_gpio_0_reg[11];
   assign h2c_gpio_0_gpio_10_f = h2c_gpio_0_reg[10];
   assign h2c_gpio_0_gpio_9_f = h2c_gpio_0_reg[9];
   assign h2c_gpio_0_gpio_8_f = h2c_gpio_0_reg[8];
   assign h2c_gpio_0_gpio_7_f = h2c_gpio_0_reg[7];
   assign h2c_gpio_0_gpio_6_f = h2c_gpio_0_reg[6];
   assign h2c_gpio_0_gpio_5_f = h2c_gpio_0_reg[5];
   assign h2c_gpio_0_gpio_4_f = h2c_gpio_0_reg[4];
   assign h2c_gpio_0_gpio_3_f = h2c_gpio_0_reg[3];
   assign h2c_gpio_0_gpio_2_f = h2c_gpio_0_reg[2];
   assign h2c_gpio_0_gpio_1_f = h2c_gpio_0_reg[1];
   assign h2c_gpio_0_gpio_0_f = h2c_gpio_0_reg[0];
   assign h2c_gpio_1_gpio_31_f = h2c_gpio_1_reg[31];
   assign h2c_gpio_1_gpio_30_f = h2c_gpio_1_reg[30];
   assign h2c_gpio_1_gpio_29_f = h2c_gpio_1_reg[29];
   assign h2c_gpio_1_gpio_28_f = h2c_gpio_1_reg[28];
   assign h2c_gpio_1_gpio_27_f = h2c_gpio_1_reg[27];
   assign h2c_gpio_1_gpio_26_f = h2c_gpio_1_reg[26];
   assign h2c_gpio_1_gpio_25_f = h2c_gpio_1_reg[25];
   assign h2c_gpio_1_gpio_24_f = h2c_gpio_1_reg[24];
   assign h2c_gpio_1_gpio_23_f = h2c_gpio_1_reg[23];
   assign h2c_gpio_1_gpio_22_f = h2c_gpio_1_reg[22];
   assign h2c_gpio_1_gpio_21_f = h2c_gpio_1_reg[21];
   assign h2c_gpio_1_gpio_20_f = h2c_gpio_1_reg[20];
   assign h2c_gpio_1_gpio_19_f = h2c_gpio_1_reg[19];
   assign h2c_gpio_1_gpio_18_f = h2c_gpio_1_reg[18];
   assign h2c_gpio_1_gpio_17_f = h2c_gpio_1_reg[17];
   assign h2c_gpio_1_gpio_16_f = h2c_gpio_1_reg[16];
   assign h2c_gpio_1_gpio_15_f = h2c_gpio_1_reg[15];
   assign h2c_gpio_1_gpio_14_f = h2c_gpio_1_reg[14];
   assign h2c_gpio_1_gpio_13_f = h2c_gpio_1_reg[13];
   assign h2c_gpio_1_gpio_12_f = h2c_gpio_1_reg[12];
   assign h2c_gpio_1_gpio_11_f = h2c_gpio_1_reg[11];
   assign h2c_gpio_1_gpio_10_f = h2c_gpio_1_reg[10];
   assign h2c_gpio_1_gpio_9_f = h2c_gpio_1_reg[9];
   assign h2c_gpio_1_gpio_8_f = h2c_gpio_1_reg[8];
   assign h2c_gpio_1_gpio_7_f = h2c_gpio_1_reg[7];
   assign h2c_gpio_1_gpio_6_f = h2c_gpio_1_reg[6];
   assign h2c_gpio_1_gpio_5_f = h2c_gpio_1_reg[5];
   assign h2c_gpio_1_gpio_4_f = h2c_gpio_1_reg[4];
   assign h2c_gpio_1_gpio_3_f = h2c_gpio_1_reg[3];
   assign h2c_gpio_1_gpio_2_f = h2c_gpio_1_reg[2];
   assign h2c_gpio_1_gpio_1_f = h2c_gpio_1_reg[1];
   assign h2c_gpio_1_gpio_0_f = h2c_gpio_1_reg[0];
   assign h2c_gpio_2_gpio_31_f = h2c_gpio_2_reg[31];
   assign h2c_gpio_2_gpio_30_f = h2c_gpio_2_reg[30];
   assign h2c_gpio_2_gpio_29_f = h2c_gpio_2_reg[29];
   assign h2c_gpio_2_gpio_28_f = h2c_gpio_2_reg[28];
   assign h2c_gpio_2_gpio_27_f = h2c_gpio_2_reg[27];
   assign h2c_gpio_2_gpio_26_f = h2c_gpio_2_reg[26];
   assign h2c_gpio_2_gpio_25_f = h2c_gpio_2_reg[25];
   assign h2c_gpio_2_gpio_24_f = h2c_gpio_2_reg[24];
   assign h2c_gpio_2_gpio_23_f = h2c_gpio_2_reg[23];
   assign h2c_gpio_2_gpio_22_f = h2c_gpio_2_reg[22];
   assign h2c_gpio_2_gpio_21_f = h2c_gpio_2_reg[21];
   assign h2c_gpio_2_gpio_20_f = h2c_gpio_2_reg[20];
   assign h2c_gpio_2_gpio_19_f = h2c_gpio_2_reg[19];
   assign h2c_gpio_2_gpio_18_f = h2c_gpio_2_reg[18];
   assign h2c_gpio_2_gpio_17_f = h2c_gpio_2_reg[17];
   assign h2c_gpio_2_gpio_16_f = h2c_gpio_2_reg[16];
   assign h2c_gpio_2_gpio_15_f = h2c_gpio_2_reg[15];
   assign h2c_gpio_2_gpio_14_f = h2c_gpio_2_reg[14];
   assign h2c_gpio_2_gpio_13_f = h2c_gpio_2_reg[13];
   assign h2c_gpio_2_gpio_12_f = h2c_gpio_2_reg[12];
   assign h2c_gpio_2_gpio_11_f = h2c_gpio_2_reg[11];
   assign h2c_gpio_2_gpio_10_f = h2c_gpio_2_reg[10];
   assign h2c_gpio_2_gpio_9_f = h2c_gpio_2_reg[9];
   assign h2c_gpio_2_gpio_8_f = h2c_gpio_2_reg[8];
   assign h2c_gpio_2_gpio_7_f = h2c_gpio_2_reg[7];
   assign h2c_gpio_2_gpio_6_f = h2c_gpio_2_reg[6];
   assign h2c_gpio_2_gpio_5_f = h2c_gpio_2_reg[5];
   assign h2c_gpio_2_gpio_4_f = h2c_gpio_2_reg[4];
   assign h2c_gpio_2_gpio_3_f = h2c_gpio_2_reg[3];
   assign h2c_gpio_2_gpio_2_f = h2c_gpio_2_reg[2];
   assign h2c_gpio_2_gpio_1_f = h2c_gpio_2_reg[1];
   assign h2c_gpio_2_gpio_0_f = h2c_gpio_2_reg[0];
   assign h2c_gpio_3_gpio_31_f = h2c_gpio_3_reg[31];
   assign h2c_gpio_3_gpio_30_f = h2c_gpio_3_reg[30];
   assign h2c_gpio_3_gpio_29_f = h2c_gpio_3_reg[29];
   assign h2c_gpio_3_gpio_28_f = h2c_gpio_3_reg[28];
   assign h2c_gpio_3_gpio_27_f = h2c_gpio_3_reg[27];
   assign h2c_gpio_3_gpio_26_f = h2c_gpio_3_reg[26];
   assign h2c_gpio_3_gpio_25_f = h2c_gpio_3_reg[25];
   assign h2c_gpio_3_gpio_24_f = h2c_gpio_3_reg[24];
   assign h2c_gpio_3_gpio_23_f = h2c_gpio_3_reg[23];
   assign h2c_gpio_3_gpio_22_f = h2c_gpio_3_reg[22];
   assign h2c_gpio_3_gpio_21_f = h2c_gpio_3_reg[21];
   assign h2c_gpio_3_gpio_20_f = h2c_gpio_3_reg[20];
   assign h2c_gpio_3_gpio_19_f = h2c_gpio_3_reg[19];
   assign h2c_gpio_3_gpio_18_f = h2c_gpio_3_reg[18];
   assign h2c_gpio_3_gpio_17_f = h2c_gpio_3_reg[17];
   assign h2c_gpio_3_gpio_16_f = h2c_gpio_3_reg[16];
   assign h2c_gpio_3_gpio_15_f = h2c_gpio_3_reg[15];
   assign h2c_gpio_3_gpio_14_f = h2c_gpio_3_reg[14];
   assign h2c_gpio_3_gpio_13_f = h2c_gpio_3_reg[13];
   assign h2c_gpio_3_gpio_12_f = h2c_gpio_3_reg[12];
   assign h2c_gpio_3_gpio_11_f = h2c_gpio_3_reg[11];
   assign h2c_gpio_3_gpio_10_f = h2c_gpio_3_reg[10];
   assign h2c_gpio_3_gpio_9_f = h2c_gpio_3_reg[9];
   assign h2c_gpio_3_gpio_8_f = h2c_gpio_3_reg[8];
   assign h2c_gpio_3_gpio_7_f = h2c_gpio_3_reg[7];
   assign h2c_gpio_3_gpio_6_f = h2c_gpio_3_reg[6];
   assign h2c_gpio_3_gpio_5_f = h2c_gpio_3_reg[5];
   assign h2c_gpio_3_gpio_4_f = h2c_gpio_3_reg[4];
   assign h2c_gpio_3_gpio_3_f = h2c_gpio_3_reg[3];
   assign h2c_gpio_3_gpio_2_f = h2c_gpio_3_reg[2];
   assign h2c_gpio_3_gpio_1_f = h2c_gpio_3_reg[1];
   assign h2c_gpio_3_gpio_0_f = h2c_gpio_3_reg[0];
   assign h2c_gpio_4_gpio_31_f = h2c_gpio_4_reg[31];
   assign h2c_gpio_4_gpio_30_f = h2c_gpio_4_reg[30];
   assign h2c_gpio_4_gpio_29_f = h2c_gpio_4_reg[29];
   assign h2c_gpio_4_gpio_28_f = h2c_gpio_4_reg[28];
   assign h2c_gpio_4_gpio_27_f = h2c_gpio_4_reg[27];
   assign h2c_gpio_4_gpio_26_f = h2c_gpio_4_reg[26];
   assign h2c_gpio_4_gpio_25_f = h2c_gpio_4_reg[25];
   assign h2c_gpio_4_gpio_24_f = h2c_gpio_4_reg[24];
   assign h2c_gpio_4_gpio_23_f = h2c_gpio_4_reg[23];
   assign h2c_gpio_4_gpio_22_f = h2c_gpio_4_reg[22];
   assign h2c_gpio_4_gpio_21_f = h2c_gpio_4_reg[21];
   assign h2c_gpio_4_gpio_20_f = h2c_gpio_4_reg[20];
   assign h2c_gpio_4_gpio_19_f = h2c_gpio_4_reg[19];
   assign h2c_gpio_4_gpio_18_f = h2c_gpio_4_reg[18];
   assign h2c_gpio_4_gpio_17_f = h2c_gpio_4_reg[17];
   assign h2c_gpio_4_gpio_16_f = h2c_gpio_4_reg[16];
   assign h2c_gpio_4_gpio_15_f = h2c_gpio_4_reg[15];
   assign h2c_gpio_4_gpio_14_f = h2c_gpio_4_reg[14];
   assign h2c_gpio_4_gpio_13_f = h2c_gpio_4_reg[13];
   assign h2c_gpio_4_gpio_12_f = h2c_gpio_4_reg[12];
   assign h2c_gpio_4_gpio_11_f = h2c_gpio_4_reg[11];
   assign h2c_gpio_4_gpio_10_f = h2c_gpio_4_reg[10];
   assign h2c_gpio_4_gpio_9_f = h2c_gpio_4_reg[9];
   assign h2c_gpio_4_gpio_8_f = h2c_gpio_4_reg[8];
   assign h2c_gpio_4_gpio_7_f = h2c_gpio_4_reg[7];
   assign h2c_gpio_4_gpio_6_f = h2c_gpio_4_reg[6];
   assign h2c_gpio_4_gpio_5_f = h2c_gpio_4_reg[5];
   assign h2c_gpio_4_gpio_4_f = h2c_gpio_4_reg[4];
   assign h2c_gpio_4_gpio_3_f = h2c_gpio_4_reg[3];
   assign h2c_gpio_4_gpio_2_f = h2c_gpio_4_reg[2];
   assign h2c_gpio_4_gpio_1_f = h2c_gpio_4_reg[1];
   assign h2c_gpio_4_gpio_0_f = h2c_gpio_4_reg[0];
   assign h2c_gpio_5_gpio_31_f = h2c_gpio_5_reg[31];
   assign h2c_gpio_5_gpio_30_f = h2c_gpio_5_reg[30];
   assign h2c_gpio_5_gpio_29_f = h2c_gpio_5_reg[29];
   assign h2c_gpio_5_gpio_28_f = h2c_gpio_5_reg[28];
   assign h2c_gpio_5_gpio_27_f = h2c_gpio_5_reg[27];
   assign h2c_gpio_5_gpio_26_f = h2c_gpio_5_reg[26];
   assign h2c_gpio_5_gpio_25_f = h2c_gpio_5_reg[25];
   assign h2c_gpio_5_gpio_24_f = h2c_gpio_5_reg[24];
   assign h2c_gpio_5_gpio_23_f = h2c_gpio_5_reg[23];
   assign h2c_gpio_5_gpio_22_f = h2c_gpio_5_reg[22];
   assign h2c_gpio_5_gpio_21_f = h2c_gpio_5_reg[21];
   assign h2c_gpio_5_gpio_20_f = h2c_gpio_5_reg[20];
   assign h2c_gpio_5_gpio_19_f = h2c_gpio_5_reg[19];
   assign h2c_gpio_5_gpio_18_f = h2c_gpio_5_reg[18];
   assign h2c_gpio_5_gpio_17_f = h2c_gpio_5_reg[17];
   assign h2c_gpio_5_gpio_16_f = h2c_gpio_5_reg[16];
   assign h2c_gpio_5_gpio_15_f = h2c_gpio_5_reg[15];
   assign h2c_gpio_5_gpio_14_f = h2c_gpio_5_reg[14];
   assign h2c_gpio_5_gpio_13_f = h2c_gpio_5_reg[13];
   assign h2c_gpio_5_gpio_12_f = h2c_gpio_5_reg[12];
   assign h2c_gpio_5_gpio_11_f = h2c_gpio_5_reg[11];
   assign h2c_gpio_5_gpio_10_f = h2c_gpio_5_reg[10];
   assign h2c_gpio_5_gpio_9_f = h2c_gpio_5_reg[9];
   assign h2c_gpio_5_gpio_8_f = h2c_gpio_5_reg[8];
   assign h2c_gpio_5_gpio_7_f = h2c_gpio_5_reg[7];
   assign h2c_gpio_5_gpio_6_f = h2c_gpio_5_reg[6];
   assign h2c_gpio_5_gpio_5_f = h2c_gpio_5_reg[5];
   assign h2c_gpio_5_gpio_4_f = h2c_gpio_5_reg[4];
   assign h2c_gpio_5_gpio_3_f = h2c_gpio_5_reg[3];
   assign h2c_gpio_5_gpio_2_f = h2c_gpio_5_reg[2];
   assign h2c_gpio_5_gpio_1_f = h2c_gpio_5_reg[1];
   assign h2c_gpio_5_gpio_0_f = h2c_gpio_5_reg[0];
   assign h2c_gpio_6_gpio_31_f = h2c_gpio_6_reg[31];
   assign h2c_gpio_6_gpio_30_f = h2c_gpio_6_reg[30];
   assign h2c_gpio_6_gpio_29_f = h2c_gpio_6_reg[29];
   assign h2c_gpio_6_gpio_28_f = h2c_gpio_6_reg[28];
   assign h2c_gpio_6_gpio_27_f = h2c_gpio_6_reg[27];
   assign h2c_gpio_6_gpio_26_f = h2c_gpio_6_reg[26];
   assign h2c_gpio_6_gpio_25_f = h2c_gpio_6_reg[25];
   assign h2c_gpio_6_gpio_24_f = h2c_gpio_6_reg[24];
   assign h2c_gpio_6_gpio_23_f = h2c_gpio_6_reg[23];
   assign h2c_gpio_6_gpio_22_f = h2c_gpio_6_reg[22];
   assign h2c_gpio_6_gpio_21_f = h2c_gpio_6_reg[21];
   assign h2c_gpio_6_gpio_20_f = h2c_gpio_6_reg[20];
   assign h2c_gpio_6_gpio_19_f = h2c_gpio_6_reg[19];
   assign h2c_gpio_6_gpio_18_f = h2c_gpio_6_reg[18];
   assign h2c_gpio_6_gpio_17_f = h2c_gpio_6_reg[17];
   assign h2c_gpio_6_gpio_16_f = h2c_gpio_6_reg[16];
   assign h2c_gpio_6_gpio_15_f = h2c_gpio_6_reg[15];
   assign h2c_gpio_6_gpio_14_f = h2c_gpio_6_reg[14];
   assign h2c_gpio_6_gpio_13_f = h2c_gpio_6_reg[13];
   assign h2c_gpio_6_gpio_12_f = h2c_gpio_6_reg[12];
   assign h2c_gpio_6_gpio_11_f = h2c_gpio_6_reg[11];
   assign h2c_gpio_6_gpio_10_f = h2c_gpio_6_reg[10];
   assign h2c_gpio_6_gpio_9_f = h2c_gpio_6_reg[9];
   assign h2c_gpio_6_gpio_8_f = h2c_gpio_6_reg[8];
   assign h2c_gpio_6_gpio_7_f = h2c_gpio_6_reg[7];
   assign h2c_gpio_6_gpio_6_f = h2c_gpio_6_reg[6];
   assign h2c_gpio_6_gpio_5_f = h2c_gpio_6_reg[5];
   assign h2c_gpio_6_gpio_4_f = h2c_gpio_6_reg[4];
   assign h2c_gpio_6_gpio_3_f = h2c_gpio_6_reg[3];
   assign h2c_gpio_6_gpio_2_f = h2c_gpio_6_reg[2];
   assign h2c_gpio_6_gpio_1_f = h2c_gpio_6_reg[1];
   assign h2c_gpio_6_gpio_0_f = h2c_gpio_6_reg[0];
   assign h2c_gpio_7_gpio_31_f = h2c_gpio_7_reg[31];
   assign h2c_gpio_7_gpio_30_f = h2c_gpio_7_reg[30];
   assign h2c_gpio_7_gpio_29_f = h2c_gpio_7_reg[29];
   assign h2c_gpio_7_gpio_28_f = h2c_gpio_7_reg[28];
   assign h2c_gpio_7_gpio_27_f = h2c_gpio_7_reg[27];
   assign h2c_gpio_7_gpio_26_f = h2c_gpio_7_reg[26];
   assign h2c_gpio_7_gpio_25_f = h2c_gpio_7_reg[25];
   assign h2c_gpio_7_gpio_24_f = h2c_gpio_7_reg[24];
   assign h2c_gpio_7_gpio_23_f = h2c_gpio_7_reg[23];
   assign h2c_gpio_7_gpio_22_f = h2c_gpio_7_reg[22];
   assign h2c_gpio_7_gpio_21_f = h2c_gpio_7_reg[21];
   assign h2c_gpio_7_gpio_20_f = h2c_gpio_7_reg[20];
   assign h2c_gpio_7_gpio_19_f = h2c_gpio_7_reg[19];
   assign h2c_gpio_7_gpio_18_f = h2c_gpio_7_reg[18];
   assign h2c_gpio_7_gpio_17_f = h2c_gpio_7_reg[17];
   assign h2c_gpio_7_gpio_16_f = h2c_gpio_7_reg[16];
   assign h2c_gpio_7_gpio_15_f = h2c_gpio_7_reg[15];
   assign h2c_gpio_7_gpio_14_f = h2c_gpio_7_reg[14];
   assign h2c_gpio_7_gpio_13_f = h2c_gpio_7_reg[13];
   assign h2c_gpio_7_gpio_12_f = h2c_gpio_7_reg[12];
   assign h2c_gpio_7_gpio_11_f = h2c_gpio_7_reg[11];
   assign h2c_gpio_7_gpio_10_f = h2c_gpio_7_reg[10];
   assign h2c_gpio_7_gpio_9_f = h2c_gpio_7_reg[9];
   assign h2c_gpio_7_gpio_8_f = h2c_gpio_7_reg[8];
   assign h2c_gpio_7_gpio_7_f = h2c_gpio_7_reg[7];
   assign h2c_gpio_7_gpio_6_f = h2c_gpio_7_reg[6];
   assign h2c_gpio_7_gpio_5_f = h2c_gpio_7_reg[5];
   assign h2c_gpio_7_gpio_4_f = h2c_gpio_7_reg[4];
   assign h2c_gpio_7_gpio_3_f = h2c_gpio_7_reg[3];
   assign h2c_gpio_7_gpio_2_f = h2c_gpio_7_reg[2];
   assign h2c_gpio_7_gpio_1_f = h2c_gpio_7_reg[1];
   assign h2c_gpio_7_gpio_0_f = h2c_gpio_7_reg[0];
   assign h2c_gpio_8_gpio_31_f = h2c_gpio_8_reg[31];
   assign h2c_gpio_8_gpio_30_f = h2c_gpio_8_reg[30];
   assign h2c_gpio_8_gpio_29_f = h2c_gpio_8_reg[29];
   assign h2c_gpio_8_gpio_28_f = h2c_gpio_8_reg[28];
   assign h2c_gpio_8_gpio_27_f = h2c_gpio_8_reg[27];
   assign h2c_gpio_8_gpio_26_f = h2c_gpio_8_reg[26];
   assign h2c_gpio_8_gpio_25_f = h2c_gpio_8_reg[25];
   assign h2c_gpio_8_gpio_24_f = h2c_gpio_8_reg[24];
   assign h2c_gpio_8_gpio_23_f = h2c_gpio_8_reg[23];
   assign h2c_gpio_8_gpio_22_f = h2c_gpio_8_reg[22];
   assign h2c_gpio_8_gpio_21_f = h2c_gpio_8_reg[21];
   assign h2c_gpio_8_gpio_20_f = h2c_gpio_8_reg[20];
   assign h2c_gpio_8_gpio_19_f = h2c_gpio_8_reg[19];
   assign h2c_gpio_8_gpio_18_f = h2c_gpio_8_reg[18];
   assign h2c_gpio_8_gpio_17_f = h2c_gpio_8_reg[17];
   assign h2c_gpio_8_gpio_16_f = h2c_gpio_8_reg[16];
   assign h2c_gpio_8_gpio_15_f = h2c_gpio_8_reg[15];
   assign h2c_gpio_8_gpio_14_f = h2c_gpio_8_reg[14];
   assign h2c_gpio_8_gpio_13_f = h2c_gpio_8_reg[13];
   assign h2c_gpio_8_gpio_12_f = h2c_gpio_8_reg[12];
   assign h2c_gpio_8_gpio_11_f = h2c_gpio_8_reg[11];
   assign h2c_gpio_8_gpio_10_f = h2c_gpio_8_reg[10];
   assign h2c_gpio_8_gpio_9_f = h2c_gpio_8_reg[9];
   assign h2c_gpio_8_gpio_8_f = h2c_gpio_8_reg[8];
   assign h2c_gpio_8_gpio_7_f = h2c_gpio_8_reg[7];
   assign h2c_gpio_8_gpio_6_f = h2c_gpio_8_reg[6];
   assign h2c_gpio_8_gpio_5_f = h2c_gpio_8_reg[5];
   assign h2c_gpio_8_gpio_4_f = h2c_gpio_8_reg[4];
   assign h2c_gpio_8_gpio_3_f = h2c_gpio_8_reg[3];
   assign h2c_gpio_8_gpio_2_f = h2c_gpio_8_reg[2];
   assign h2c_gpio_8_gpio_1_f = h2c_gpio_8_reg[1];
   assign h2c_gpio_8_gpio_0_f = h2c_gpio_8_reg[0];
   assign h2c_gpio_9_gpio_31_f = h2c_gpio_9_reg[31];
   assign h2c_gpio_9_gpio_30_f = h2c_gpio_9_reg[30];
   assign h2c_gpio_9_gpio_29_f = h2c_gpio_9_reg[29];
   assign h2c_gpio_9_gpio_28_f = h2c_gpio_9_reg[28];
   assign h2c_gpio_9_gpio_27_f = h2c_gpio_9_reg[27];
   assign h2c_gpio_9_gpio_26_f = h2c_gpio_9_reg[26];
   assign h2c_gpio_9_gpio_25_f = h2c_gpio_9_reg[25];
   assign h2c_gpio_9_gpio_24_f = h2c_gpio_9_reg[24];
   assign h2c_gpio_9_gpio_23_f = h2c_gpio_9_reg[23];
   assign h2c_gpio_9_gpio_22_f = h2c_gpio_9_reg[22];
   assign h2c_gpio_9_gpio_21_f = h2c_gpio_9_reg[21];
   assign h2c_gpio_9_gpio_20_f = h2c_gpio_9_reg[20];
   assign h2c_gpio_9_gpio_19_f = h2c_gpio_9_reg[19];
   assign h2c_gpio_9_gpio_18_f = h2c_gpio_9_reg[18];
   assign h2c_gpio_9_gpio_17_f = h2c_gpio_9_reg[17];
   assign h2c_gpio_9_gpio_16_f = h2c_gpio_9_reg[16];
   assign h2c_gpio_9_gpio_15_f = h2c_gpio_9_reg[15];
   assign h2c_gpio_9_gpio_14_f = h2c_gpio_9_reg[14];
   assign h2c_gpio_9_gpio_13_f = h2c_gpio_9_reg[13];
   assign h2c_gpio_9_gpio_12_f = h2c_gpio_9_reg[12];
   assign h2c_gpio_9_gpio_11_f = h2c_gpio_9_reg[11];
   assign h2c_gpio_9_gpio_10_f = h2c_gpio_9_reg[10];
   assign h2c_gpio_9_gpio_9_f = h2c_gpio_9_reg[9];
   assign h2c_gpio_9_gpio_8_f = h2c_gpio_9_reg[8];
   assign h2c_gpio_9_gpio_7_f = h2c_gpio_9_reg[7];
   assign h2c_gpio_9_gpio_6_f = h2c_gpio_9_reg[6];
   assign h2c_gpio_9_gpio_5_f = h2c_gpio_9_reg[5];
   assign h2c_gpio_9_gpio_4_f = h2c_gpio_9_reg[4];
   assign h2c_gpio_9_gpio_3_f = h2c_gpio_9_reg[3];
   assign h2c_gpio_9_gpio_2_f = h2c_gpio_9_reg[2];
   assign h2c_gpio_9_gpio_1_f = h2c_gpio_9_reg[1];
   assign h2c_gpio_9_gpio_0_f = h2c_gpio_9_reg[0];
   assign h2c_gpio_10_gpio_31_f = h2c_gpio_10_reg[31];
   assign h2c_gpio_10_gpio_30_f = h2c_gpio_10_reg[30];
   assign h2c_gpio_10_gpio_29_f = h2c_gpio_10_reg[29];
   assign h2c_gpio_10_gpio_28_f = h2c_gpio_10_reg[28];
   assign h2c_gpio_10_gpio_27_f = h2c_gpio_10_reg[27];
   assign h2c_gpio_10_gpio_26_f = h2c_gpio_10_reg[26];
   assign h2c_gpio_10_gpio_25_f = h2c_gpio_10_reg[25];
   assign h2c_gpio_10_gpio_24_f = h2c_gpio_10_reg[24];
   assign h2c_gpio_10_gpio_23_f = h2c_gpio_10_reg[23];
   assign h2c_gpio_10_gpio_22_f = h2c_gpio_10_reg[22];
   assign h2c_gpio_10_gpio_21_f = h2c_gpio_10_reg[21];
   assign h2c_gpio_10_gpio_20_f = h2c_gpio_10_reg[20];
   assign h2c_gpio_10_gpio_19_f = h2c_gpio_10_reg[19];
   assign h2c_gpio_10_gpio_18_f = h2c_gpio_10_reg[18];
   assign h2c_gpio_10_gpio_17_f = h2c_gpio_10_reg[17];
   assign h2c_gpio_10_gpio_16_f = h2c_gpio_10_reg[16];
   assign h2c_gpio_10_gpio_15_f = h2c_gpio_10_reg[15];
   assign h2c_gpio_10_gpio_14_f = h2c_gpio_10_reg[14];
   assign h2c_gpio_10_gpio_13_f = h2c_gpio_10_reg[13];
   assign h2c_gpio_10_gpio_12_f = h2c_gpio_10_reg[12];
   assign h2c_gpio_10_gpio_11_f = h2c_gpio_10_reg[11];
   assign h2c_gpio_10_gpio_10_f = h2c_gpio_10_reg[10];
   assign h2c_gpio_10_gpio_9_f = h2c_gpio_10_reg[9];
   assign h2c_gpio_10_gpio_8_f = h2c_gpio_10_reg[8];
   assign h2c_gpio_10_gpio_7_f = h2c_gpio_10_reg[7];
   assign h2c_gpio_10_gpio_6_f = h2c_gpio_10_reg[6];
   assign h2c_gpio_10_gpio_5_f = h2c_gpio_10_reg[5];
   assign h2c_gpio_10_gpio_4_f = h2c_gpio_10_reg[4];
   assign h2c_gpio_10_gpio_3_f = h2c_gpio_10_reg[3];
   assign h2c_gpio_10_gpio_2_f = h2c_gpio_10_reg[2];
   assign h2c_gpio_10_gpio_1_f = h2c_gpio_10_reg[1];
   assign h2c_gpio_10_gpio_0_f = h2c_gpio_10_reg[0];
   assign h2c_gpio_11_gpio_31_f = h2c_gpio_11_reg[31];
   assign h2c_gpio_11_gpio_30_f = h2c_gpio_11_reg[30];
   assign h2c_gpio_11_gpio_29_f = h2c_gpio_11_reg[29];
   assign h2c_gpio_11_gpio_28_f = h2c_gpio_11_reg[28];
   assign h2c_gpio_11_gpio_27_f = h2c_gpio_11_reg[27];
   assign h2c_gpio_11_gpio_26_f = h2c_gpio_11_reg[26];
   assign h2c_gpio_11_gpio_25_f = h2c_gpio_11_reg[25];
   assign h2c_gpio_11_gpio_24_f = h2c_gpio_11_reg[24];
   assign h2c_gpio_11_gpio_23_f = h2c_gpio_11_reg[23];
   assign h2c_gpio_11_gpio_22_f = h2c_gpio_11_reg[22];
   assign h2c_gpio_11_gpio_21_f = h2c_gpio_11_reg[21];
   assign h2c_gpio_11_gpio_20_f = h2c_gpio_11_reg[20];
   assign h2c_gpio_11_gpio_19_f = h2c_gpio_11_reg[19];
   assign h2c_gpio_11_gpio_18_f = h2c_gpio_11_reg[18];
   assign h2c_gpio_11_gpio_17_f = h2c_gpio_11_reg[17];
   assign h2c_gpio_11_gpio_16_f = h2c_gpio_11_reg[16];
   assign h2c_gpio_11_gpio_15_f = h2c_gpio_11_reg[15];
   assign h2c_gpio_11_gpio_14_f = h2c_gpio_11_reg[14];
   assign h2c_gpio_11_gpio_13_f = h2c_gpio_11_reg[13];
   assign h2c_gpio_11_gpio_12_f = h2c_gpio_11_reg[12];
   assign h2c_gpio_11_gpio_11_f = h2c_gpio_11_reg[11];
   assign h2c_gpio_11_gpio_10_f = h2c_gpio_11_reg[10];
   assign h2c_gpio_11_gpio_9_f = h2c_gpio_11_reg[9];
   assign h2c_gpio_11_gpio_8_f = h2c_gpio_11_reg[8];
   assign h2c_gpio_11_gpio_7_f = h2c_gpio_11_reg[7];
   assign h2c_gpio_11_gpio_6_f = h2c_gpio_11_reg[6];
   assign h2c_gpio_11_gpio_5_f = h2c_gpio_11_reg[5];
   assign h2c_gpio_11_gpio_4_f = h2c_gpio_11_reg[4];
   assign h2c_gpio_11_gpio_3_f = h2c_gpio_11_reg[3];
   assign h2c_gpio_11_gpio_2_f = h2c_gpio_11_reg[2];
   assign h2c_gpio_11_gpio_1_f = h2c_gpio_11_reg[1];
   assign h2c_gpio_11_gpio_0_f = h2c_gpio_11_reg[0];
   assign h2c_gpio_12_gpio_31_f = h2c_gpio_12_reg[31];
   assign h2c_gpio_12_gpio_30_f = h2c_gpio_12_reg[30];
   assign h2c_gpio_12_gpio_29_f = h2c_gpio_12_reg[29];
   assign h2c_gpio_12_gpio_28_f = h2c_gpio_12_reg[28];
   assign h2c_gpio_12_gpio_27_f = h2c_gpio_12_reg[27];
   assign h2c_gpio_12_gpio_26_f = h2c_gpio_12_reg[26];
   assign h2c_gpio_12_gpio_25_f = h2c_gpio_12_reg[25];
   assign h2c_gpio_12_gpio_24_f = h2c_gpio_12_reg[24];
   assign h2c_gpio_12_gpio_23_f = h2c_gpio_12_reg[23];
   assign h2c_gpio_12_gpio_22_f = h2c_gpio_12_reg[22];
   assign h2c_gpio_12_gpio_21_f = h2c_gpio_12_reg[21];
   assign h2c_gpio_12_gpio_20_f = h2c_gpio_12_reg[20];
   assign h2c_gpio_12_gpio_19_f = h2c_gpio_12_reg[19];
   assign h2c_gpio_12_gpio_18_f = h2c_gpio_12_reg[18];
   assign h2c_gpio_12_gpio_17_f = h2c_gpio_12_reg[17];
   assign h2c_gpio_12_gpio_16_f = h2c_gpio_12_reg[16];
   assign h2c_gpio_12_gpio_15_f = h2c_gpio_12_reg[15];
   assign h2c_gpio_12_gpio_14_f = h2c_gpio_12_reg[14];
   assign h2c_gpio_12_gpio_13_f = h2c_gpio_12_reg[13];
   assign h2c_gpio_12_gpio_12_f = h2c_gpio_12_reg[12];
   assign h2c_gpio_12_gpio_11_f = h2c_gpio_12_reg[11];
   assign h2c_gpio_12_gpio_10_f = h2c_gpio_12_reg[10];
   assign h2c_gpio_12_gpio_9_f = h2c_gpio_12_reg[9];
   assign h2c_gpio_12_gpio_8_f = h2c_gpio_12_reg[8];
   assign h2c_gpio_12_gpio_7_f = h2c_gpio_12_reg[7];
   assign h2c_gpio_12_gpio_6_f = h2c_gpio_12_reg[6];
   assign h2c_gpio_12_gpio_5_f = h2c_gpio_12_reg[5];
   assign h2c_gpio_12_gpio_4_f = h2c_gpio_12_reg[4];
   assign h2c_gpio_12_gpio_3_f = h2c_gpio_12_reg[3];
   assign h2c_gpio_12_gpio_2_f = h2c_gpio_12_reg[2];
   assign h2c_gpio_12_gpio_1_f = h2c_gpio_12_reg[1];
   assign h2c_gpio_12_gpio_0_f = h2c_gpio_12_reg[0];
   assign h2c_gpio_13_gpio_31_f = h2c_gpio_13_reg[31];
   assign h2c_gpio_13_gpio_30_f = h2c_gpio_13_reg[30];
   assign h2c_gpio_13_gpio_29_f = h2c_gpio_13_reg[29];
   assign h2c_gpio_13_gpio_28_f = h2c_gpio_13_reg[28];
   assign h2c_gpio_13_gpio_27_f = h2c_gpio_13_reg[27];
   assign h2c_gpio_13_gpio_26_f = h2c_gpio_13_reg[26];
   assign h2c_gpio_13_gpio_25_f = h2c_gpio_13_reg[25];
   assign h2c_gpio_13_gpio_24_f = h2c_gpio_13_reg[24];
   assign h2c_gpio_13_gpio_23_f = h2c_gpio_13_reg[23];
   assign h2c_gpio_13_gpio_22_f = h2c_gpio_13_reg[22];
   assign h2c_gpio_13_gpio_21_f = h2c_gpio_13_reg[21];
   assign h2c_gpio_13_gpio_20_f = h2c_gpio_13_reg[20];
   assign h2c_gpio_13_gpio_19_f = h2c_gpio_13_reg[19];
   assign h2c_gpio_13_gpio_18_f = h2c_gpio_13_reg[18];
   assign h2c_gpio_13_gpio_17_f = h2c_gpio_13_reg[17];
   assign h2c_gpio_13_gpio_16_f = h2c_gpio_13_reg[16];
   assign h2c_gpio_13_gpio_15_f = h2c_gpio_13_reg[15];
   assign h2c_gpio_13_gpio_14_f = h2c_gpio_13_reg[14];
   assign h2c_gpio_13_gpio_13_f = h2c_gpio_13_reg[13];
   assign h2c_gpio_13_gpio_12_f = h2c_gpio_13_reg[12];
   assign h2c_gpio_13_gpio_11_f = h2c_gpio_13_reg[11];
   assign h2c_gpio_13_gpio_10_f = h2c_gpio_13_reg[10];
   assign h2c_gpio_13_gpio_9_f = h2c_gpio_13_reg[9];
   assign h2c_gpio_13_gpio_8_f = h2c_gpio_13_reg[8];
   assign h2c_gpio_13_gpio_7_f = h2c_gpio_13_reg[7];
   assign h2c_gpio_13_gpio_6_f = h2c_gpio_13_reg[6];
   assign h2c_gpio_13_gpio_5_f = h2c_gpio_13_reg[5];
   assign h2c_gpio_13_gpio_4_f = h2c_gpio_13_reg[4];
   assign h2c_gpio_13_gpio_3_f = h2c_gpio_13_reg[3];
   assign h2c_gpio_13_gpio_2_f = h2c_gpio_13_reg[2];
   assign h2c_gpio_13_gpio_1_f = h2c_gpio_13_reg[1];
   assign h2c_gpio_13_gpio_0_f = h2c_gpio_13_reg[0];
   assign h2c_gpio_14_gpio_31_f = h2c_gpio_14_reg[31];
   assign h2c_gpio_14_gpio_30_f = h2c_gpio_14_reg[30];
   assign h2c_gpio_14_gpio_29_f = h2c_gpio_14_reg[29];
   assign h2c_gpio_14_gpio_28_f = h2c_gpio_14_reg[28];
   assign h2c_gpio_14_gpio_27_f = h2c_gpio_14_reg[27];
   assign h2c_gpio_14_gpio_26_f = h2c_gpio_14_reg[26];
   assign h2c_gpio_14_gpio_25_f = h2c_gpio_14_reg[25];
   assign h2c_gpio_14_gpio_24_f = h2c_gpio_14_reg[24];
   assign h2c_gpio_14_gpio_23_f = h2c_gpio_14_reg[23];
   assign h2c_gpio_14_gpio_22_f = h2c_gpio_14_reg[22];
   assign h2c_gpio_14_gpio_21_f = h2c_gpio_14_reg[21];
   assign h2c_gpio_14_gpio_20_f = h2c_gpio_14_reg[20];
   assign h2c_gpio_14_gpio_19_f = h2c_gpio_14_reg[19];
   assign h2c_gpio_14_gpio_18_f = h2c_gpio_14_reg[18];
   assign h2c_gpio_14_gpio_17_f = h2c_gpio_14_reg[17];
   assign h2c_gpio_14_gpio_16_f = h2c_gpio_14_reg[16];
   assign h2c_gpio_14_gpio_15_f = h2c_gpio_14_reg[15];
   assign h2c_gpio_14_gpio_14_f = h2c_gpio_14_reg[14];
   assign h2c_gpio_14_gpio_13_f = h2c_gpio_14_reg[13];
   assign h2c_gpio_14_gpio_12_f = h2c_gpio_14_reg[12];
   assign h2c_gpio_14_gpio_11_f = h2c_gpio_14_reg[11];
   assign h2c_gpio_14_gpio_10_f = h2c_gpio_14_reg[10];
   assign h2c_gpio_14_gpio_9_f = h2c_gpio_14_reg[9];
   assign h2c_gpio_14_gpio_8_f = h2c_gpio_14_reg[8];
   assign h2c_gpio_14_gpio_7_f = h2c_gpio_14_reg[7];
   assign h2c_gpio_14_gpio_6_f = h2c_gpio_14_reg[6];
   assign h2c_gpio_14_gpio_5_f = h2c_gpio_14_reg[5];
   assign h2c_gpio_14_gpio_4_f = h2c_gpio_14_reg[4];
   assign h2c_gpio_14_gpio_3_f = h2c_gpio_14_reg[3];
   assign h2c_gpio_14_gpio_2_f = h2c_gpio_14_reg[2];
   assign h2c_gpio_14_gpio_1_f = h2c_gpio_14_reg[1];
   assign h2c_gpio_14_gpio_0_f = h2c_gpio_14_reg[0];
   assign h2c_gpio_15_gpio_31_f = h2c_gpio_15_reg[31];
   assign h2c_gpio_15_gpio_30_f = h2c_gpio_15_reg[30];
   assign h2c_gpio_15_gpio_29_f = h2c_gpio_15_reg[29];
   assign h2c_gpio_15_gpio_28_f = h2c_gpio_15_reg[28];
   assign h2c_gpio_15_gpio_27_f = h2c_gpio_15_reg[27];
   assign h2c_gpio_15_gpio_26_f = h2c_gpio_15_reg[26];
   assign h2c_gpio_15_gpio_25_f = h2c_gpio_15_reg[25];
   assign h2c_gpio_15_gpio_24_f = h2c_gpio_15_reg[24];
   assign h2c_gpio_15_gpio_23_f = h2c_gpio_15_reg[23];
   assign h2c_gpio_15_gpio_22_f = h2c_gpio_15_reg[22];
   assign h2c_gpio_15_gpio_21_f = h2c_gpio_15_reg[21];
   assign h2c_gpio_15_gpio_20_f = h2c_gpio_15_reg[20];
   assign h2c_gpio_15_gpio_19_f = h2c_gpio_15_reg[19];
   assign h2c_gpio_15_gpio_18_f = h2c_gpio_15_reg[18];
   assign h2c_gpio_15_gpio_17_f = h2c_gpio_15_reg[17];
   assign h2c_gpio_15_gpio_16_f = h2c_gpio_15_reg[16];
   assign h2c_gpio_15_gpio_15_f = h2c_gpio_15_reg[15];
   assign h2c_gpio_15_gpio_14_f = h2c_gpio_15_reg[14];
   assign h2c_gpio_15_gpio_13_f = h2c_gpio_15_reg[13];
   assign h2c_gpio_15_gpio_12_f = h2c_gpio_15_reg[12];
   assign h2c_gpio_15_gpio_11_f = h2c_gpio_15_reg[11];
   assign h2c_gpio_15_gpio_10_f = h2c_gpio_15_reg[10];
   assign h2c_gpio_15_gpio_9_f = h2c_gpio_15_reg[9];
   assign h2c_gpio_15_gpio_8_f = h2c_gpio_15_reg[8];
   assign h2c_gpio_15_gpio_7_f = h2c_gpio_15_reg[7];
   assign h2c_gpio_15_gpio_6_f = h2c_gpio_15_reg[6];
   assign h2c_gpio_15_gpio_5_f = h2c_gpio_15_reg[5];
   assign h2c_gpio_15_gpio_4_f = h2c_gpio_15_reg[4];
   assign h2c_gpio_15_gpio_3_f = h2c_gpio_15_reg[3];
   assign h2c_gpio_15_gpio_2_f = h2c_gpio_15_reg[2];
   assign h2c_gpio_15_gpio_1_f = h2c_gpio_15_reg[1];
   assign h2c_gpio_15_gpio_0_f = h2c_gpio_15_reg[0];
   assign rd_req_desc_0_size_txn_size_f = rd_req_desc_0_size_reg[31:0];
   assign rd_req_desc_0_axsize_axsize_f = rd_req_desc_0_axsize_reg[2:0];
   assign rd_req_desc_0_attr_axsnoop_f = rd_req_desc_0_attr_reg[27:24];
   assign rd_req_desc_0_attr_axdomain_f = rd_req_desc_0_attr_reg[23:22];
   assign rd_req_desc_0_attr_axbar_f = rd_req_desc_0_attr_reg[21:20];
   assign rd_req_desc_0_attr_axregion_f = rd_req_desc_0_attr_reg[18:15];
   assign rd_req_desc_0_attr_axqos_f = rd_req_desc_0_attr_reg[14:11];
   assign rd_req_desc_0_attr_axprot_f = rd_req_desc_0_attr_reg[10:8];
   assign rd_req_desc_0_attr_axcache_f = rd_req_desc_0_attr_reg[7:4];
   assign rd_req_desc_0_attr_axlock_f = rd_req_desc_0_attr_reg[2];
   assign rd_req_desc_0_attr_axburst_f = rd_req_desc_0_attr_reg[1:0];
   assign rd_req_desc_0_axaddr_0_addr_f = rd_req_desc_0_axaddr_0_reg[31:0];
   assign rd_req_desc_0_axaddr_1_addr_f = rd_req_desc_0_axaddr_1_reg[31:0];
   assign rd_req_desc_0_axaddr_2_addr_f = rd_req_desc_0_axaddr_2_reg[31:0];
   assign rd_req_desc_0_axaddr_3_addr_f = rd_req_desc_0_axaddr_3_reg[31:0];
   assign rd_req_desc_0_axid_0_axid_f = rd_req_desc_0_axid_0_reg[31:0];
   assign rd_req_desc_0_axid_1_axid_f = rd_req_desc_0_axid_1_reg[31:0];
   assign rd_req_desc_0_axid_2_axid_f = rd_req_desc_0_axid_2_reg[31:0];
   assign rd_req_desc_0_axid_3_axid_f = rd_req_desc_0_axid_3_reg[31:0];
   assign rd_req_desc_0_axuser_0_axuser_f = rd_req_desc_0_axuser_0_reg[31:0];
   assign rd_req_desc_0_axuser_1_axuser_f = rd_req_desc_0_axuser_1_reg[31:0];
   assign rd_req_desc_0_axuser_2_axuser_f = rd_req_desc_0_axuser_2_reg[31:0];
   assign rd_req_desc_0_axuser_3_axuser_f = rd_req_desc_0_axuser_3_reg[31:0];
   assign rd_req_desc_0_axuser_4_axuser_f = rd_req_desc_0_axuser_4_reg[31:0];
   assign rd_req_desc_0_axuser_5_axuser_f = rd_req_desc_0_axuser_5_reg[31:0];
   assign rd_req_desc_0_axuser_6_axuser_f = rd_req_desc_0_axuser_6_reg[31:0];
   assign rd_req_desc_0_axuser_7_axuser_f = rd_req_desc_0_axuser_7_reg[31:0];
   assign rd_req_desc_0_axuser_8_axuser_f = rd_req_desc_0_axuser_8_reg[31:0];
   assign rd_req_desc_0_axuser_9_axuser_f = rd_req_desc_0_axuser_9_reg[31:0];
   assign rd_req_desc_0_axuser_10_axuser_f = rd_req_desc_0_axuser_10_reg[31:0];
   assign rd_req_desc_0_axuser_11_axuser_f = rd_req_desc_0_axuser_11_reg[31:0];
   assign rd_req_desc_0_axuser_12_axuser_f = rd_req_desc_0_axuser_12_reg[31:0];
   assign rd_req_desc_0_axuser_13_axuser_f = rd_req_desc_0_axuser_13_reg[31:0];
   assign rd_req_desc_0_axuser_14_axuser_f = rd_req_desc_0_axuser_14_reg[31:0];
   assign rd_req_desc_0_axuser_15_axuser_f = rd_req_desc_0_axuser_15_reg[31:0];
   assign rd_resp_desc_0_data_offset_addr_f = rd_resp_desc_0_data_offset_reg[13:0];
   assign rd_resp_desc_0_data_size_size_f = rd_resp_desc_0_data_size_reg[31:0];
   assign rd_resp_desc_0_data_host_addr_0_addr_f = rd_resp_desc_0_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_0_data_host_addr_1_addr_f = rd_resp_desc_0_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_0_data_host_addr_2_addr_f = rd_resp_desc_0_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_0_data_host_addr_3_addr_f = rd_resp_desc_0_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_0_resp_resp_f = rd_resp_desc_0_resp_reg[4:0];
   assign rd_resp_desc_0_xid_0_xid_f = rd_resp_desc_0_xid_0_reg[31:0];
   assign rd_resp_desc_0_xid_1_xid_f = rd_resp_desc_0_xid_1_reg[31:0];
   assign rd_resp_desc_0_xid_2_xid_f = rd_resp_desc_0_xid_2_reg[31:0];
   assign rd_resp_desc_0_xid_3_xid_f = rd_resp_desc_0_xid_3_reg[31:0];
   assign rd_resp_desc_0_xuser_0_xuser_f = rd_resp_desc_0_xuser_0_reg[31:0];
   assign rd_resp_desc_0_xuser_1_xuser_f = rd_resp_desc_0_xuser_1_reg[31:0];
   assign rd_resp_desc_0_xuser_2_xuser_f = rd_resp_desc_0_xuser_2_reg[31:0];
   assign rd_resp_desc_0_xuser_3_xuser_f = rd_resp_desc_0_xuser_3_reg[31:0];
   assign rd_resp_desc_0_xuser_4_xuser_f = rd_resp_desc_0_xuser_4_reg[31:0];
   assign rd_resp_desc_0_xuser_5_xuser_f = rd_resp_desc_0_xuser_5_reg[31:0];
   assign rd_resp_desc_0_xuser_6_xuser_f = rd_resp_desc_0_xuser_6_reg[31:0];
   assign rd_resp_desc_0_xuser_7_xuser_f = rd_resp_desc_0_xuser_7_reg[31:0];
   assign rd_resp_desc_0_xuser_8_xuser_f = rd_resp_desc_0_xuser_8_reg[31:0];
   assign rd_resp_desc_0_xuser_9_xuser_f = rd_resp_desc_0_xuser_9_reg[31:0];
   assign rd_resp_desc_0_xuser_10_xuser_f = rd_resp_desc_0_xuser_10_reg[31:0];
   assign rd_resp_desc_0_xuser_11_xuser_f = rd_resp_desc_0_xuser_11_reg[31:0];
   assign rd_resp_desc_0_xuser_12_xuser_f = rd_resp_desc_0_xuser_12_reg[31:0];
   assign rd_resp_desc_0_xuser_13_xuser_f = rd_resp_desc_0_xuser_13_reg[31:0];
   assign rd_resp_desc_0_xuser_14_xuser_f = rd_resp_desc_0_xuser_14_reg[31:0];
   assign rd_resp_desc_0_xuser_15_xuser_f = rd_resp_desc_0_xuser_15_reg[31:0];
   assign wr_req_desc_0_txn_type_wr_strb_f = wr_req_desc_0_txn_type_reg[1];
   assign wr_req_desc_0_size_txn_size_f = wr_req_desc_0_size_reg[31:0];
   assign wr_req_desc_0_data_offset_addr_f = wr_req_desc_0_data_offset_reg[13:0];
   assign wr_req_desc_0_data_host_addr_0_addr_f = wr_req_desc_0_data_host_addr_0_reg[31:0];
   assign wr_req_desc_0_data_host_addr_1_addr_f = wr_req_desc_0_data_host_addr_1_reg[31:0];
   assign wr_req_desc_0_data_host_addr_2_addr_f = wr_req_desc_0_data_host_addr_2_reg[31:0];
   assign wr_req_desc_0_data_host_addr_3_addr_f = wr_req_desc_0_data_host_addr_3_reg[31:0];
   assign wr_req_desc_0_wstrb_host_addr_0_addr_f = wr_req_desc_0_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_0_wstrb_host_addr_1_addr_f = wr_req_desc_0_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_0_wstrb_host_addr_2_addr_f = wr_req_desc_0_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_0_wstrb_host_addr_3_addr_f = wr_req_desc_0_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_0_axsize_axsize_f = wr_req_desc_0_axsize_reg[2:0];
   assign wr_req_desc_0_attr_axsnoop_f = wr_req_desc_0_attr_reg[27:24];
   assign wr_req_desc_0_attr_axdomain_f = wr_req_desc_0_attr_reg[23:22];
   assign wr_req_desc_0_attr_axbar_f = wr_req_desc_0_attr_reg[21:20];
   assign wr_req_desc_0_attr_awunique_f = wr_req_desc_0_attr_reg[19];
   assign wr_req_desc_0_attr_axregion_f = wr_req_desc_0_attr_reg[18:15];
   assign wr_req_desc_0_attr_axqos_f = wr_req_desc_0_attr_reg[14:11];
   assign wr_req_desc_0_attr_axprot_f = wr_req_desc_0_attr_reg[10:8];
   assign wr_req_desc_0_attr_axcache_f = wr_req_desc_0_attr_reg[7:4];
   assign wr_req_desc_0_attr_axlock_f = wr_req_desc_0_attr_reg[2];
   assign wr_req_desc_0_attr_axburst_f = wr_req_desc_0_attr_reg[1:0];
   assign wr_req_desc_0_axaddr_0_addr_f = wr_req_desc_0_axaddr_0_reg[31:0];
   assign wr_req_desc_0_axaddr_1_addr_f = wr_req_desc_0_axaddr_1_reg[31:0];
   assign wr_req_desc_0_axaddr_2_addr_f = wr_req_desc_0_axaddr_2_reg[31:0];
   assign wr_req_desc_0_axaddr_3_addr_f = wr_req_desc_0_axaddr_3_reg[31:0];
   assign wr_req_desc_0_axid_0_axid_f = wr_req_desc_0_axid_0_reg[31:0];
   assign wr_req_desc_0_axid_1_axid_f = wr_req_desc_0_axid_1_reg[31:0];
   assign wr_req_desc_0_axid_2_axid_f = wr_req_desc_0_axid_2_reg[31:0];
   assign wr_req_desc_0_axid_3_axid_f = wr_req_desc_0_axid_3_reg[31:0];
   assign wr_req_desc_0_axuser_0_axuser_f = wr_req_desc_0_axuser_0_reg[31:0];
   assign wr_req_desc_0_axuser_1_axuser_f = wr_req_desc_0_axuser_1_reg[31:0];
   assign wr_req_desc_0_axuser_2_axuser_f = wr_req_desc_0_axuser_2_reg[31:0];
   assign wr_req_desc_0_axuser_3_axuser_f = wr_req_desc_0_axuser_3_reg[31:0];
   assign wr_req_desc_0_axuser_4_axuser_f = wr_req_desc_0_axuser_4_reg[31:0];
   assign wr_req_desc_0_axuser_5_axuser_f = wr_req_desc_0_axuser_5_reg[31:0];
   assign wr_req_desc_0_axuser_6_axuser_f = wr_req_desc_0_axuser_6_reg[31:0];
   assign wr_req_desc_0_axuser_7_axuser_f = wr_req_desc_0_axuser_7_reg[31:0];
   assign wr_req_desc_0_axuser_8_axuser_f = wr_req_desc_0_axuser_8_reg[31:0];
   assign wr_req_desc_0_axuser_9_axuser_f = wr_req_desc_0_axuser_9_reg[31:0];
   assign wr_req_desc_0_axuser_10_axuser_f = wr_req_desc_0_axuser_10_reg[31:0];
   assign wr_req_desc_0_axuser_11_axuser_f = wr_req_desc_0_axuser_11_reg[31:0];
   assign wr_req_desc_0_axuser_12_axuser_f = wr_req_desc_0_axuser_12_reg[31:0];
   assign wr_req_desc_0_axuser_13_axuser_f = wr_req_desc_0_axuser_13_reg[31:0];
   assign wr_req_desc_0_axuser_14_axuser_f = wr_req_desc_0_axuser_14_reg[31:0];
   assign wr_req_desc_0_axuser_15_axuser_f = wr_req_desc_0_axuser_15_reg[31:0];
   assign wr_req_desc_0_wuser_0_wuser_f = wr_req_desc_0_wuser_0_reg[31:0];
   assign wr_req_desc_0_wuser_1_wuser_f = wr_req_desc_0_wuser_1_reg[31:0];
   assign wr_req_desc_0_wuser_2_wuser_f = wr_req_desc_0_wuser_2_reg[31:0];
   assign wr_req_desc_0_wuser_3_wuser_f = wr_req_desc_0_wuser_3_reg[31:0];
   assign wr_req_desc_0_wuser_4_wuser_f = wr_req_desc_0_wuser_4_reg[31:0];
   assign wr_req_desc_0_wuser_5_wuser_f = wr_req_desc_0_wuser_5_reg[31:0];
   assign wr_req_desc_0_wuser_6_wuser_f = wr_req_desc_0_wuser_6_reg[31:0];
   assign wr_req_desc_0_wuser_7_wuser_f = wr_req_desc_0_wuser_7_reg[31:0];
   assign wr_req_desc_0_wuser_8_wuser_f = wr_req_desc_0_wuser_8_reg[31:0];
   assign wr_req_desc_0_wuser_9_wuser_f = wr_req_desc_0_wuser_9_reg[31:0];
   assign wr_req_desc_0_wuser_10_wuser_f = wr_req_desc_0_wuser_10_reg[31:0];
   assign wr_req_desc_0_wuser_11_wuser_f = wr_req_desc_0_wuser_11_reg[31:0];
   assign wr_req_desc_0_wuser_12_wuser_f = wr_req_desc_0_wuser_12_reg[31:0];
   assign wr_req_desc_0_wuser_13_wuser_f = wr_req_desc_0_wuser_13_reg[31:0];
   assign wr_req_desc_0_wuser_14_wuser_f = wr_req_desc_0_wuser_14_reg[31:0];
   assign wr_req_desc_0_wuser_15_wuser_f = wr_req_desc_0_wuser_15_reg[31:0];
   assign wr_resp_desc_0_resp_resp_f = wr_resp_desc_0_resp_reg[4:0];
   assign wr_resp_desc_0_xid_0_xid_f = wr_resp_desc_0_xid_0_reg[31:0];
   assign wr_resp_desc_0_xid_1_xid_f = wr_resp_desc_0_xid_1_reg[31:0];
   assign wr_resp_desc_0_xid_2_xid_f = wr_resp_desc_0_xid_2_reg[31:0];
   assign wr_resp_desc_0_xid_3_xid_f = wr_resp_desc_0_xid_3_reg[31:0];
   assign wr_resp_desc_0_xuser_0_xuser_f = wr_resp_desc_0_xuser_0_reg[31:0];
   assign wr_resp_desc_0_xuser_1_xuser_f = wr_resp_desc_0_xuser_1_reg[31:0];
   assign wr_resp_desc_0_xuser_2_xuser_f = wr_resp_desc_0_xuser_2_reg[31:0];
   assign wr_resp_desc_0_xuser_3_xuser_f = wr_resp_desc_0_xuser_3_reg[31:0];
   assign wr_resp_desc_0_xuser_4_xuser_f = wr_resp_desc_0_xuser_4_reg[31:0];
   assign wr_resp_desc_0_xuser_5_xuser_f = wr_resp_desc_0_xuser_5_reg[31:0];
   assign wr_resp_desc_0_xuser_6_xuser_f = wr_resp_desc_0_xuser_6_reg[31:0];
   assign wr_resp_desc_0_xuser_7_xuser_f = wr_resp_desc_0_xuser_7_reg[31:0];
   assign wr_resp_desc_0_xuser_8_xuser_f = wr_resp_desc_0_xuser_8_reg[31:0];
   assign wr_resp_desc_0_xuser_9_xuser_f = wr_resp_desc_0_xuser_9_reg[31:0];
   assign wr_resp_desc_0_xuser_10_xuser_f = wr_resp_desc_0_xuser_10_reg[31:0];
   assign wr_resp_desc_0_xuser_11_xuser_f = wr_resp_desc_0_xuser_11_reg[31:0];
   assign wr_resp_desc_0_xuser_12_xuser_f = wr_resp_desc_0_xuser_12_reg[31:0];
   assign wr_resp_desc_0_xuser_13_xuser_f = wr_resp_desc_0_xuser_13_reg[31:0];
   assign wr_resp_desc_0_xuser_14_xuser_f = wr_resp_desc_0_xuser_14_reg[31:0];
   assign wr_resp_desc_0_xuser_15_xuser_f = wr_resp_desc_0_xuser_15_reg[31:0];
   assign sn_req_desc_0_attr_acsnoop_f = sn_req_desc_0_attr_reg[27:24];
   assign sn_req_desc_0_attr_acprot_f = sn_req_desc_0_attr_reg[10:8];
   assign sn_req_desc_0_acaddr_0_addr_f = sn_req_desc_0_acaddr_0_reg[31:0];
   assign sn_req_desc_0_acaddr_1_addr_f = sn_req_desc_0_acaddr_1_reg[31:0];
   assign sn_req_desc_0_acaddr_2_addr_f = sn_req_desc_0_acaddr_2_reg[31:0];
   assign sn_req_desc_0_acaddr_3_addr_f = sn_req_desc_0_acaddr_3_reg[31:0];
   assign sn_resp_desc_0_resp_resp_f = sn_resp_desc_0_resp_reg[4:0];
   assign rd_req_desc_1_size_txn_size_f = rd_req_desc_1_size_reg[31:0];
   assign rd_req_desc_1_axsize_axsize_f = rd_req_desc_1_axsize_reg[2:0];
   assign rd_req_desc_1_attr_axsnoop_f = rd_req_desc_1_attr_reg[27:24];
   assign rd_req_desc_1_attr_axdomain_f = rd_req_desc_1_attr_reg[23:22];
   assign rd_req_desc_1_attr_axbar_f = rd_req_desc_1_attr_reg[21:20];
   assign rd_req_desc_1_attr_axregion_f = rd_req_desc_1_attr_reg[18:15];
   assign rd_req_desc_1_attr_axqos_f = rd_req_desc_1_attr_reg[14:11];
   assign rd_req_desc_1_attr_axprot_f = rd_req_desc_1_attr_reg[10:8];
   assign rd_req_desc_1_attr_axcache_f = rd_req_desc_1_attr_reg[7:4];
   assign rd_req_desc_1_attr_axlock_f = rd_req_desc_1_attr_reg[2];
   assign rd_req_desc_1_attr_axburst_f = rd_req_desc_1_attr_reg[1:0];
   assign rd_req_desc_1_axaddr_0_addr_f = rd_req_desc_1_axaddr_0_reg[31:0];
   assign rd_req_desc_1_axaddr_1_addr_f = rd_req_desc_1_axaddr_1_reg[31:0];
   assign rd_req_desc_1_axaddr_2_addr_f = rd_req_desc_1_axaddr_2_reg[31:0];
   assign rd_req_desc_1_axaddr_3_addr_f = rd_req_desc_1_axaddr_3_reg[31:0];
   assign rd_req_desc_1_axid_0_axid_f = rd_req_desc_1_axid_0_reg[31:0];
   assign rd_req_desc_1_axid_1_axid_f = rd_req_desc_1_axid_1_reg[31:0];
   assign rd_req_desc_1_axid_2_axid_f = rd_req_desc_1_axid_2_reg[31:0];
   assign rd_req_desc_1_axid_3_axid_f = rd_req_desc_1_axid_3_reg[31:0];
   assign rd_req_desc_1_axuser_0_axuser_f = rd_req_desc_1_axuser_0_reg[31:0];
   assign rd_req_desc_1_axuser_1_axuser_f = rd_req_desc_1_axuser_1_reg[31:0];
   assign rd_req_desc_1_axuser_2_axuser_f = rd_req_desc_1_axuser_2_reg[31:0];
   assign rd_req_desc_1_axuser_3_axuser_f = rd_req_desc_1_axuser_3_reg[31:0];
   assign rd_req_desc_1_axuser_4_axuser_f = rd_req_desc_1_axuser_4_reg[31:0];
   assign rd_req_desc_1_axuser_5_axuser_f = rd_req_desc_1_axuser_5_reg[31:0];
   assign rd_req_desc_1_axuser_6_axuser_f = rd_req_desc_1_axuser_6_reg[31:0];
   assign rd_req_desc_1_axuser_7_axuser_f = rd_req_desc_1_axuser_7_reg[31:0];
   assign rd_req_desc_1_axuser_8_axuser_f = rd_req_desc_1_axuser_8_reg[31:0];
   assign rd_req_desc_1_axuser_9_axuser_f = rd_req_desc_1_axuser_9_reg[31:0];
   assign rd_req_desc_1_axuser_10_axuser_f = rd_req_desc_1_axuser_10_reg[31:0];
   assign rd_req_desc_1_axuser_11_axuser_f = rd_req_desc_1_axuser_11_reg[31:0];
   assign rd_req_desc_1_axuser_12_axuser_f = rd_req_desc_1_axuser_12_reg[31:0];
   assign rd_req_desc_1_axuser_13_axuser_f = rd_req_desc_1_axuser_13_reg[31:0];
   assign rd_req_desc_1_axuser_14_axuser_f = rd_req_desc_1_axuser_14_reg[31:0];
   assign rd_req_desc_1_axuser_15_axuser_f = rd_req_desc_1_axuser_15_reg[31:0];
   assign rd_resp_desc_1_data_offset_addr_f = rd_resp_desc_1_data_offset_reg[13:0];
   assign rd_resp_desc_1_data_size_size_f = rd_resp_desc_1_data_size_reg[31:0];
   assign rd_resp_desc_1_data_host_addr_0_addr_f = rd_resp_desc_1_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_1_data_host_addr_1_addr_f = rd_resp_desc_1_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_1_data_host_addr_2_addr_f = rd_resp_desc_1_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_1_data_host_addr_3_addr_f = rd_resp_desc_1_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_1_resp_resp_f = rd_resp_desc_1_resp_reg[4:0];
   assign rd_resp_desc_1_xid_0_xid_f = rd_resp_desc_1_xid_0_reg[31:0];
   assign rd_resp_desc_1_xid_1_xid_f = rd_resp_desc_1_xid_1_reg[31:0];
   assign rd_resp_desc_1_xid_2_xid_f = rd_resp_desc_1_xid_2_reg[31:0];
   assign rd_resp_desc_1_xid_3_xid_f = rd_resp_desc_1_xid_3_reg[31:0];
   assign rd_resp_desc_1_xuser_0_xuser_f = rd_resp_desc_1_xuser_0_reg[31:0];
   assign rd_resp_desc_1_xuser_1_xuser_f = rd_resp_desc_1_xuser_1_reg[31:0];
   assign rd_resp_desc_1_xuser_2_xuser_f = rd_resp_desc_1_xuser_2_reg[31:0];
   assign rd_resp_desc_1_xuser_3_xuser_f = rd_resp_desc_1_xuser_3_reg[31:0];
   assign rd_resp_desc_1_xuser_4_xuser_f = rd_resp_desc_1_xuser_4_reg[31:0];
   assign rd_resp_desc_1_xuser_5_xuser_f = rd_resp_desc_1_xuser_5_reg[31:0];
   assign rd_resp_desc_1_xuser_6_xuser_f = rd_resp_desc_1_xuser_6_reg[31:0];
   assign rd_resp_desc_1_xuser_7_xuser_f = rd_resp_desc_1_xuser_7_reg[31:0];
   assign rd_resp_desc_1_xuser_8_xuser_f = rd_resp_desc_1_xuser_8_reg[31:0];
   assign rd_resp_desc_1_xuser_9_xuser_f = rd_resp_desc_1_xuser_9_reg[31:0];
   assign rd_resp_desc_1_xuser_10_xuser_f = rd_resp_desc_1_xuser_10_reg[31:0];
   assign rd_resp_desc_1_xuser_11_xuser_f = rd_resp_desc_1_xuser_11_reg[31:0];
   assign rd_resp_desc_1_xuser_12_xuser_f = rd_resp_desc_1_xuser_12_reg[31:0];
   assign rd_resp_desc_1_xuser_13_xuser_f = rd_resp_desc_1_xuser_13_reg[31:0];
   assign rd_resp_desc_1_xuser_14_xuser_f = rd_resp_desc_1_xuser_14_reg[31:0];
   assign rd_resp_desc_1_xuser_15_xuser_f = rd_resp_desc_1_xuser_15_reg[31:0];
   assign wr_req_desc_1_txn_type_wr_strb_f = wr_req_desc_1_txn_type_reg[1];
   assign wr_req_desc_1_size_txn_size_f = wr_req_desc_1_size_reg[31:0];
   assign wr_req_desc_1_data_offset_addr_f = wr_req_desc_1_data_offset_reg[13:0];
   assign wr_req_desc_1_data_host_addr_0_addr_f = wr_req_desc_1_data_host_addr_0_reg[31:0];
   assign wr_req_desc_1_data_host_addr_1_addr_f = wr_req_desc_1_data_host_addr_1_reg[31:0];
   assign wr_req_desc_1_data_host_addr_2_addr_f = wr_req_desc_1_data_host_addr_2_reg[31:0];
   assign wr_req_desc_1_data_host_addr_3_addr_f = wr_req_desc_1_data_host_addr_3_reg[31:0];
   assign wr_req_desc_1_wstrb_host_addr_0_addr_f = wr_req_desc_1_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_1_wstrb_host_addr_1_addr_f = wr_req_desc_1_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_1_wstrb_host_addr_2_addr_f = wr_req_desc_1_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_1_wstrb_host_addr_3_addr_f = wr_req_desc_1_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_1_axsize_axsize_f = wr_req_desc_1_axsize_reg[2:0];
   assign wr_req_desc_1_attr_axsnoop_f = wr_req_desc_1_attr_reg[27:24];
   assign wr_req_desc_1_attr_axdomain_f = wr_req_desc_1_attr_reg[23:22];
   assign wr_req_desc_1_attr_axbar_f = wr_req_desc_1_attr_reg[21:20];
   assign wr_req_desc_1_attr_awunique_f = wr_req_desc_1_attr_reg[19];
   assign wr_req_desc_1_attr_axregion_f = wr_req_desc_1_attr_reg[18:15];
   assign wr_req_desc_1_attr_axqos_f = wr_req_desc_1_attr_reg[14:11];
   assign wr_req_desc_1_attr_axprot_f = wr_req_desc_1_attr_reg[10:8];
   assign wr_req_desc_1_attr_axcache_f = wr_req_desc_1_attr_reg[7:4];
   assign wr_req_desc_1_attr_axlock_f = wr_req_desc_1_attr_reg[2];
   assign wr_req_desc_1_attr_axburst_f = wr_req_desc_1_attr_reg[1:0];
   assign wr_req_desc_1_axaddr_0_addr_f = wr_req_desc_1_axaddr_0_reg[31:0];
   assign wr_req_desc_1_axaddr_1_addr_f = wr_req_desc_1_axaddr_1_reg[31:0];
   assign wr_req_desc_1_axaddr_2_addr_f = wr_req_desc_1_axaddr_2_reg[31:0];
   assign wr_req_desc_1_axaddr_3_addr_f = wr_req_desc_1_axaddr_3_reg[31:0];
   assign wr_req_desc_1_axid_0_axid_f = wr_req_desc_1_axid_0_reg[31:0];
   assign wr_req_desc_1_axid_1_axid_f = wr_req_desc_1_axid_1_reg[31:0];
   assign wr_req_desc_1_axid_2_axid_f = wr_req_desc_1_axid_2_reg[31:0];
   assign wr_req_desc_1_axid_3_axid_f = wr_req_desc_1_axid_3_reg[31:0];
   assign wr_req_desc_1_axuser_0_axuser_f = wr_req_desc_1_axuser_0_reg[31:0];
   assign wr_req_desc_1_axuser_1_axuser_f = wr_req_desc_1_axuser_1_reg[31:0];
   assign wr_req_desc_1_axuser_2_axuser_f = wr_req_desc_1_axuser_2_reg[31:0];
   assign wr_req_desc_1_axuser_3_axuser_f = wr_req_desc_1_axuser_3_reg[31:0];
   assign wr_req_desc_1_axuser_4_axuser_f = wr_req_desc_1_axuser_4_reg[31:0];
   assign wr_req_desc_1_axuser_5_axuser_f = wr_req_desc_1_axuser_5_reg[31:0];
   assign wr_req_desc_1_axuser_6_axuser_f = wr_req_desc_1_axuser_6_reg[31:0];
   assign wr_req_desc_1_axuser_7_axuser_f = wr_req_desc_1_axuser_7_reg[31:0];
   assign wr_req_desc_1_axuser_8_axuser_f = wr_req_desc_1_axuser_8_reg[31:0];
   assign wr_req_desc_1_axuser_9_axuser_f = wr_req_desc_1_axuser_9_reg[31:0];
   assign wr_req_desc_1_axuser_10_axuser_f = wr_req_desc_1_axuser_10_reg[31:0];
   assign wr_req_desc_1_axuser_11_axuser_f = wr_req_desc_1_axuser_11_reg[31:0];
   assign wr_req_desc_1_axuser_12_axuser_f = wr_req_desc_1_axuser_12_reg[31:0];
   assign wr_req_desc_1_axuser_13_axuser_f = wr_req_desc_1_axuser_13_reg[31:0];
   assign wr_req_desc_1_axuser_14_axuser_f = wr_req_desc_1_axuser_14_reg[31:0];
   assign wr_req_desc_1_axuser_15_axuser_f = wr_req_desc_1_axuser_15_reg[31:0];
   assign wr_req_desc_1_wuser_0_wuser_f = wr_req_desc_1_wuser_0_reg[31:0];
   assign wr_req_desc_1_wuser_1_wuser_f = wr_req_desc_1_wuser_1_reg[31:0];
   assign wr_req_desc_1_wuser_2_wuser_f = wr_req_desc_1_wuser_2_reg[31:0];
   assign wr_req_desc_1_wuser_3_wuser_f = wr_req_desc_1_wuser_3_reg[31:0];
   assign wr_req_desc_1_wuser_4_wuser_f = wr_req_desc_1_wuser_4_reg[31:0];
   assign wr_req_desc_1_wuser_5_wuser_f = wr_req_desc_1_wuser_5_reg[31:0];
   assign wr_req_desc_1_wuser_6_wuser_f = wr_req_desc_1_wuser_6_reg[31:0];
   assign wr_req_desc_1_wuser_7_wuser_f = wr_req_desc_1_wuser_7_reg[31:0];
   assign wr_req_desc_1_wuser_8_wuser_f = wr_req_desc_1_wuser_8_reg[31:0];
   assign wr_req_desc_1_wuser_9_wuser_f = wr_req_desc_1_wuser_9_reg[31:0];
   assign wr_req_desc_1_wuser_10_wuser_f = wr_req_desc_1_wuser_10_reg[31:0];
   assign wr_req_desc_1_wuser_11_wuser_f = wr_req_desc_1_wuser_11_reg[31:0];
   assign wr_req_desc_1_wuser_12_wuser_f = wr_req_desc_1_wuser_12_reg[31:0];
   assign wr_req_desc_1_wuser_13_wuser_f = wr_req_desc_1_wuser_13_reg[31:0];
   assign wr_req_desc_1_wuser_14_wuser_f = wr_req_desc_1_wuser_14_reg[31:0];
   assign wr_req_desc_1_wuser_15_wuser_f = wr_req_desc_1_wuser_15_reg[31:0];
   assign wr_resp_desc_1_resp_resp_f = wr_resp_desc_1_resp_reg[4:0];
   assign wr_resp_desc_1_xid_0_xid_f = wr_resp_desc_1_xid_0_reg[31:0];
   assign wr_resp_desc_1_xid_1_xid_f = wr_resp_desc_1_xid_1_reg[31:0];
   assign wr_resp_desc_1_xid_2_xid_f = wr_resp_desc_1_xid_2_reg[31:0];
   assign wr_resp_desc_1_xid_3_xid_f = wr_resp_desc_1_xid_3_reg[31:0];
   assign wr_resp_desc_1_xuser_0_xuser_f = wr_resp_desc_1_xuser_0_reg[31:0];
   assign wr_resp_desc_1_xuser_1_xuser_f = wr_resp_desc_1_xuser_1_reg[31:0];
   assign wr_resp_desc_1_xuser_2_xuser_f = wr_resp_desc_1_xuser_2_reg[31:0];
   assign wr_resp_desc_1_xuser_3_xuser_f = wr_resp_desc_1_xuser_3_reg[31:0];
   assign wr_resp_desc_1_xuser_4_xuser_f = wr_resp_desc_1_xuser_4_reg[31:0];
   assign wr_resp_desc_1_xuser_5_xuser_f = wr_resp_desc_1_xuser_5_reg[31:0];
   assign wr_resp_desc_1_xuser_6_xuser_f = wr_resp_desc_1_xuser_6_reg[31:0];
   assign wr_resp_desc_1_xuser_7_xuser_f = wr_resp_desc_1_xuser_7_reg[31:0];
   assign wr_resp_desc_1_xuser_8_xuser_f = wr_resp_desc_1_xuser_8_reg[31:0];
   assign wr_resp_desc_1_xuser_9_xuser_f = wr_resp_desc_1_xuser_9_reg[31:0];
   assign wr_resp_desc_1_xuser_10_xuser_f = wr_resp_desc_1_xuser_10_reg[31:0];
   assign wr_resp_desc_1_xuser_11_xuser_f = wr_resp_desc_1_xuser_11_reg[31:0];
   assign wr_resp_desc_1_xuser_12_xuser_f = wr_resp_desc_1_xuser_12_reg[31:0];
   assign wr_resp_desc_1_xuser_13_xuser_f = wr_resp_desc_1_xuser_13_reg[31:0];
   assign wr_resp_desc_1_xuser_14_xuser_f = wr_resp_desc_1_xuser_14_reg[31:0];
   assign wr_resp_desc_1_xuser_15_xuser_f = wr_resp_desc_1_xuser_15_reg[31:0];
   assign sn_req_desc_1_attr_acsnoop_f = sn_req_desc_1_attr_reg[27:24];
   assign sn_req_desc_1_attr_acprot_f = sn_req_desc_1_attr_reg[10:8];
   assign sn_req_desc_1_acaddr_0_addr_f = sn_req_desc_1_acaddr_0_reg[31:0];
   assign sn_req_desc_1_acaddr_1_addr_f = sn_req_desc_1_acaddr_1_reg[31:0];
   assign sn_req_desc_1_acaddr_2_addr_f = sn_req_desc_1_acaddr_2_reg[31:0];
   assign sn_req_desc_1_acaddr_3_addr_f = sn_req_desc_1_acaddr_3_reg[31:0];
   assign sn_resp_desc_1_resp_resp_f = sn_resp_desc_1_resp_reg[4:0];
   assign rd_req_desc_2_size_txn_size_f = rd_req_desc_2_size_reg[31:0];
   assign rd_req_desc_2_axsize_axsize_f = rd_req_desc_2_axsize_reg[2:0];
   assign rd_req_desc_2_attr_axsnoop_f = rd_req_desc_2_attr_reg[27:24];
   assign rd_req_desc_2_attr_axdomain_f = rd_req_desc_2_attr_reg[23:22];
   assign rd_req_desc_2_attr_axbar_f = rd_req_desc_2_attr_reg[21:20];
   assign rd_req_desc_2_attr_axregion_f = rd_req_desc_2_attr_reg[18:15];
   assign rd_req_desc_2_attr_axqos_f = rd_req_desc_2_attr_reg[14:11];
   assign rd_req_desc_2_attr_axprot_f = rd_req_desc_2_attr_reg[10:8];
   assign rd_req_desc_2_attr_axcache_f = rd_req_desc_2_attr_reg[7:4];
   assign rd_req_desc_2_attr_axlock_f = rd_req_desc_2_attr_reg[2];
   assign rd_req_desc_2_attr_axburst_f = rd_req_desc_2_attr_reg[1:0];
   assign rd_req_desc_2_axaddr_0_addr_f = rd_req_desc_2_axaddr_0_reg[31:0];
   assign rd_req_desc_2_axaddr_1_addr_f = rd_req_desc_2_axaddr_1_reg[31:0];
   assign rd_req_desc_2_axaddr_2_addr_f = rd_req_desc_2_axaddr_2_reg[31:0];
   assign rd_req_desc_2_axaddr_3_addr_f = rd_req_desc_2_axaddr_3_reg[31:0];
   assign rd_req_desc_2_axid_0_axid_f = rd_req_desc_2_axid_0_reg[31:0];
   assign rd_req_desc_2_axid_1_axid_f = rd_req_desc_2_axid_1_reg[31:0];
   assign rd_req_desc_2_axid_2_axid_f = rd_req_desc_2_axid_2_reg[31:0];
   assign rd_req_desc_2_axid_3_axid_f = rd_req_desc_2_axid_3_reg[31:0];
   assign rd_req_desc_2_axuser_0_axuser_f = rd_req_desc_2_axuser_0_reg[31:0];
   assign rd_req_desc_2_axuser_1_axuser_f = rd_req_desc_2_axuser_1_reg[31:0];
   assign rd_req_desc_2_axuser_2_axuser_f = rd_req_desc_2_axuser_2_reg[31:0];
   assign rd_req_desc_2_axuser_3_axuser_f = rd_req_desc_2_axuser_3_reg[31:0];
   assign rd_req_desc_2_axuser_4_axuser_f = rd_req_desc_2_axuser_4_reg[31:0];
   assign rd_req_desc_2_axuser_5_axuser_f = rd_req_desc_2_axuser_5_reg[31:0];
   assign rd_req_desc_2_axuser_6_axuser_f = rd_req_desc_2_axuser_6_reg[31:0];
   assign rd_req_desc_2_axuser_7_axuser_f = rd_req_desc_2_axuser_7_reg[31:0];
   assign rd_req_desc_2_axuser_8_axuser_f = rd_req_desc_2_axuser_8_reg[31:0];
   assign rd_req_desc_2_axuser_9_axuser_f = rd_req_desc_2_axuser_9_reg[31:0];
   assign rd_req_desc_2_axuser_10_axuser_f = rd_req_desc_2_axuser_10_reg[31:0];
   assign rd_req_desc_2_axuser_11_axuser_f = rd_req_desc_2_axuser_11_reg[31:0];
   assign rd_req_desc_2_axuser_12_axuser_f = rd_req_desc_2_axuser_12_reg[31:0];
   assign rd_req_desc_2_axuser_13_axuser_f = rd_req_desc_2_axuser_13_reg[31:0];
   assign rd_req_desc_2_axuser_14_axuser_f = rd_req_desc_2_axuser_14_reg[31:0];
   assign rd_req_desc_2_axuser_15_axuser_f = rd_req_desc_2_axuser_15_reg[31:0];
   assign rd_resp_desc_2_data_offset_addr_f = rd_resp_desc_2_data_offset_reg[13:0];
   assign rd_resp_desc_2_data_size_size_f = rd_resp_desc_2_data_size_reg[31:0];
   assign rd_resp_desc_2_data_host_addr_0_addr_f = rd_resp_desc_2_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_2_data_host_addr_1_addr_f = rd_resp_desc_2_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_2_data_host_addr_2_addr_f = rd_resp_desc_2_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_2_data_host_addr_3_addr_f = rd_resp_desc_2_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_2_resp_resp_f = rd_resp_desc_2_resp_reg[4:0];
   assign rd_resp_desc_2_xid_0_xid_f = rd_resp_desc_2_xid_0_reg[31:0];
   assign rd_resp_desc_2_xid_1_xid_f = rd_resp_desc_2_xid_1_reg[31:0];
   assign rd_resp_desc_2_xid_2_xid_f = rd_resp_desc_2_xid_2_reg[31:0];
   assign rd_resp_desc_2_xid_3_xid_f = rd_resp_desc_2_xid_3_reg[31:0];
   assign rd_resp_desc_2_xuser_0_xuser_f = rd_resp_desc_2_xuser_0_reg[31:0];
   assign rd_resp_desc_2_xuser_1_xuser_f = rd_resp_desc_2_xuser_1_reg[31:0];
   assign rd_resp_desc_2_xuser_2_xuser_f = rd_resp_desc_2_xuser_2_reg[31:0];
   assign rd_resp_desc_2_xuser_3_xuser_f = rd_resp_desc_2_xuser_3_reg[31:0];
   assign rd_resp_desc_2_xuser_4_xuser_f = rd_resp_desc_2_xuser_4_reg[31:0];
   assign rd_resp_desc_2_xuser_5_xuser_f = rd_resp_desc_2_xuser_5_reg[31:0];
   assign rd_resp_desc_2_xuser_6_xuser_f = rd_resp_desc_2_xuser_6_reg[31:0];
   assign rd_resp_desc_2_xuser_7_xuser_f = rd_resp_desc_2_xuser_7_reg[31:0];
   assign rd_resp_desc_2_xuser_8_xuser_f = rd_resp_desc_2_xuser_8_reg[31:0];
   assign rd_resp_desc_2_xuser_9_xuser_f = rd_resp_desc_2_xuser_9_reg[31:0];
   assign rd_resp_desc_2_xuser_10_xuser_f = rd_resp_desc_2_xuser_10_reg[31:0];
   assign rd_resp_desc_2_xuser_11_xuser_f = rd_resp_desc_2_xuser_11_reg[31:0];
   assign rd_resp_desc_2_xuser_12_xuser_f = rd_resp_desc_2_xuser_12_reg[31:0];
   assign rd_resp_desc_2_xuser_13_xuser_f = rd_resp_desc_2_xuser_13_reg[31:0];
   assign rd_resp_desc_2_xuser_14_xuser_f = rd_resp_desc_2_xuser_14_reg[31:0];
   assign rd_resp_desc_2_xuser_15_xuser_f = rd_resp_desc_2_xuser_15_reg[31:0];
   assign wr_req_desc_2_txn_type_wr_strb_f = wr_req_desc_2_txn_type_reg[1];
   assign wr_req_desc_2_size_txn_size_f = wr_req_desc_2_size_reg[31:0];
   assign wr_req_desc_2_data_offset_addr_f = wr_req_desc_2_data_offset_reg[13:0];
   assign wr_req_desc_2_data_host_addr_0_addr_f = wr_req_desc_2_data_host_addr_0_reg[31:0];
   assign wr_req_desc_2_data_host_addr_1_addr_f = wr_req_desc_2_data_host_addr_1_reg[31:0];
   assign wr_req_desc_2_data_host_addr_2_addr_f = wr_req_desc_2_data_host_addr_2_reg[31:0];
   assign wr_req_desc_2_data_host_addr_3_addr_f = wr_req_desc_2_data_host_addr_3_reg[31:0];
   assign wr_req_desc_2_wstrb_host_addr_0_addr_f = wr_req_desc_2_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_2_wstrb_host_addr_1_addr_f = wr_req_desc_2_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_2_wstrb_host_addr_2_addr_f = wr_req_desc_2_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_2_wstrb_host_addr_3_addr_f = wr_req_desc_2_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_2_axsize_axsize_f = wr_req_desc_2_axsize_reg[2:0];
   assign wr_req_desc_2_attr_axsnoop_f = wr_req_desc_2_attr_reg[27:24];
   assign wr_req_desc_2_attr_axdomain_f = wr_req_desc_2_attr_reg[23:22];
   assign wr_req_desc_2_attr_axbar_f = wr_req_desc_2_attr_reg[21:20];
   assign wr_req_desc_2_attr_awunique_f = wr_req_desc_2_attr_reg[19];
   assign wr_req_desc_2_attr_axregion_f = wr_req_desc_2_attr_reg[18:15];
   assign wr_req_desc_2_attr_axqos_f = wr_req_desc_2_attr_reg[14:11];
   assign wr_req_desc_2_attr_axprot_f = wr_req_desc_2_attr_reg[10:8];
   assign wr_req_desc_2_attr_axcache_f = wr_req_desc_2_attr_reg[7:4];
   assign wr_req_desc_2_attr_axlock_f = wr_req_desc_2_attr_reg[2];
   assign wr_req_desc_2_attr_axburst_f = wr_req_desc_2_attr_reg[1:0];
   assign wr_req_desc_2_axaddr_0_addr_f = wr_req_desc_2_axaddr_0_reg[31:0];
   assign wr_req_desc_2_axaddr_1_addr_f = wr_req_desc_2_axaddr_1_reg[31:0];
   assign wr_req_desc_2_axaddr_2_addr_f = wr_req_desc_2_axaddr_2_reg[31:0];
   assign wr_req_desc_2_axaddr_3_addr_f = wr_req_desc_2_axaddr_3_reg[31:0];
   assign wr_req_desc_2_axid_0_axid_f = wr_req_desc_2_axid_0_reg[31:0];
   assign wr_req_desc_2_axid_1_axid_f = wr_req_desc_2_axid_1_reg[31:0];
   assign wr_req_desc_2_axid_2_axid_f = wr_req_desc_2_axid_2_reg[31:0];
   assign wr_req_desc_2_axid_3_axid_f = wr_req_desc_2_axid_3_reg[31:0];
   assign wr_req_desc_2_axuser_0_axuser_f = wr_req_desc_2_axuser_0_reg[31:0];
   assign wr_req_desc_2_axuser_1_axuser_f = wr_req_desc_2_axuser_1_reg[31:0];
   assign wr_req_desc_2_axuser_2_axuser_f = wr_req_desc_2_axuser_2_reg[31:0];
   assign wr_req_desc_2_axuser_3_axuser_f = wr_req_desc_2_axuser_3_reg[31:0];
   assign wr_req_desc_2_axuser_4_axuser_f = wr_req_desc_2_axuser_4_reg[31:0];
   assign wr_req_desc_2_axuser_5_axuser_f = wr_req_desc_2_axuser_5_reg[31:0];
   assign wr_req_desc_2_axuser_6_axuser_f = wr_req_desc_2_axuser_6_reg[31:0];
   assign wr_req_desc_2_axuser_7_axuser_f = wr_req_desc_2_axuser_7_reg[31:0];
   assign wr_req_desc_2_axuser_8_axuser_f = wr_req_desc_2_axuser_8_reg[31:0];
   assign wr_req_desc_2_axuser_9_axuser_f = wr_req_desc_2_axuser_9_reg[31:0];
   assign wr_req_desc_2_axuser_10_axuser_f = wr_req_desc_2_axuser_10_reg[31:0];
   assign wr_req_desc_2_axuser_11_axuser_f = wr_req_desc_2_axuser_11_reg[31:0];
   assign wr_req_desc_2_axuser_12_axuser_f = wr_req_desc_2_axuser_12_reg[31:0];
   assign wr_req_desc_2_axuser_13_axuser_f = wr_req_desc_2_axuser_13_reg[31:0];
   assign wr_req_desc_2_axuser_14_axuser_f = wr_req_desc_2_axuser_14_reg[31:0];
   assign wr_req_desc_2_axuser_15_axuser_f = wr_req_desc_2_axuser_15_reg[31:0];
   assign wr_req_desc_2_wuser_0_wuser_f = wr_req_desc_2_wuser_0_reg[31:0];
   assign wr_req_desc_2_wuser_1_wuser_f = wr_req_desc_2_wuser_1_reg[31:0];
   assign wr_req_desc_2_wuser_2_wuser_f = wr_req_desc_2_wuser_2_reg[31:0];
   assign wr_req_desc_2_wuser_3_wuser_f = wr_req_desc_2_wuser_3_reg[31:0];
   assign wr_req_desc_2_wuser_4_wuser_f = wr_req_desc_2_wuser_4_reg[31:0];
   assign wr_req_desc_2_wuser_5_wuser_f = wr_req_desc_2_wuser_5_reg[31:0];
   assign wr_req_desc_2_wuser_6_wuser_f = wr_req_desc_2_wuser_6_reg[31:0];
   assign wr_req_desc_2_wuser_7_wuser_f = wr_req_desc_2_wuser_7_reg[31:0];
   assign wr_req_desc_2_wuser_8_wuser_f = wr_req_desc_2_wuser_8_reg[31:0];
   assign wr_req_desc_2_wuser_9_wuser_f = wr_req_desc_2_wuser_9_reg[31:0];
   assign wr_req_desc_2_wuser_10_wuser_f = wr_req_desc_2_wuser_10_reg[31:0];
   assign wr_req_desc_2_wuser_11_wuser_f = wr_req_desc_2_wuser_11_reg[31:0];
   assign wr_req_desc_2_wuser_12_wuser_f = wr_req_desc_2_wuser_12_reg[31:0];
   assign wr_req_desc_2_wuser_13_wuser_f = wr_req_desc_2_wuser_13_reg[31:0];
   assign wr_req_desc_2_wuser_14_wuser_f = wr_req_desc_2_wuser_14_reg[31:0];
   assign wr_req_desc_2_wuser_15_wuser_f = wr_req_desc_2_wuser_15_reg[31:0];
   assign wr_resp_desc_2_resp_resp_f = wr_resp_desc_2_resp_reg[4:0];
   assign wr_resp_desc_2_xid_0_xid_f = wr_resp_desc_2_xid_0_reg[31:0];
   assign wr_resp_desc_2_xid_1_xid_f = wr_resp_desc_2_xid_1_reg[31:0];
   assign wr_resp_desc_2_xid_2_xid_f = wr_resp_desc_2_xid_2_reg[31:0];
   assign wr_resp_desc_2_xid_3_xid_f = wr_resp_desc_2_xid_3_reg[31:0];
   assign wr_resp_desc_2_xuser_0_xuser_f = wr_resp_desc_2_xuser_0_reg[31:0];
   assign wr_resp_desc_2_xuser_1_xuser_f = wr_resp_desc_2_xuser_1_reg[31:0];
   assign wr_resp_desc_2_xuser_2_xuser_f = wr_resp_desc_2_xuser_2_reg[31:0];
   assign wr_resp_desc_2_xuser_3_xuser_f = wr_resp_desc_2_xuser_3_reg[31:0];
   assign wr_resp_desc_2_xuser_4_xuser_f = wr_resp_desc_2_xuser_4_reg[31:0];
   assign wr_resp_desc_2_xuser_5_xuser_f = wr_resp_desc_2_xuser_5_reg[31:0];
   assign wr_resp_desc_2_xuser_6_xuser_f = wr_resp_desc_2_xuser_6_reg[31:0];
   assign wr_resp_desc_2_xuser_7_xuser_f = wr_resp_desc_2_xuser_7_reg[31:0];
   assign wr_resp_desc_2_xuser_8_xuser_f = wr_resp_desc_2_xuser_8_reg[31:0];
   assign wr_resp_desc_2_xuser_9_xuser_f = wr_resp_desc_2_xuser_9_reg[31:0];
   assign wr_resp_desc_2_xuser_10_xuser_f = wr_resp_desc_2_xuser_10_reg[31:0];
   assign wr_resp_desc_2_xuser_11_xuser_f = wr_resp_desc_2_xuser_11_reg[31:0];
   assign wr_resp_desc_2_xuser_12_xuser_f = wr_resp_desc_2_xuser_12_reg[31:0];
   assign wr_resp_desc_2_xuser_13_xuser_f = wr_resp_desc_2_xuser_13_reg[31:0];
   assign wr_resp_desc_2_xuser_14_xuser_f = wr_resp_desc_2_xuser_14_reg[31:0];
   assign wr_resp_desc_2_xuser_15_xuser_f = wr_resp_desc_2_xuser_15_reg[31:0];
   assign sn_req_desc_2_attr_acsnoop_f = sn_req_desc_2_attr_reg[27:24];
   assign sn_req_desc_2_attr_acprot_f = sn_req_desc_2_attr_reg[10:8];
   assign sn_req_desc_2_acaddr_0_addr_f = sn_req_desc_2_acaddr_0_reg[31:0];
   assign sn_req_desc_2_acaddr_1_addr_f = sn_req_desc_2_acaddr_1_reg[31:0];
   assign sn_req_desc_2_acaddr_2_addr_f = sn_req_desc_2_acaddr_2_reg[31:0];
   assign sn_req_desc_2_acaddr_3_addr_f = sn_req_desc_2_acaddr_3_reg[31:0];
   assign sn_resp_desc_2_resp_resp_f = sn_resp_desc_2_resp_reg[4:0];
   assign rd_req_desc_3_size_txn_size_f = rd_req_desc_3_size_reg[31:0];
   assign rd_req_desc_3_axsize_axsize_f = rd_req_desc_3_axsize_reg[2:0];
   assign rd_req_desc_3_attr_axsnoop_f = rd_req_desc_3_attr_reg[27:24];
   assign rd_req_desc_3_attr_axdomain_f = rd_req_desc_3_attr_reg[23:22];
   assign rd_req_desc_3_attr_axbar_f = rd_req_desc_3_attr_reg[21:20];
   assign rd_req_desc_3_attr_axregion_f = rd_req_desc_3_attr_reg[18:15];
   assign rd_req_desc_3_attr_axqos_f = rd_req_desc_3_attr_reg[14:11];
   assign rd_req_desc_3_attr_axprot_f = rd_req_desc_3_attr_reg[10:8];
   assign rd_req_desc_3_attr_axcache_f = rd_req_desc_3_attr_reg[7:4];
   assign rd_req_desc_3_attr_axlock_f = rd_req_desc_3_attr_reg[2];
   assign rd_req_desc_3_attr_axburst_f = rd_req_desc_3_attr_reg[1:0];
   assign rd_req_desc_3_axaddr_0_addr_f = rd_req_desc_3_axaddr_0_reg[31:0];
   assign rd_req_desc_3_axaddr_1_addr_f = rd_req_desc_3_axaddr_1_reg[31:0];
   assign rd_req_desc_3_axaddr_2_addr_f = rd_req_desc_3_axaddr_2_reg[31:0];
   assign rd_req_desc_3_axaddr_3_addr_f = rd_req_desc_3_axaddr_3_reg[31:0];
   assign rd_req_desc_3_axid_0_axid_f = rd_req_desc_3_axid_0_reg[31:0];
   assign rd_req_desc_3_axid_1_axid_f = rd_req_desc_3_axid_1_reg[31:0];
   assign rd_req_desc_3_axid_2_axid_f = rd_req_desc_3_axid_2_reg[31:0];
   assign rd_req_desc_3_axid_3_axid_f = rd_req_desc_3_axid_3_reg[31:0];
   assign rd_req_desc_3_axuser_0_axuser_f = rd_req_desc_3_axuser_0_reg[31:0];
   assign rd_req_desc_3_axuser_1_axuser_f = rd_req_desc_3_axuser_1_reg[31:0];
   assign rd_req_desc_3_axuser_2_axuser_f = rd_req_desc_3_axuser_2_reg[31:0];
   assign rd_req_desc_3_axuser_3_axuser_f = rd_req_desc_3_axuser_3_reg[31:0];
   assign rd_req_desc_3_axuser_4_axuser_f = rd_req_desc_3_axuser_4_reg[31:0];
   assign rd_req_desc_3_axuser_5_axuser_f = rd_req_desc_3_axuser_5_reg[31:0];
   assign rd_req_desc_3_axuser_6_axuser_f = rd_req_desc_3_axuser_6_reg[31:0];
   assign rd_req_desc_3_axuser_7_axuser_f = rd_req_desc_3_axuser_7_reg[31:0];
   assign rd_req_desc_3_axuser_8_axuser_f = rd_req_desc_3_axuser_8_reg[31:0];
   assign rd_req_desc_3_axuser_9_axuser_f = rd_req_desc_3_axuser_9_reg[31:0];
   assign rd_req_desc_3_axuser_10_axuser_f = rd_req_desc_3_axuser_10_reg[31:0];
   assign rd_req_desc_3_axuser_11_axuser_f = rd_req_desc_3_axuser_11_reg[31:0];
   assign rd_req_desc_3_axuser_12_axuser_f = rd_req_desc_3_axuser_12_reg[31:0];
   assign rd_req_desc_3_axuser_13_axuser_f = rd_req_desc_3_axuser_13_reg[31:0];
   assign rd_req_desc_3_axuser_14_axuser_f = rd_req_desc_3_axuser_14_reg[31:0];
   assign rd_req_desc_3_axuser_15_axuser_f = rd_req_desc_3_axuser_15_reg[31:0];
   assign rd_resp_desc_3_data_offset_addr_f = rd_resp_desc_3_data_offset_reg[13:0];
   assign rd_resp_desc_3_data_size_size_f = rd_resp_desc_3_data_size_reg[31:0];
   assign rd_resp_desc_3_data_host_addr_0_addr_f = rd_resp_desc_3_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_3_data_host_addr_1_addr_f = rd_resp_desc_3_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_3_data_host_addr_2_addr_f = rd_resp_desc_3_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_3_data_host_addr_3_addr_f = rd_resp_desc_3_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_3_resp_resp_f = rd_resp_desc_3_resp_reg[4:0];
   assign rd_resp_desc_3_xid_0_xid_f = rd_resp_desc_3_xid_0_reg[31:0];
   assign rd_resp_desc_3_xid_1_xid_f = rd_resp_desc_3_xid_1_reg[31:0];
   assign rd_resp_desc_3_xid_2_xid_f = rd_resp_desc_3_xid_2_reg[31:0];
   assign rd_resp_desc_3_xid_3_xid_f = rd_resp_desc_3_xid_3_reg[31:0];
   assign rd_resp_desc_3_xuser_0_xuser_f = rd_resp_desc_3_xuser_0_reg[31:0];
   assign rd_resp_desc_3_xuser_1_xuser_f = rd_resp_desc_3_xuser_1_reg[31:0];
   assign rd_resp_desc_3_xuser_2_xuser_f = rd_resp_desc_3_xuser_2_reg[31:0];
   assign rd_resp_desc_3_xuser_3_xuser_f = rd_resp_desc_3_xuser_3_reg[31:0];
   assign rd_resp_desc_3_xuser_4_xuser_f = rd_resp_desc_3_xuser_4_reg[31:0];
   assign rd_resp_desc_3_xuser_5_xuser_f = rd_resp_desc_3_xuser_5_reg[31:0];
   assign rd_resp_desc_3_xuser_6_xuser_f = rd_resp_desc_3_xuser_6_reg[31:0];
   assign rd_resp_desc_3_xuser_7_xuser_f = rd_resp_desc_3_xuser_7_reg[31:0];
   assign rd_resp_desc_3_xuser_8_xuser_f = rd_resp_desc_3_xuser_8_reg[31:0];
   assign rd_resp_desc_3_xuser_9_xuser_f = rd_resp_desc_3_xuser_9_reg[31:0];
   assign rd_resp_desc_3_xuser_10_xuser_f = rd_resp_desc_3_xuser_10_reg[31:0];
   assign rd_resp_desc_3_xuser_11_xuser_f = rd_resp_desc_3_xuser_11_reg[31:0];
   assign rd_resp_desc_3_xuser_12_xuser_f = rd_resp_desc_3_xuser_12_reg[31:0];
   assign rd_resp_desc_3_xuser_13_xuser_f = rd_resp_desc_3_xuser_13_reg[31:0];
   assign rd_resp_desc_3_xuser_14_xuser_f = rd_resp_desc_3_xuser_14_reg[31:0];
   assign rd_resp_desc_3_xuser_15_xuser_f = rd_resp_desc_3_xuser_15_reg[31:0];
   assign wr_req_desc_3_txn_type_wr_strb_f = wr_req_desc_3_txn_type_reg[1];
   assign wr_req_desc_3_size_txn_size_f = wr_req_desc_3_size_reg[31:0];
   assign wr_req_desc_3_data_offset_addr_f = wr_req_desc_3_data_offset_reg[13:0];
   assign wr_req_desc_3_data_host_addr_0_addr_f = wr_req_desc_3_data_host_addr_0_reg[31:0];
   assign wr_req_desc_3_data_host_addr_1_addr_f = wr_req_desc_3_data_host_addr_1_reg[31:0];
   assign wr_req_desc_3_data_host_addr_2_addr_f = wr_req_desc_3_data_host_addr_2_reg[31:0];
   assign wr_req_desc_3_data_host_addr_3_addr_f = wr_req_desc_3_data_host_addr_3_reg[31:0];
   assign wr_req_desc_3_wstrb_host_addr_0_addr_f = wr_req_desc_3_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_3_wstrb_host_addr_1_addr_f = wr_req_desc_3_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_3_wstrb_host_addr_2_addr_f = wr_req_desc_3_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_3_wstrb_host_addr_3_addr_f = wr_req_desc_3_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_3_axsize_axsize_f = wr_req_desc_3_axsize_reg[2:0];
   assign wr_req_desc_3_attr_axsnoop_f = wr_req_desc_3_attr_reg[27:24];
   assign wr_req_desc_3_attr_axdomain_f = wr_req_desc_3_attr_reg[23:22];
   assign wr_req_desc_3_attr_axbar_f = wr_req_desc_3_attr_reg[21:20];
   assign wr_req_desc_3_attr_awunique_f = wr_req_desc_3_attr_reg[19];
   assign wr_req_desc_3_attr_axregion_f = wr_req_desc_3_attr_reg[18:15];
   assign wr_req_desc_3_attr_axqos_f = wr_req_desc_3_attr_reg[14:11];
   assign wr_req_desc_3_attr_axprot_f = wr_req_desc_3_attr_reg[10:8];
   assign wr_req_desc_3_attr_axcache_f = wr_req_desc_3_attr_reg[7:4];
   assign wr_req_desc_3_attr_axlock_f = wr_req_desc_3_attr_reg[2];
   assign wr_req_desc_3_attr_axburst_f = wr_req_desc_3_attr_reg[1:0];
   assign wr_req_desc_3_axaddr_0_addr_f = wr_req_desc_3_axaddr_0_reg[31:0];
   assign wr_req_desc_3_axaddr_1_addr_f = wr_req_desc_3_axaddr_1_reg[31:0];
   assign wr_req_desc_3_axaddr_2_addr_f = wr_req_desc_3_axaddr_2_reg[31:0];
   assign wr_req_desc_3_axaddr_3_addr_f = wr_req_desc_3_axaddr_3_reg[31:0];
   assign wr_req_desc_3_axid_0_axid_f = wr_req_desc_3_axid_0_reg[31:0];
   assign wr_req_desc_3_axid_1_axid_f = wr_req_desc_3_axid_1_reg[31:0];
   assign wr_req_desc_3_axid_2_axid_f = wr_req_desc_3_axid_2_reg[31:0];
   assign wr_req_desc_3_axid_3_axid_f = wr_req_desc_3_axid_3_reg[31:0];
   assign wr_req_desc_3_axuser_0_axuser_f = wr_req_desc_3_axuser_0_reg[31:0];
   assign wr_req_desc_3_axuser_1_axuser_f = wr_req_desc_3_axuser_1_reg[31:0];
   assign wr_req_desc_3_axuser_2_axuser_f = wr_req_desc_3_axuser_2_reg[31:0];
   assign wr_req_desc_3_axuser_3_axuser_f = wr_req_desc_3_axuser_3_reg[31:0];
   assign wr_req_desc_3_axuser_4_axuser_f = wr_req_desc_3_axuser_4_reg[31:0];
   assign wr_req_desc_3_axuser_5_axuser_f = wr_req_desc_3_axuser_5_reg[31:0];
   assign wr_req_desc_3_axuser_6_axuser_f = wr_req_desc_3_axuser_6_reg[31:0];
   assign wr_req_desc_3_axuser_7_axuser_f = wr_req_desc_3_axuser_7_reg[31:0];
   assign wr_req_desc_3_axuser_8_axuser_f = wr_req_desc_3_axuser_8_reg[31:0];
   assign wr_req_desc_3_axuser_9_axuser_f = wr_req_desc_3_axuser_9_reg[31:0];
   assign wr_req_desc_3_axuser_10_axuser_f = wr_req_desc_3_axuser_10_reg[31:0];
   assign wr_req_desc_3_axuser_11_axuser_f = wr_req_desc_3_axuser_11_reg[31:0];
   assign wr_req_desc_3_axuser_12_axuser_f = wr_req_desc_3_axuser_12_reg[31:0];
   assign wr_req_desc_3_axuser_13_axuser_f = wr_req_desc_3_axuser_13_reg[31:0];
   assign wr_req_desc_3_axuser_14_axuser_f = wr_req_desc_3_axuser_14_reg[31:0];
   assign wr_req_desc_3_axuser_15_axuser_f = wr_req_desc_3_axuser_15_reg[31:0];
   assign wr_req_desc_3_wuser_0_wuser_f = wr_req_desc_3_wuser_0_reg[31:0];
   assign wr_req_desc_3_wuser_1_wuser_f = wr_req_desc_3_wuser_1_reg[31:0];
   assign wr_req_desc_3_wuser_2_wuser_f = wr_req_desc_3_wuser_2_reg[31:0];
   assign wr_req_desc_3_wuser_3_wuser_f = wr_req_desc_3_wuser_3_reg[31:0];
   assign wr_req_desc_3_wuser_4_wuser_f = wr_req_desc_3_wuser_4_reg[31:0];
   assign wr_req_desc_3_wuser_5_wuser_f = wr_req_desc_3_wuser_5_reg[31:0];
   assign wr_req_desc_3_wuser_6_wuser_f = wr_req_desc_3_wuser_6_reg[31:0];
   assign wr_req_desc_3_wuser_7_wuser_f = wr_req_desc_3_wuser_7_reg[31:0];
   assign wr_req_desc_3_wuser_8_wuser_f = wr_req_desc_3_wuser_8_reg[31:0];
   assign wr_req_desc_3_wuser_9_wuser_f = wr_req_desc_3_wuser_9_reg[31:0];
   assign wr_req_desc_3_wuser_10_wuser_f = wr_req_desc_3_wuser_10_reg[31:0];
   assign wr_req_desc_3_wuser_11_wuser_f = wr_req_desc_3_wuser_11_reg[31:0];
   assign wr_req_desc_3_wuser_12_wuser_f = wr_req_desc_3_wuser_12_reg[31:0];
   assign wr_req_desc_3_wuser_13_wuser_f = wr_req_desc_3_wuser_13_reg[31:0];
   assign wr_req_desc_3_wuser_14_wuser_f = wr_req_desc_3_wuser_14_reg[31:0];
   assign wr_req_desc_3_wuser_15_wuser_f = wr_req_desc_3_wuser_15_reg[31:0];
   assign wr_resp_desc_3_resp_resp_f = wr_resp_desc_3_resp_reg[4:0];
   assign wr_resp_desc_3_xid_0_xid_f = wr_resp_desc_3_xid_0_reg[31:0];
   assign wr_resp_desc_3_xid_1_xid_f = wr_resp_desc_3_xid_1_reg[31:0];
   assign wr_resp_desc_3_xid_2_xid_f = wr_resp_desc_3_xid_2_reg[31:0];
   assign wr_resp_desc_3_xid_3_xid_f = wr_resp_desc_3_xid_3_reg[31:0];
   assign wr_resp_desc_3_xuser_0_xuser_f = wr_resp_desc_3_xuser_0_reg[31:0];
   assign wr_resp_desc_3_xuser_1_xuser_f = wr_resp_desc_3_xuser_1_reg[31:0];
   assign wr_resp_desc_3_xuser_2_xuser_f = wr_resp_desc_3_xuser_2_reg[31:0];
   assign wr_resp_desc_3_xuser_3_xuser_f = wr_resp_desc_3_xuser_3_reg[31:0];
   assign wr_resp_desc_3_xuser_4_xuser_f = wr_resp_desc_3_xuser_4_reg[31:0];
   assign wr_resp_desc_3_xuser_5_xuser_f = wr_resp_desc_3_xuser_5_reg[31:0];
   assign wr_resp_desc_3_xuser_6_xuser_f = wr_resp_desc_3_xuser_6_reg[31:0];
   assign wr_resp_desc_3_xuser_7_xuser_f = wr_resp_desc_3_xuser_7_reg[31:0];
   assign wr_resp_desc_3_xuser_8_xuser_f = wr_resp_desc_3_xuser_8_reg[31:0];
   assign wr_resp_desc_3_xuser_9_xuser_f = wr_resp_desc_3_xuser_9_reg[31:0];
   assign wr_resp_desc_3_xuser_10_xuser_f = wr_resp_desc_3_xuser_10_reg[31:0];
   assign wr_resp_desc_3_xuser_11_xuser_f = wr_resp_desc_3_xuser_11_reg[31:0];
   assign wr_resp_desc_3_xuser_12_xuser_f = wr_resp_desc_3_xuser_12_reg[31:0];
   assign wr_resp_desc_3_xuser_13_xuser_f = wr_resp_desc_3_xuser_13_reg[31:0];
   assign wr_resp_desc_3_xuser_14_xuser_f = wr_resp_desc_3_xuser_14_reg[31:0];
   assign wr_resp_desc_3_xuser_15_xuser_f = wr_resp_desc_3_xuser_15_reg[31:0];
   assign sn_req_desc_3_attr_acsnoop_f = sn_req_desc_3_attr_reg[27:24];
   assign sn_req_desc_3_attr_acprot_f = sn_req_desc_3_attr_reg[10:8];
   assign sn_req_desc_3_acaddr_0_addr_f = sn_req_desc_3_acaddr_0_reg[31:0];
   assign sn_req_desc_3_acaddr_1_addr_f = sn_req_desc_3_acaddr_1_reg[31:0];
   assign sn_req_desc_3_acaddr_2_addr_f = sn_req_desc_3_acaddr_2_reg[31:0];
   assign sn_req_desc_3_acaddr_3_addr_f = sn_req_desc_3_acaddr_3_reg[31:0];
   assign sn_resp_desc_3_resp_resp_f = sn_resp_desc_3_resp_reg[4:0];
   assign rd_req_desc_4_size_txn_size_f = rd_req_desc_4_size_reg[31:0];
   assign rd_req_desc_4_axsize_axsize_f = rd_req_desc_4_axsize_reg[2:0];
   assign rd_req_desc_4_attr_axsnoop_f = rd_req_desc_4_attr_reg[27:24];
   assign rd_req_desc_4_attr_axdomain_f = rd_req_desc_4_attr_reg[23:22];
   assign rd_req_desc_4_attr_axbar_f = rd_req_desc_4_attr_reg[21:20];
   assign rd_req_desc_4_attr_axregion_f = rd_req_desc_4_attr_reg[18:15];
   assign rd_req_desc_4_attr_axqos_f = rd_req_desc_4_attr_reg[14:11];
   assign rd_req_desc_4_attr_axprot_f = rd_req_desc_4_attr_reg[10:8];
   assign rd_req_desc_4_attr_axcache_f = rd_req_desc_4_attr_reg[7:4];
   assign rd_req_desc_4_attr_axlock_f = rd_req_desc_4_attr_reg[2];
   assign rd_req_desc_4_attr_axburst_f = rd_req_desc_4_attr_reg[1:0];
   assign rd_req_desc_4_axaddr_0_addr_f = rd_req_desc_4_axaddr_0_reg[31:0];
   assign rd_req_desc_4_axaddr_1_addr_f = rd_req_desc_4_axaddr_1_reg[31:0];
   assign rd_req_desc_4_axaddr_2_addr_f = rd_req_desc_4_axaddr_2_reg[31:0];
   assign rd_req_desc_4_axaddr_3_addr_f = rd_req_desc_4_axaddr_3_reg[31:0];
   assign rd_req_desc_4_axid_0_axid_f = rd_req_desc_4_axid_0_reg[31:0];
   assign rd_req_desc_4_axid_1_axid_f = rd_req_desc_4_axid_1_reg[31:0];
   assign rd_req_desc_4_axid_2_axid_f = rd_req_desc_4_axid_2_reg[31:0];
   assign rd_req_desc_4_axid_3_axid_f = rd_req_desc_4_axid_3_reg[31:0];
   assign rd_req_desc_4_axuser_0_axuser_f = rd_req_desc_4_axuser_0_reg[31:0];
   assign rd_req_desc_4_axuser_1_axuser_f = rd_req_desc_4_axuser_1_reg[31:0];
   assign rd_req_desc_4_axuser_2_axuser_f = rd_req_desc_4_axuser_2_reg[31:0];
   assign rd_req_desc_4_axuser_3_axuser_f = rd_req_desc_4_axuser_3_reg[31:0];
   assign rd_req_desc_4_axuser_4_axuser_f = rd_req_desc_4_axuser_4_reg[31:0];
   assign rd_req_desc_4_axuser_5_axuser_f = rd_req_desc_4_axuser_5_reg[31:0];
   assign rd_req_desc_4_axuser_6_axuser_f = rd_req_desc_4_axuser_6_reg[31:0];
   assign rd_req_desc_4_axuser_7_axuser_f = rd_req_desc_4_axuser_7_reg[31:0];
   assign rd_req_desc_4_axuser_8_axuser_f = rd_req_desc_4_axuser_8_reg[31:0];
   assign rd_req_desc_4_axuser_9_axuser_f = rd_req_desc_4_axuser_9_reg[31:0];
   assign rd_req_desc_4_axuser_10_axuser_f = rd_req_desc_4_axuser_10_reg[31:0];
   assign rd_req_desc_4_axuser_11_axuser_f = rd_req_desc_4_axuser_11_reg[31:0];
   assign rd_req_desc_4_axuser_12_axuser_f = rd_req_desc_4_axuser_12_reg[31:0];
   assign rd_req_desc_4_axuser_13_axuser_f = rd_req_desc_4_axuser_13_reg[31:0];
   assign rd_req_desc_4_axuser_14_axuser_f = rd_req_desc_4_axuser_14_reg[31:0];
   assign rd_req_desc_4_axuser_15_axuser_f = rd_req_desc_4_axuser_15_reg[31:0];
   assign rd_resp_desc_4_data_offset_addr_f = rd_resp_desc_4_data_offset_reg[13:0];
   assign rd_resp_desc_4_data_size_size_f = rd_resp_desc_4_data_size_reg[31:0];
   assign rd_resp_desc_4_data_host_addr_0_addr_f = rd_resp_desc_4_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_4_data_host_addr_1_addr_f = rd_resp_desc_4_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_4_data_host_addr_2_addr_f = rd_resp_desc_4_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_4_data_host_addr_3_addr_f = rd_resp_desc_4_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_4_resp_resp_f = rd_resp_desc_4_resp_reg[4:0];
   assign rd_resp_desc_4_xid_0_xid_f = rd_resp_desc_4_xid_0_reg[31:0];
   assign rd_resp_desc_4_xid_1_xid_f = rd_resp_desc_4_xid_1_reg[31:0];
   assign rd_resp_desc_4_xid_2_xid_f = rd_resp_desc_4_xid_2_reg[31:0];
   assign rd_resp_desc_4_xid_3_xid_f = rd_resp_desc_4_xid_3_reg[31:0];
   assign rd_resp_desc_4_xuser_0_xuser_f = rd_resp_desc_4_xuser_0_reg[31:0];
   assign rd_resp_desc_4_xuser_1_xuser_f = rd_resp_desc_4_xuser_1_reg[31:0];
   assign rd_resp_desc_4_xuser_2_xuser_f = rd_resp_desc_4_xuser_2_reg[31:0];
   assign rd_resp_desc_4_xuser_3_xuser_f = rd_resp_desc_4_xuser_3_reg[31:0];
   assign rd_resp_desc_4_xuser_4_xuser_f = rd_resp_desc_4_xuser_4_reg[31:0];
   assign rd_resp_desc_4_xuser_5_xuser_f = rd_resp_desc_4_xuser_5_reg[31:0];
   assign rd_resp_desc_4_xuser_6_xuser_f = rd_resp_desc_4_xuser_6_reg[31:0];
   assign rd_resp_desc_4_xuser_7_xuser_f = rd_resp_desc_4_xuser_7_reg[31:0];
   assign rd_resp_desc_4_xuser_8_xuser_f = rd_resp_desc_4_xuser_8_reg[31:0];
   assign rd_resp_desc_4_xuser_9_xuser_f = rd_resp_desc_4_xuser_9_reg[31:0];
   assign rd_resp_desc_4_xuser_10_xuser_f = rd_resp_desc_4_xuser_10_reg[31:0];
   assign rd_resp_desc_4_xuser_11_xuser_f = rd_resp_desc_4_xuser_11_reg[31:0];
   assign rd_resp_desc_4_xuser_12_xuser_f = rd_resp_desc_4_xuser_12_reg[31:0];
   assign rd_resp_desc_4_xuser_13_xuser_f = rd_resp_desc_4_xuser_13_reg[31:0];
   assign rd_resp_desc_4_xuser_14_xuser_f = rd_resp_desc_4_xuser_14_reg[31:0];
   assign rd_resp_desc_4_xuser_15_xuser_f = rd_resp_desc_4_xuser_15_reg[31:0];
   assign wr_req_desc_4_txn_type_wr_strb_f = wr_req_desc_4_txn_type_reg[1];
   assign wr_req_desc_4_size_txn_size_f = wr_req_desc_4_size_reg[31:0];
   assign wr_req_desc_4_data_offset_addr_f = wr_req_desc_4_data_offset_reg[13:0];
   assign wr_req_desc_4_data_host_addr_0_addr_f = wr_req_desc_4_data_host_addr_0_reg[31:0];
   assign wr_req_desc_4_data_host_addr_1_addr_f = wr_req_desc_4_data_host_addr_1_reg[31:0];
   assign wr_req_desc_4_data_host_addr_2_addr_f = wr_req_desc_4_data_host_addr_2_reg[31:0];
   assign wr_req_desc_4_data_host_addr_3_addr_f = wr_req_desc_4_data_host_addr_3_reg[31:0];
   assign wr_req_desc_4_wstrb_host_addr_0_addr_f = wr_req_desc_4_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_4_wstrb_host_addr_1_addr_f = wr_req_desc_4_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_4_wstrb_host_addr_2_addr_f = wr_req_desc_4_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_4_wstrb_host_addr_3_addr_f = wr_req_desc_4_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_4_axsize_axsize_f = wr_req_desc_4_axsize_reg[2:0];
   assign wr_req_desc_4_attr_axsnoop_f = wr_req_desc_4_attr_reg[27:24];
   assign wr_req_desc_4_attr_axdomain_f = wr_req_desc_4_attr_reg[23:22];
   assign wr_req_desc_4_attr_axbar_f = wr_req_desc_4_attr_reg[21:20];
   assign wr_req_desc_4_attr_awunique_f = wr_req_desc_4_attr_reg[19];
   assign wr_req_desc_4_attr_axregion_f = wr_req_desc_4_attr_reg[18:15];
   assign wr_req_desc_4_attr_axqos_f = wr_req_desc_4_attr_reg[14:11];
   assign wr_req_desc_4_attr_axprot_f = wr_req_desc_4_attr_reg[10:8];
   assign wr_req_desc_4_attr_axcache_f = wr_req_desc_4_attr_reg[7:4];
   assign wr_req_desc_4_attr_axlock_f = wr_req_desc_4_attr_reg[2];
   assign wr_req_desc_4_attr_axburst_f = wr_req_desc_4_attr_reg[1:0];
   assign wr_req_desc_4_axaddr_0_addr_f = wr_req_desc_4_axaddr_0_reg[31:0];
   assign wr_req_desc_4_axaddr_1_addr_f = wr_req_desc_4_axaddr_1_reg[31:0];
   assign wr_req_desc_4_axaddr_2_addr_f = wr_req_desc_4_axaddr_2_reg[31:0];
   assign wr_req_desc_4_axaddr_3_addr_f = wr_req_desc_4_axaddr_3_reg[31:0];
   assign wr_req_desc_4_axid_0_axid_f = wr_req_desc_4_axid_0_reg[31:0];
   assign wr_req_desc_4_axid_1_axid_f = wr_req_desc_4_axid_1_reg[31:0];
   assign wr_req_desc_4_axid_2_axid_f = wr_req_desc_4_axid_2_reg[31:0];
   assign wr_req_desc_4_axid_3_axid_f = wr_req_desc_4_axid_3_reg[31:0];
   assign wr_req_desc_4_axuser_0_axuser_f = wr_req_desc_4_axuser_0_reg[31:0];
   assign wr_req_desc_4_axuser_1_axuser_f = wr_req_desc_4_axuser_1_reg[31:0];
   assign wr_req_desc_4_axuser_2_axuser_f = wr_req_desc_4_axuser_2_reg[31:0];
   assign wr_req_desc_4_axuser_3_axuser_f = wr_req_desc_4_axuser_3_reg[31:0];
   assign wr_req_desc_4_axuser_4_axuser_f = wr_req_desc_4_axuser_4_reg[31:0];
   assign wr_req_desc_4_axuser_5_axuser_f = wr_req_desc_4_axuser_5_reg[31:0];
   assign wr_req_desc_4_axuser_6_axuser_f = wr_req_desc_4_axuser_6_reg[31:0];
   assign wr_req_desc_4_axuser_7_axuser_f = wr_req_desc_4_axuser_7_reg[31:0];
   assign wr_req_desc_4_axuser_8_axuser_f = wr_req_desc_4_axuser_8_reg[31:0];
   assign wr_req_desc_4_axuser_9_axuser_f = wr_req_desc_4_axuser_9_reg[31:0];
   assign wr_req_desc_4_axuser_10_axuser_f = wr_req_desc_4_axuser_10_reg[31:0];
   assign wr_req_desc_4_axuser_11_axuser_f = wr_req_desc_4_axuser_11_reg[31:0];
   assign wr_req_desc_4_axuser_12_axuser_f = wr_req_desc_4_axuser_12_reg[31:0];
   assign wr_req_desc_4_axuser_13_axuser_f = wr_req_desc_4_axuser_13_reg[31:0];
   assign wr_req_desc_4_axuser_14_axuser_f = wr_req_desc_4_axuser_14_reg[31:0];
   assign wr_req_desc_4_axuser_15_axuser_f = wr_req_desc_4_axuser_15_reg[31:0];
   assign wr_req_desc_4_wuser_0_wuser_f = wr_req_desc_4_wuser_0_reg[31:0];
   assign wr_req_desc_4_wuser_1_wuser_f = wr_req_desc_4_wuser_1_reg[31:0];
   assign wr_req_desc_4_wuser_2_wuser_f = wr_req_desc_4_wuser_2_reg[31:0];
   assign wr_req_desc_4_wuser_3_wuser_f = wr_req_desc_4_wuser_3_reg[31:0];
   assign wr_req_desc_4_wuser_4_wuser_f = wr_req_desc_4_wuser_4_reg[31:0];
   assign wr_req_desc_4_wuser_5_wuser_f = wr_req_desc_4_wuser_5_reg[31:0];
   assign wr_req_desc_4_wuser_6_wuser_f = wr_req_desc_4_wuser_6_reg[31:0];
   assign wr_req_desc_4_wuser_7_wuser_f = wr_req_desc_4_wuser_7_reg[31:0];
   assign wr_req_desc_4_wuser_8_wuser_f = wr_req_desc_4_wuser_8_reg[31:0];
   assign wr_req_desc_4_wuser_9_wuser_f = wr_req_desc_4_wuser_9_reg[31:0];
   assign wr_req_desc_4_wuser_10_wuser_f = wr_req_desc_4_wuser_10_reg[31:0];
   assign wr_req_desc_4_wuser_11_wuser_f = wr_req_desc_4_wuser_11_reg[31:0];
   assign wr_req_desc_4_wuser_12_wuser_f = wr_req_desc_4_wuser_12_reg[31:0];
   assign wr_req_desc_4_wuser_13_wuser_f = wr_req_desc_4_wuser_13_reg[31:0];
   assign wr_req_desc_4_wuser_14_wuser_f = wr_req_desc_4_wuser_14_reg[31:0];
   assign wr_req_desc_4_wuser_15_wuser_f = wr_req_desc_4_wuser_15_reg[31:0];
   assign wr_resp_desc_4_resp_resp_f = wr_resp_desc_4_resp_reg[4:0];
   assign wr_resp_desc_4_xid_0_xid_f = wr_resp_desc_4_xid_0_reg[31:0];
   assign wr_resp_desc_4_xid_1_xid_f = wr_resp_desc_4_xid_1_reg[31:0];
   assign wr_resp_desc_4_xid_2_xid_f = wr_resp_desc_4_xid_2_reg[31:0];
   assign wr_resp_desc_4_xid_3_xid_f = wr_resp_desc_4_xid_3_reg[31:0];
   assign wr_resp_desc_4_xuser_0_xuser_f = wr_resp_desc_4_xuser_0_reg[31:0];
   assign wr_resp_desc_4_xuser_1_xuser_f = wr_resp_desc_4_xuser_1_reg[31:0];
   assign wr_resp_desc_4_xuser_2_xuser_f = wr_resp_desc_4_xuser_2_reg[31:0];
   assign wr_resp_desc_4_xuser_3_xuser_f = wr_resp_desc_4_xuser_3_reg[31:0];
   assign wr_resp_desc_4_xuser_4_xuser_f = wr_resp_desc_4_xuser_4_reg[31:0];
   assign wr_resp_desc_4_xuser_5_xuser_f = wr_resp_desc_4_xuser_5_reg[31:0];
   assign wr_resp_desc_4_xuser_6_xuser_f = wr_resp_desc_4_xuser_6_reg[31:0];
   assign wr_resp_desc_4_xuser_7_xuser_f = wr_resp_desc_4_xuser_7_reg[31:0];
   assign wr_resp_desc_4_xuser_8_xuser_f = wr_resp_desc_4_xuser_8_reg[31:0];
   assign wr_resp_desc_4_xuser_9_xuser_f = wr_resp_desc_4_xuser_9_reg[31:0];
   assign wr_resp_desc_4_xuser_10_xuser_f = wr_resp_desc_4_xuser_10_reg[31:0];
   assign wr_resp_desc_4_xuser_11_xuser_f = wr_resp_desc_4_xuser_11_reg[31:0];
   assign wr_resp_desc_4_xuser_12_xuser_f = wr_resp_desc_4_xuser_12_reg[31:0];
   assign wr_resp_desc_4_xuser_13_xuser_f = wr_resp_desc_4_xuser_13_reg[31:0];
   assign wr_resp_desc_4_xuser_14_xuser_f = wr_resp_desc_4_xuser_14_reg[31:0];
   assign wr_resp_desc_4_xuser_15_xuser_f = wr_resp_desc_4_xuser_15_reg[31:0];
   assign sn_req_desc_4_attr_acsnoop_f = sn_req_desc_4_attr_reg[27:24];
   assign sn_req_desc_4_attr_acprot_f = sn_req_desc_4_attr_reg[10:8];
   assign sn_req_desc_4_acaddr_0_addr_f = sn_req_desc_4_acaddr_0_reg[31:0];
   assign sn_req_desc_4_acaddr_1_addr_f = sn_req_desc_4_acaddr_1_reg[31:0];
   assign sn_req_desc_4_acaddr_2_addr_f = sn_req_desc_4_acaddr_2_reg[31:0];
   assign sn_req_desc_4_acaddr_3_addr_f = sn_req_desc_4_acaddr_3_reg[31:0];
   assign sn_resp_desc_4_resp_resp_f = sn_resp_desc_4_resp_reg[4:0];
   assign rd_req_desc_5_size_txn_size_f = rd_req_desc_5_size_reg[31:0];
   assign rd_req_desc_5_axsize_axsize_f = rd_req_desc_5_axsize_reg[2:0];
   assign rd_req_desc_5_attr_axsnoop_f = rd_req_desc_5_attr_reg[27:24];
   assign rd_req_desc_5_attr_axdomain_f = rd_req_desc_5_attr_reg[23:22];
   assign rd_req_desc_5_attr_axbar_f = rd_req_desc_5_attr_reg[21:20];
   assign rd_req_desc_5_attr_axregion_f = rd_req_desc_5_attr_reg[18:15];
   assign rd_req_desc_5_attr_axqos_f = rd_req_desc_5_attr_reg[14:11];
   assign rd_req_desc_5_attr_axprot_f = rd_req_desc_5_attr_reg[10:8];
   assign rd_req_desc_5_attr_axcache_f = rd_req_desc_5_attr_reg[7:4];
   assign rd_req_desc_5_attr_axlock_f = rd_req_desc_5_attr_reg[2];
   assign rd_req_desc_5_attr_axburst_f = rd_req_desc_5_attr_reg[1:0];
   assign rd_req_desc_5_axaddr_0_addr_f = rd_req_desc_5_axaddr_0_reg[31:0];
   assign rd_req_desc_5_axaddr_1_addr_f = rd_req_desc_5_axaddr_1_reg[31:0];
   assign rd_req_desc_5_axaddr_2_addr_f = rd_req_desc_5_axaddr_2_reg[31:0];
   assign rd_req_desc_5_axaddr_3_addr_f = rd_req_desc_5_axaddr_3_reg[31:0];
   assign rd_req_desc_5_axid_0_axid_f = rd_req_desc_5_axid_0_reg[31:0];
   assign rd_req_desc_5_axid_1_axid_f = rd_req_desc_5_axid_1_reg[31:0];
   assign rd_req_desc_5_axid_2_axid_f = rd_req_desc_5_axid_2_reg[31:0];
   assign rd_req_desc_5_axid_3_axid_f = rd_req_desc_5_axid_3_reg[31:0];
   assign rd_req_desc_5_axuser_0_axuser_f = rd_req_desc_5_axuser_0_reg[31:0];
   assign rd_req_desc_5_axuser_1_axuser_f = rd_req_desc_5_axuser_1_reg[31:0];
   assign rd_req_desc_5_axuser_2_axuser_f = rd_req_desc_5_axuser_2_reg[31:0];
   assign rd_req_desc_5_axuser_3_axuser_f = rd_req_desc_5_axuser_3_reg[31:0];
   assign rd_req_desc_5_axuser_4_axuser_f = rd_req_desc_5_axuser_4_reg[31:0];
   assign rd_req_desc_5_axuser_5_axuser_f = rd_req_desc_5_axuser_5_reg[31:0];
   assign rd_req_desc_5_axuser_6_axuser_f = rd_req_desc_5_axuser_6_reg[31:0];
   assign rd_req_desc_5_axuser_7_axuser_f = rd_req_desc_5_axuser_7_reg[31:0];
   assign rd_req_desc_5_axuser_8_axuser_f = rd_req_desc_5_axuser_8_reg[31:0];
   assign rd_req_desc_5_axuser_9_axuser_f = rd_req_desc_5_axuser_9_reg[31:0];
   assign rd_req_desc_5_axuser_10_axuser_f = rd_req_desc_5_axuser_10_reg[31:0];
   assign rd_req_desc_5_axuser_11_axuser_f = rd_req_desc_5_axuser_11_reg[31:0];
   assign rd_req_desc_5_axuser_12_axuser_f = rd_req_desc_5_axuser_12_reg[31:0];
   assign rd_req_desc_5_axuser_13_axuser_f = rd_req_desc_5_axuser_13_reg[31:0];
   assign rd_req_desc_5_axuser_14_axuser_f = rd_req_desc_5_axuser_14_reg[31:0];
   assign rd_req_desc_5_axuser_15_axuser_f = rd_req_desc_5_axuser_15_reg[31:0];
   assign rd_resp_desc_5_data_offset_addr_f = rd_resp_desc_5_data_offset_reg[13:0];
   assign rd_resp_desc_5_data_size_size_f = rd_resp_desc_5_data_size_reg[31:0];
   assign rd_resp_desc_5_data_host_addr_0_addr_f = rd_resp_desc_5_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_5_data_host_addr_1_addr_f = rd_resp_desc_5_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_5_data_host_addr_2_addr_f = rd_resp_desc_5_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_5_data_host_addr_3_addr_f = rd_resp_desc_5_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_5_resp_resp_f = rd_resp_desc_5_resp_reg[4:0];
   assign rd_resp_desc_5_xid_0_xid_f = rd_resp_desc_5_xid_0_reg[31:0];
   assign rd_resp_desc_5_xid_1_xid_f = rd_resp_desc_5_xid_1_reg[31:0];
   assign rd_resp_desc_5_xid_2_xid_f = rd_resp_desc_5_xid_2_reg[31:0];
   assign rd_resp_desc_5_xid_3_xid_f = rd_resp_desc_5_xid_3_reg[31:0];
   assign rd_resp_desc_5_xuser_0_xuser_f = rd_resp_desc_5_xuser_0_reg[31:0];
   assign rd_resp_desc_5_xuser_1_xuser_f = rd_resp_desc_5_xuser_1_reg[31:0];
   assign rd_resp_desc_5_xuser_2_xuser_f = rd_resp_desc_5_xuser_2_reg[31:0];
   assign rd_resp_desc_5_xuser_3_xuser_f = rd_resp_desc_5_xuser_3_reg[31:0];
   assign rd_resp_desc_5_xuser_4_xuser_f = rd_resp_desc_5_xuser_4_reg[31:0];
   assign rd_resp_desc_5_xuser_5_xuser_f = rd_resp_desc_5_xuser_5_reg[31:0];
   assign rd_resp_desc_5_xuser_6_xuser_f = rd_resp_desc_5_xuser_6_reg[31:0];
   assign rd_resp_desc_5_xuser_7_xuser_f = rd_resp_desc_5_xuser_7_reg[31:0];
   assign rd_resp_desc_5_xuser_8_xuser_f = rd_resp_desc_5_xuser_8_reg[31:0];
   assign rd_resp_desc_5_xuser_9_xuser_f = rd_resp_desc_5_xuser_9_reg[31:0];
   assign rd_resp_desc_5_xuser_10_xuser_f = rd_resp_desc_5_xuser_10_reg[31:0];
   assign rd_resp_desc_5_xuser_11_xuser_f = rd_resp_desc_5_xuser_11_reg[31:0];
   assign rd_resp_desc_5_xuser_12_xuser_f = rd_resp_desc_5_xuser_12_reg[31:0];
   assign rd_resp_desc_5_xuser_13_xuser_f = rd_resp_desc_5_xuser_13_reg[31:0];
   assign rd_resp_desc_5_xuser_14_xuser_f = rd_resp_desc_5_xuser_14_reg[31:0];
   assign rd_resp_desc_5_xuser_15_xuser_f = rd_resp_desc_5_xuser_15_reg[31:0];
   assign wr_req_desc_5_txn_type_wr_strb_f = wr_req_desc_5_txn_type_reg[1];
   assign wr_req_desc_5_size_txn_size_f = wr_req_desc_5_size_reg[31:0];
   assign wr_req_desc_5_data_offset_addr_f = wr_req_desc_5_data_offset_reg[13:0];
   assign wr_req_desc_5_data_host_addr_0_addr_f = wr_req_desc_5_data_host_addr_0_reg[31:0];
   assign wr_req_desc_5_data_host_addr_1_addr_f = wr_req_desc_5_data_host_addr_1_reg[31:0];
   assign wr_req_desc_5_data_host_addr_2_addr_f = wr_req_desc_5_data_host_addr_2_reg[31:0];
   assign wr_req_desc_5_data_host_addr_3_addr_f = wr_req_desc_5_data_host_addr_3_reg[31:0];
   assign wr_req_desc_5_wstrb_host_addr_0_addr_f = wr_req_desc_5_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_5_wstrb_host_addr_1_addr_f = wr_req_desc_5_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_5_wstrb_host_addr_2_addr_f = wr_req_desc_5_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_5_wstrb_host_addr_3_addr_f = wr_req_desc_5_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_5_axsize_axsize_f = wr_req_desc_5_axsize_reg[2:0];
   assign wr_req_desc_5_attr_axsnoop_f = wr_req_desc_5_attr_reg[27:24];
   assign wr_req_desc_5_attr_axdomain_f = wr_req_desc_5_attr_reg[23:22];
   assign wr_req_desc_5_attr_axbar_f = wr_req_desc_5_attr_reg[21:20];
   assign wr_req_desc_5_attr_awunique_f = wr_req_desc_5_attr_reg[19];
   assign wr_req_desc_5_attr_axregion_f = wr_req_desc_5_attr_reg[18:15];
   assign wr_req_desc_5_attr_axqos_f = wr_req_desc_5_attr_reg[14:11];
   assign wr_req_desc_5_attr_axprot_f = wr_req_desc_5_attr_reg[10:8];
   assign wr_req_desc_5_attr_axcache_f = wr_req_desc_5_attr_reg[7:4];
   assign wr_req_desc_5_attr_axlock_f = wr_req_desc_5_attr_reg[2];
   assign wr_req_desc_5_attr_axburst_f = wr_req_desc_5_attr_reg[1:0];
   assign wr_req_desc_5_axaddr_0_addr_f = wr_req_desc_5_axaddr_0_reg[31:0];
   assign wr_req_desc_5_axaddr_1_addr_f = wr_req_desc_5_axaddr_1_reg[31:0];
   assign wr_req_desc_5_axaddr_2_addr_f = wr_req_desc_5_axaddr_2_reg[31:0];
   assign wr_req_desc_5_axaddr_3_addr_f = wr_req_desc_5_axaddr_3_reg[31:0];
   assign wr_req_desc_5_axid_0_axid_f = wr_req_desc_5_axid_0_reg[31:0];
   assign wr_req_desc_5_axid_1_axid_f = wr_req_desc_5_axid_1_reg[31:0];
   assign wr_req_desc_5_axid_2_axid_f = wr_req_desc_5_axid_2_reg[31:0];
   assign wr_req_desc_5_axid_3_axid_f = wr_req_desc_5_axid_3_reg[31:0];
   assign wr_req_desc_5_axuser_0_axuser_f = wr_req_desc_5_axuser_0_reg[31:0];
   assign wr_req_desc_5_axuser_1_axuser_f = wr_req_desc_5_axuser_1_reg[31:0];
   assign wr_req_desc_5_axuser_2_axuser_f = wr_req_desc_5_axuser_2_reg[31:0];
   assign wr_req_desc_5_axuser_3_axuser_f = wr_req_desc_5_axuser_3_reg[31:0];
   assign wr_req_desc_5_axuser_4_axuser_f = wr_req_desc_5_axuser_4_reg[31:0];
   assign wr_req_desc_5_axuser_5_axuser_f = wr_req_desc_5_axuser_5_reg[31:0];
   assign wr_req_desc_5_axuser_6_axuser_f = wr_req_desc_5_axuser_6_reg[31:0];
   assign wr_req_desc_5_axuser_7_axuser_f = wr_req_desc_5_axuser_7_reg[31:0];
   assign wr_req_desc_5_axuser_8_axuser_f = wr_req_desc_5_axuser_8_reg[31:0];
   assign wr_req_desc_5_axuser_9_axuser_f = wr_req_desc_5_axuser_9_reg[31:0];
   assign wr_req_desc_5_axuser_10_axuser_f = wr_req_desc_5_axuser_10_reg[31:0];
   assign wr_req_desc_5_axuser_11_axuser_f = wr_req_desc_5_axuser_11_reg[31:0];
   assign wr_req_desc_5_axuser_12_axuser_f = wr_req_desc_5_axuser_12_reg[31:0];
   assign wr_req_desc_5_axuser_13_axuser_f = wr_req_desc_5_axuser_13_reg[31:0];
   assign wr_req_desc_5_axuser_14_axuser_f = wr_req_desc_5_axuser_14_reg[31:0];
   assign wr_req_desc_5_axuser_15_axuser_f = wr_req_desc_5_axuser_15_reg[31:0];
   assign wr_req_desc_5_wuser_0_wuser_f = wr_req_desc_5_wuser_0_reg[31:0];
   assign wr_req_desc_5_wuser_1_wuser_f = wr_req_desc_5_wuser_1_reg[31:0];
   assign wr_req_desc_5_wuser_2_wuser_f = wr_req_desc_5_wuser_2_reg[31:0];
   assign wr_req_desc_5_wuser_3_wuser_f = wr_req_desc_5_wuser_3_reg[31:0];
   assign wr_req_desc_5_wuser_4_wuser_f = wr_req_desc_5_wuser_4_reg[31:0];
   assign wr_req_desc_5_wuser_5_wuser_f = wr_req_desc_5_wuser_5_reg[31:0];
   assign wr_req_desc_5_wuser_6_wuser_f = wr_req_desc_5_wuser_6_reg[31:0];
   assign wr_req_desc_5_wuser_7_wuser_f = wr_req_desc_5_wuser_7_reg[31:0];
   assign wr_req_desc_5_wuser_8_wuser_f = wr_req_desc_5_wuser_8_reg[31:0];
   assign wr_req_desc_5_wuser_9_wuser_f = wr_req_desc_5_wuser_9_reg[31:0];
   assign wr_req_desc_5_wuser_10_wuser_f = wr_req_desc_5_wuser_10_reg[31:0];
   assign wr_req_desc_5_wuser_11_wuser_f = wr_req_desc_5_wuser_11_reg[31:0];
   assign wr_req_desc_5_wuser_12_wuser_f = wr_req_desc_5_wuser_12_reg[31:0];
   assign wr_req_desc_5_wuser_13_wuser_f = wr_req_desc_5_wuser_13_reg[31:0];
   assign wr_req_desc_5_wuser_14_wuser_f = wr_req_desc_5_wuser_14_reg[31:0];
   assign wr_req_desc_5_wuser_15_wuser_f = wr_req_desc_5_wuser_15_reg[31:0];
   assign wr_resp_desc_5_resp_resp_f = wr_resp_desc_5_resp_reg[4:0];
   assign wr_resp_desc_5_xid_0_xid_f = wr_resp_desc_5_xid_0_reg[31:0];
   assign wr_resp_desc_5_xid_1_xid_f = wr_resp_desc_5_xid_1_reg[31:0];
   assign wr_resp_desc_5_xid_2_xid_f = wr_resp_desc_5_xid_2_reg[31:0];
   assign wr_resp_desc_5_xid_3_xid_f = wr_resp_desc_5_xid_3_reg[31:0];
   assign wr_resp_desc_5_xuser_0_xuser_f = wr_resp_desc_5_xuser_0_reg[31:0];
   assign wr_resp_desc_5_xuser_1_xuser_f = wr_resp_desc_5_xuser_1_reg[31:0];
   assign wr_resp_desc_5_xuser_2_xuser_f = wr_resp_desc_5_xuser_2_reg[31:0];
   assign wr_resp_desc_5_xuser_3_xuser_f = wr_resp_desc_5_xuser_3_reg[31:0];
   assign wr_resp_desc_5_xuser_4_xuser_f = wr_resp_desc_5_xuser_4_reg[31:0];
   assign wr_resp_desc_5_xuser_5_xuser_f = wr_resp_desc_5_xuser_5_reg[31:0];
   assign wr_resp_desc_5_xuser_6_xuser_f = wr_resp_desc_5_xuser_6_reg[31:0];
   assign wr_resp_desc_5_xuser_7_xuser_f = wr_resp_desc_5_xuser_7_reg[31:0];
   assign wr_resp_desc_5_xuser_8_xuser_f = wr_resp_desc_5_xuser_8_reg[31:0];
   assign wr_resp_desc_5_xuser_9_xuser_f = wr_resp_desc_5_xuser_9_reg[31:0];
   assign wr_resp_desc_5_xuser_10_xuser_f = wr_resp_desc_5_xuser_10_reg[31:0];
   assign wr_resp_desc_5_xuser_11_xuser_f = wr_resp_desc_5_xuser_11_reg[31:0];
   assign wr_resp_desc_5_xuser_12_xuser_f = wr_resp_desc_5_xuser_12_reg[31:0];
   assign wr_resp_desc_5_xuser_13_xuser_f = wr_resp_desc_5_xuser_13_reg[31:0];
   assign wr_resp_desc_5_xuser_14_xuser_f = wr_resp_desc_5_xuser_14_reg[31:0];
   assign wr_resp_desc_5_xuser_15_xuser_f = wr_resp_desc_5_xuser_15_reg[31:0];
   assign sn_req_desc_5_attr_acsnoop_f = sn_req_desc_5_attr_reg[27:24];
   assign sn_req_desc_5_attr_acprot_f = sn_req_desc_5_attr_reg[10:8];
   assign sn_req_desc_5_acaddr_0_addr_f = sn_req_desc_5_acaddr_0_reg[31:0];
   assign sn_req_desc_5_acaddr_1_addr_f = sn_req_desc_5_acaddr_1_reg[31:0];
   assign sn_req_desc_5_acaddr_2_addr_f = sn_req_desc_5_acaddr_2_reg[31:0];
   assign sn_req_desc_5_acaddr_3_addr_f = sn_req_desc_5_acaddr_3_reg[31:0];
   assign sn_resp_desc_5_resp_resp_f = sn_resp_desc_5_resp_reg[4:0];
   assign rd_req_desc_6_size_txn_size_f = rd_req_desc_6_size_reg[31:0];
   assign rd_req_desc_6_axsize_axsize_f = rd_req_desc_6_axsize_reg[2:0];
   assign rd_req_desc_6_attr_axsnoop_f = rd_req_desc_6_attr_reg[27:24];
   assign rd_req_desc_6_attr_axdomain_f = rd_req_desc_6_attr_reg[23:22];
   assign rd_req_desc_6_attr_axbar_f = rd_req_desc_6_attr_reg[21:20];
   assign rd_req_desc_6_attr_axregion_f = rd_req_desc_6_attr_reg[18:15];
   assign rd_req_desc_6_attr_axqos_f = rd_req_desc_6_attr_reg[14:11];
   assign rd_req_desc_6_attr_axprot_f = rd_req_desc_6_attr_reg[10:8];
   assign rd_req_desc_6_attr_axcache_f = rd_req_desc_6_attr_reg[7:4];
   assign rd_req_desc_6_attr_axlock_f = rd_req_desc_6_attr_reg[2];
   assign rd_req_desc_6_attr_axburst_f = rd_req_desc_6_attr_reg[1:0];
   assign rd_req_desc_6_axaddr_0_addr_f = rd_req_desc_6_axaddr_0_reg[31:0];
   assign rd_req_desc_6_axaddr_1_addr_f = rd_req_desc_6_axaddr_1_reg[31:0];
   assign rd_req_desc_6_axaddr_2_addr_f = rd_req_desc_6_axaddr_2_reg[31:0];
   assign rd_req_desc_6_axaddr_3_addr_f = rd_req_desc_6_axaddr_3_reg[31:0];
   assign rd_req_desc_6_axid_0_axid_f = rd_req_desc_6_axid_0_reg[31:0];
   assign rd_req_desc_6_axid_1_axid_f = rd_req_desc_6_axid_1_reg[31:0];
   assign rd_req_desc_6_axid_2_axid_f = rd_req_desc_6_axid_2_reg[31:0];
   assign rd_req_desc_6_axid_3_axid_f = rd_req_desc_6_axid_3_reg[31:0];
   assign rd_req_desc_6_axuser_0_axuser_f = rd_req_desc_6_axuser_0_reg[31:0];
   assign rd_req_desc_6_axuser_1_axuser_f = rd_req_desc_6_axuser_1_reg[31:0];
   assign rd_req_desc_6_axuser_2_axuser_f = rd_req_desc_6_axuser_2_reg[31:0];
   assign rd_req_desc_6_axuser_3_axuser_f = rd_req_desc_6_axuser_3_reg[31:0];
   assign rd_req_desc_6_axuser_4_axuser_f = rd_req_desc_6_axuser_4_reg[31:0];
   assign rd_req_desc_6_axuser_5_axuser_f = rd_req_desc_6_axuser_5_reg[31:0];
   assign rd_req_desc_6_axuser_6_axuser_f = rd_req_desc_6_axuser_6_reg[31:0];
   assign rd_req_desc_6_axuser_7_axuser_f = rd_req_desc_6_axuser_7_reg[31:0];
   assign rd_req_desc_6_axuser_8_axuser_f = rd_req_desc_6_axuser_8_reg[31:0];
   assign rd_req_desc_6_axuser_9_axuser_f = rd_req_desc_6_axuser_9_reg[31:0];
   assign rd_req_desc_6_axuser_10_axuser_f = rd_req_desc_6_axuser_10_reg[31:0];
   assign rd_req_desc_6_axuser_11_axuser_f = rd_req_desc_6_axuser_11_reg[31:0];
   assign rd_req_desc_6_axuser_12_axuser_f = rd_req_desc_6_axuser_12_reg[31:0];
   assign rd_req_desc_6_axuser_13_axuser_f = rd_req_desc_6_axuser_13_reg[31:0];
   assign rd_req_desc_6_axuser_14_axuser_f = rd_req_desc_6_axuser_14_reg[31:0];
   assign rd_req_desc_6_axuser_15_axuser_f = rd_req_desc_6_axuser_15_reg[31:0];
   assign rd_resp_desc_6_data_offset_addr_f = rd_resp_desc_6_data_offset_reg[13:0];
   assign rd_resp_desc_6_data_size_size_f = rd_resp_desc_6_data_size_reg[31:0];
   assign rd_resp_desc_6_data_host_addr_0_addr_f = rd_resp_desc_6_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_6_data_host_addr_1_addr_f = rd_resp_desc_6_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_6_data_host_addr_2_addr_f = rd_resp_desc_6_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_6_data_host_addr_3_addr_f = rd_resp_desc_6_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_6_resp_resp_f = rd_resp_desc_6_resp_reg[4:0];
   assign rd_resp_desc_6_xid_0_xid_f = rd_resp_desc_6_xid_0_reg[31:0];
   assign rd_resp_desc_6_xid_1_xid_f = rd_resp_desc_6_xid_1_reg[31:0];
   assign rd_resp_desc_6_xid_2_xid_f = rd_resp_desc_6_xid_2_reg[31:0];
   assign rd_resp_desc_6_xid_3_xid_f = rd_resp_desc_6_xid_3_reg[31:0];
   assign rd_resp_desc_6_xuser_0_xuser_f = rd_resp_desc_6_xuser_0_reg[31:0];
   assign rd_resp_desc_6_xuser_1_xuser_f = rd_resp_desc_6_xuser_1_reg[31:0];
   assign rd_resp_desc_6_xuser_2_xuser_f = rd_resp_desc_6_xuser_2_reg[31:0];
   assign rd_resp_desc_6_xuser_3_xuser_f = rd_resp_desc_6_xuser_3_reg[31:0];
   assign rd_resp_desc_6_xuser_4_xuser_f = rd_resp_desc_6_xuser_4_reg[31:0];
   assign rd_resp_desc_6_xuser_5_xuser_f = rd_resp_desc_6_xuser_5_reg[31:0];
   assign rd_resp_desc_6_xuser_6_xuser_f = rd_resp_desc_6_xuser_6_reg[31:0];
   assign rd_resp_desc_6_xuser_7_xuser_f = rd_resp_desc_6_xuser_7_reg[31:0];
   assign rd_resp_desc_6_xuser_8_xuser_f = rd_resp_desc_6_xuser_8_reg[31:0];
   assign rd_resp_desc_6_xuser_9_xuser_f = rd_resp_desc_6_xuser_9_reg[31:0];
   assign rd_resp_desc_6_xuser_10_xuser_f = rd_resp_desc_6_xuser_10_reg[31:0];
   assign rd_resp_desc_6_xuser_11_xuser_f = rd_resp_desc_6_xuser_11_reg[31:0];
   assign rd_resp_desc_6_xuser_12_xuser_f = rd_resp_desc_6_xuser_12_reg[31:0];
   assign rd_resp_desc_6_xuser_13_xuser_f = rd_resp_desc_6_xuser_13_reg[31:0];
   assign rd_resp_desc_6_xuser_14_xuser_f = rd_resp_desc_6_xuser_14_reg[31:0];
   assign rd_resp_desc_6_xuser_15_xuser_f = rd_resp_desc_6_xuser_15_reg[31:0];
   assign wr_req_desc_6_txn_type_wr_strb_f = wr_req_desc_6_txn_type_reg[1];
   assign wr_req_desc_6_size_txn_size_f = wr_req_desc_6_size_reg[31:0];
   assign wr_req_desc_6_data_offset_addr_f = wr_req_desc_6_data_offset_reg[13:0];
   assign wr_req_desc_6_data_host_addr_0_addr_f = wr_req_desc_6_data_host_addr_0_reg[31:0];
   assign wr_req_desc_6_data_host_addr_1_addr_f = wr_req_desc_6_data_host_addr_1_reg[31:0];
   assign wr_req_desc_6_data_host_addr_2_addr_f = wr_req_desc_6_data_host_addr_2_reg[31:0];
   assign wr_req_desc_6_data_host_addr_3_addr_f = wr_req_desc_6_data_host_addr_3_reg[31:0];
   assign wr_req_desc_6_wstrb_host_addr_0_addr_f = wr_req_desc_6_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_6_wstrb_host_addr_1_addr_f = wr_req_desc_6_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_6_wstrb_host_addr_2_addr_f = wr_req_desc_6_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_6_wstrb_host_addr_3_addr_f = wr_req_desc_6_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_6_axsize_axsize_f = wr_req_desc_6_axsize_reg[2:0];
   assign wr_req_desc_6_attr_axsnoop_f = wr_req_desc_6_attr_reg[27:24];
   assign wr_req_desc_6_attr_axdomain_f = wr_req_desc_6_attr_reg[23:22];
   assign wr_req_desc_6_attr_axbar_f = wr_req_desc_6_attr_reg[21:20];
   assign wr_req_desc_6_attr_awunique_f = wr_req_desc_6_attr_reg[19];
   assign wr_req_desc_6_attr_axregion_f = wr_req_desc_6_attr_reg[18:15];
   assign wr_req_desc_6_attr_axqos_f = wr_req_desc_6_attr_reg[14:11];
   assign wr_req_desc_6_attr_axprot_f = wr_req_desc_6_attr_reg[10:8];
   assign wr_req_desc_6_attr_axcache_f = wr_req_desc_6_attr_reg[7:4];
   assign wr_req_desc_6_attr_axlock_f = wr_req_desc_6_attr_reg[2];
   assign wr_req_desc_6_attr_axburst_f = wr_req_desc_6_attr_reg[1:0];
   assign wr_req_desc_6_axaddr_0_addr_f = wr_req_desc_6_axaddr_0_reg[31:0];
   assign wr_req_desc_6_axaddr_1_addr_f = wr_req_desc_6_axaddr_1_reg[31:0];
   assign wr_req_desc_6_axaddr_2_addr_f = wr_req_desc_6_axaddr_2_reg[31:0];
   assign wr_req_desc_6_axaddr_3_addr_f = wr_req_desc_6_axaddr_3_reg[31:0];
   assign wr_req_desc_6_axid_0_axid_f = wr_req_desc_6_axid_0_reg[31:0];
   assign wr_req_desc_6_axid_1_axid_f = wr_req_desc_6_axid_1_reg[31:0];
   assign wr_req_desc_6_axid_2_axid_f = wr_req_desc_6_axid_2_reg[31:0];
   assign wr_req_desc_6_axid_3_axid_f = wr_req_desc_6_axid_3_reg[31:0];
   assign wr_req_desc_6_axuser_0_axuser_f = wr_req_desc_6_axuser_0_reg[31:0];
   assign wr_req_desc_6_axuser_1_axuser_f = wr_req_desc_6_axuser_1_reg[31:0];
   assign wr_req_desc_6_axuser_2_axuser_f = wr_req_desc_6_axuser_2_reg[31:0];
   assign wr_req_desc_6_axuser_3_axuser_f = wr_req_desc_6_axuser_3_reg[31:0];
   assign wr_req_desc_6_axuser_4_axuser_f = wr_req_desc_6_axuser_4_reg[31:0];
   assign wr_req_desc_6_axuser_5_axuser_f = wr_req_desc_6_axuser_5_reg[31:0];
   assign wr_req_desc_6_axuser_6_axuser_f = wr_req_desc_6_axuser_6_reg[31:0];
   assign wr_req_desc_6_axuser_7_axuser_f = wr_req_desc_6_axuser_7_reg[31:0];
   assign wr_req_desc_6_axuser_8_axuser_f = wr_req_desc_6_axuser_8_reg[31:0];
   assign wr_req_desc_6_axuser_9_axuser_f = wr_req_desc_6_axuser_9_reg[31:0];
   assign wr_req_desc_6_axuser_10_axuser_f = wr_req_desc_6_axuser_10_reg[31:0];
   assign wr_req_desc_6_axuser_11_axuser_f = wr_req_desc_6_axuser_11_reg[31:0];
   assign wr_req_desc_6_axuser_12_axuser_f = wr_req_desc_6_axuser_12_reg[31:0];
   assign wr_req_desc_6_axuser_13_axuser_f = wr_req_desc_6_axuser_13_reg[31:0];
   assign wr_req_desc_6_axuser_14_axuser_f = wr_req_desc_6_axuser_14_reg[31:0];
   assign wr_req_desc_6_axuser_15_axuser_f = wr_req_desc_6_axuser_15_reg[31:0];
   assign wr_req_desc_6_wuser_0_wuser_f = wr_req_desc_6_wuser_0_reg[31:0];
   assign wr_req_desc_6_wuser_1_wuser_f = wr_req_desc_6_wuser_1_reg[31:0];
   assign wr_req_desc_6_wuser_2_wuser_f = wr_req_desc_6_wuser_2_reg[31:0];
   assign wr_req_desc_6_wuser_3_wuser_f = wr_req_desc_6_wuser_3_reg[31:0];
   assign wr_req_desc_6_wuser_4_wuser_f = wr_req_desc_6_wuser_4_reg[31:0];
   assign wr_req_desc_6_wuser_5_wuser_f = wr_req_desc_6_wuser_5_reg[31:0];
   assign wr_req_desc_6_wuser_6_wuser_f = wr_req_desc_6_wuser_6_reg[31:0];
   assign wr_req_desc_6_wuser_7_wuser_f = wr_req_desc_6_wuser_7_reg[31:0];
   assign wr_req_desc_6_wuser_8_wuser_f = wr_req_desc_6_wuser_8_reg[31:0];
   assign wr_req_desc_6_wuser_9_wuser_f = wr_req_desc_6_wuser_9_reg[31:0];
   assign wr_req_desc_6_wuser_10_wuser_f = wr_req_desc_6_wuser_10_reg[31:0];
   assign wr_req_desc_6_wuser_11_wuser_f = wr_req_desc_6_wuser_11_reg[31:0];
   assign wr_req_desc_6_wuser_12_wuser_f = wr_req_desc_6_wuser_12_reg[31:0];
   assign wr_req_desc_6_wuser_13_wuser_f = wr_req_desc_6_wuser_13_reg[31:0];
   assign wr_req_desc_6_wuser_14_wuser_f = wr_req_desc_6_wuser_14_reg[31:0];
   assign wr_req_desc_6_wuser_15_wuser_f = wr_req_desc_6_wuser_15_reg[31:0];
   assign wr_resp_desc_6_resp_resp_f = wr_resp_desc_6_resp_reg[4:0];
   assign wr_resp_desc_6_xid_0_xid_f = wr_resp_desc_6_xid_0_reg[31:0];
   assign wr_resp_desc_6_xid_1_xid_f = wr_resp_desc_6_xid_1_reg[31:0];
   assign wr_resp_desc_6_xid_2_xid_f = wr_resp_desc_6_xid_2_reg[31:0];
   assign wr_resp_desc_6_xid_3_xid_f = wr_resp_desc_6_xid_3_reg[31:0];
   assign wr_resp_desc_6_xuser_0_xuser_f = wr_resp_desc_6_xuser_0_reg[31:0];
   assign wr_resp_desc_6_xuser_1_xuser_f = wr_resp_desc_6_xuser_1_reg[31:0];
   assign wr_resp_desc_6_xuser_2_xuser_f = wr_resp_desc_6_xuser_2_reg[31:0];
   assign wr_resp_desc_6_xuser_3_xuser_f = wr_resp_desc_6_xuser_3_reg[31:0];
   assign wr_resp_desc_6_xuser_4_xuser_f = wr_resp_desc_6_xuser_4_reg[31:0];
   assign wr_resp_desc_6_xuser_5_xuser_f = wr_resp_desc_6_xuser_5_reg[31:0];
   assign wr_resp_desc_6_xuser_6_xuser_f = wr_resp_desc_6_xuser_6_reg[31:0];
   assign wr_resp_desc_6_xuser_7_xuser_f = wr_resp_desc_6_xuser_7_reg[31:0];
   assign wr_resp_desc_6_xuser_8_xuser_f = wr_resp_desc_6_xuser_8_reg[31:0];
   assign wr_resp_desc_6_xuser_9_xuser_f = wr_resp_desc_6_xuser_9_reg[31:0];
   assign wr_resp_desc_6_xuser_10_xuser_f = wr_resp_desc_6_xuser_10_reg[31:0];
   assign wr_resp_desc_6_xuser_11_xuser_f = wr_resp_desc_6_xuser_11_reg[31:0];
   assign wr_resp_desc_6_xuser_12_xuser_f = wr_resp_desc_6_xuser_12_reg[31:0];
   assign wr_resp_desc_6_xuser_13_xuser_f = wr_resp_desc_6_xuser_13_reg[31:0];
   assign wr_resp_desc_6_xuser_14_xuser_f = wr_resp_desc_6_xuser_14_reg[31:0];
   assign wr_resp_desc_6_xuser_15_xuser_f = wr_resp_desc_6_xuser_15_reg[31:0];
   assign sn_req_desc_6_attr_acsnoop_f = sn_req_desc_6_attr_reg[27:24];
   assign sn_req_desc_6_attr_acprot_f = sn_req_desc_6_attr_reg[10:8];
   assign sn_req_desc_6_acaddr_0_addr_f = sn_req_desc_6_acaddr_0_reg[31:0];
   assign sn_req_desc_6_acaddr_1_addr_f = sn_req_desc_6_acaddr_1_reg[31:0];
   assign sn_req_desc_6_acaddr_2_addr_f = sn_req_desc_6_acaddr_2_reg[31:0];
   assign sn_req_desc_6_acaddr_3_addr_f = sn_req_desc_6_acaddr_3_reg[31:0];
   assign sn_resp_desc_6_resp_resp_f = sn_resp_desc_6_resp_reg[4:0];
   assign rd_req_desc_7_size_txn_size_f = rd_req_desc_7_size_reg[31:0];
   assign rd_req_desc_7_axsize_axsize_f = rd_req_desc_7_axsize_reg[2:0];
   assign rd_req_desc_7_attr_axsnoop_f = rd_req_desc_7_attr_reg[27:24];
   assign rd_req_desc_7_attr_axdomain_f = rd_req_desc_7_attr_reg[23:22];
   assign rd_req_desc_7_attr_axbar_f = rd_req_desc_7_attr_reg[21:20];
   assign rd_req_desc_7_attr_axregion_f = rd_req_desc_7_attr_reg[18:15];
   assign rd_req_desc_7_attr_axqos_f = rd_req_desc_7_attr_reg[14:11];
   assign rd_req_desc_7_attr_axprot_f = rd_req_desc_7_attr_reg[10:8];
   assign rd_req_desc_7_attr_axcache_f = rd_req_desc_7_attr_reg[7:4];
   assign rd_req_desc_7_attr_axlock_f = rd_req_desc_7_attr_reg[2];
   assign rd_req_desc_7_attr_axburst_f = rd_req_desc_7_attr_reg[1:0];
   assign rd_req_desc_7_axaddr_0_addr_f = rd_req_desc_7_axaddr_0_reg[31:0];
   assign rd_req_desc_7_axaddr_1_addr_f = rd_req_desc_7_axaddr_1_reg[31:0];
   assign rd_req_desc_7_axaddr_2_addr_f = rd_req_desc_7_axaddr_2_reg[31:0];
   assign rd_req_desc_7_axaddr_3_addr_f = rd_req_desc_7_axaddr_3_reg[31:0];
   assign rd_req_desc_7_axid_0_axid_f = rd_req_desc_7_axid_0_reg[31:0];
   assign rd_req_desc_7_axid_1_axid_f = rd_req_desc_7_axid_1_reg[31:0];
   assign rd_req_desc_7_axid_2_axid_f = rd_req_desc_7_axid_2_reg[31:0];
   assign rd_req_desc_7_axid_3_axid_f = rd_req_desc_7_axid_3_reg[31:0];
   assign rd_req_desc_7_axuser_0_axuser_f = rd_req_desc_7_axuser_0_reg[31:0];
   assign rd_req_desc_7_axuser_1_axuser_f = rd_req_desc_7_axuser_1_reg[31:0];
   assign rd_req_desc_7_axuser_2_axuser_f = rd_req_desc_7_axuser_2_reg[31:0];
   assign rd_req_desc_7_axuser_3_axuser_f = rd_req_desc_7_axuser_3_reg[31:0];
   assign rd_req_desc_7_axuser_4_axuser_f = rd_req_desc_7_axuser_4_reg[31:0];
   assign rd_req_desc_7_axuser_5_axuser_f = rd_req_desc_7_axuser_5_reg[31:0];
   assign rd_req_desc_7_axuser_6_axuser_f = rd_req_desc_7_axuser_6_reg[31:0];
   assign rd_req_desc_7_axuser_7_axuser_f = rd_req_desc_7_axuser_7_reg[31:0];
   assign rd_req_desc_7_axuser_8_axuser_f = rd_req_desc_7_axuser_8_reg[31:0];
   assign rd_req_desc_7_axuser_9_axuser_f = rd_req_desc_7_axuser_9_reg[31:0];
   assign rd_req_desc_7_axuser_10_axuser_f = rd_req_desc_7_axuser_10_reg[31:0];
   assign rd_req_desc_7_axuser_11_axuser_f = rd_req_desc_7_axuser_11_reg[31:0];
   assign rd_req_desc_7_axuser_12_axuser_f = rd_req_desc_7_axuser_12_reg[31:0];
   assign rd_req_desc_7_axuser_13_axuser_f = rd_req_desc_7_axuser_13_reg[31:0];
   assign rd_req_desc_7_axuser_14_axuser_f = rd_req_desc_7_axuser_14_reg[31:0];
   assign rd_req_desc_7_axuser_15_axuser_f = rd_req_desc_7_axuser_15_reg[31:0];
   assign rd_resp_desc_7_data_offset_addr_f = rd_resp_desc_7_data_offset_reg[13:0];
   assign rd_resp_desc_7_data_size_size_f = rd_resp_desc_7_data_size_reg[31:0];
   assign rd_resp_desc_7_data_host_addr_0_addr_f = rd_resp_desc_7_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_7_data_host_addr_1_addr_f = rd_resp_desc_7_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_7_data_host_addr_2_addr_f = rd_resp_desc_7_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_7_data_host_addr_3_addr_f = rd_resp_desc_7_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_7_resp_resp_f = rd_resp_desc_7_resp_reg[4:0];
   assign rd_resp_desc_7_xid_0_xid_f = rd_resp_desc_7_xid_0_reg[31:0];
   assign rd_resp_desc_7_xid_1_xid_f = rd_resp_desc_7_xid_1_reg[31:0];
   assign rd_resp_desc_7_xid_2_xid_f = rd_resp_desc_7_xid_2_reg[31:0];
   assign rd_resp_desc_7_xid_3_xid_f = rd_resp_desc_7_xid_3_reg[31:0];
   assign rd_resp_desc_7_xuser_0_xuser_f = rd_resp_desc_7_xuser_0_reg[31:0];
   assign rd_resp_desc_7_xuser_1_xuser_f = rd_resp_desc_7_xuser_1_reg[31:0];
   assign rd_resp_desc_7_xuser_2_xuser_f = rd_resp_desc_7_xuser_2_reg[31:0];
   assign rd_resp_desc_7_xuser_3_xuser_f = rd_resp_desc_7_xuser_3_reg[31:0];
   assign rd_resp_desc_7_xuser_4_xuser_f = rd_resp_desc_7_xuser_4_reg[31:0];
   assign rd_resp_desc_7_xuser_5_xuser_f = rd_resp_desc_7_xuser_5_reg[31:0];
   assign rd_resp_desc_7_xuser_6_xuser_f = rd_resp_desc_7_xuser_6_reg[31:0];
   assign rd_resp_desc_7_xuser_7_xuser_f = rd_resp_desc_7_xuser_7_reg[31:0];
   assign rd_resp_desc_7_xuser_8_xuser_f = rd_resp_desc_7_xuser_8_reg[31:0];
   assign rd_resp_desc_7_xuser_9_xuser_f = rd_resp_desc_7_xuser_9_reg[31:0];
   assign rd_resp_desc_7_xuser_10_xuser_f = rd_resp_desc_7_xuser_10_reg[31:0];
   assign rd_resp_desc_7_xuser_11_xuser_f = rd_resp_desc_7_xuser_11_reg[31:0];
   assign rd_resp_desc_7_xuser_12_xuser_f = rd_resp_desc_7_xuser_12_reg[31:0];
   assign rd_resp_desc_7_xuser_13_xuser_f = rd_resp_desc_7_xuser_13_reg[31:0];
   assign rd_resp_desc_7_xuser_14_xuser_f = rd_resp_desc_7_xuser_14_reg[31:0];
   assign rd_resp_desc_7_xuser_15_xuser_f = rd_resp_desc_7_xuser_15_reg[31:0];
   assign wr_req_desc_7_txn_type_wr_strb_f = wr_req_desc_7_txn_type_reg[1];
   assign wr_req_desc_7_size_txn_size_f = wr_req_desc_7_size_reg[31:0];
   assign wr_req_desc_7_data_offset_addr_f = wr_req_desc_7_data_offset_reg[13:0];
   assign wr_req_desc_7_data_host_addr_0_addr_f = wr_req_desc_7_data_host_addr_0_reg[31:0];
   assign wr_req_desc_7_data_host_addr_1_addr_f = wr_req_desc_7_data_host_addr_1_reg[31:0];
   assign wr_req_desc_7_data_host_addr_2_addr_f = wr_req_desc_7_data_host_addr_2_reg[31:0];
   assign wr_req_desc_7_data_host_addr_3_addr_f = wr_req_desc_7_data_host_addr_3_reg[31:0];
   assign wr_req_desc_7_wstrb_host_addr_0_addr_f = wr_req_desc_7_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_7_wstrb_host_addr_1_addr_f = wr_req_desc_7_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_7_wstrb_host_addr_2_addr_f = wr_req_desc_7_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_7_wstrb_host_addr_3_addr_f = wr_req_desc_7_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_7_axsize_axsize_f = wr_req_desc_7_axsize_reg[2:0];
   assign wr_req_desc_7_attr_axsnoop_f = wr_req_desc_7_attr_reg[27:24];
   assign wr_req_desc_7_attr_axdomain_f = wr_req_desc_7_attr_reg[23:22];
   assign wr_req_desc_7_attr_axbar_f = wr_req_desc_7_attr_reg[21:20];
   assign wr_req_desc_7_attr_awunique_f = wr_req_desc_7_attr_reg[19];
   assign wr_req_desc_7_attr_axregion_f = wr_req_desc_7_attr_reg[18:15];
   assign wr_req_desc_7_attr_axqos_f = wr_req_desc_7_attr_reg[14:11];
   assign wr_req_desc_7_attr_axprot_f = wr_req_desc_7_attr_reg[10:8];
   assign wr_req_desc_7_attr_axcache_f = wr_req_desc_7_attr_reg[7:4];
   assign wr_req_desc_7_attr_axlock_f = wr_req_desc_7_attr_reg[2];
   assign wr_req_desc_7_attr_axburst_f = wr_req_desc_7_attr_reg[1:0];
   assign wr_req_desc_7_axaddr_0_addr_f = wr_req_desc_7_axaddr_0_reg[31:0];
   assign wr_req_desc_7_axaddr_1_addr_f = wr_req_desc_7_axaddr_1_reg[31:0];
   assign wr_req_desc_7_axaddr_2_addr_f = wr_req_desc_7_axaddr_2_reg[31:0];
   assign wr_req_desc_7_axaddr_3_addr_f = wr_req_desc_7_axaddr_3_reg[31:0];
   assign wr_req_desc_7_axid_0_axid_f = wr_req_desc_7_axid_0_reg[31:0];
   assign wr_req_desc_7_axid_1_axid_f = wr_req_desc_7_axid_1_reg[31:0];
   assign wr_req_desc_7_axid_2_axid_f = wr_req_desc_7_axid_2_reg[31:0];
   assign wr_req_desc_7_axid_3_axid_f = wr_req_desc_7_axid_3_reg[31:0];
   assign wr_req_desc_7_axuser_0_axuser_f = wr_req_desc_7_axuser_0_reg[31:0];
   assign wr_req_desc_7_axuser_1_axuser_f = wr_req_desc_7_axuser_1_reg[31:0];
   assign wr_req_desc_7_axuser_2_axuser_f = wr_req_desc_7_axuser_2_reg[31:0];
   assign wr_req_desc_7_axuser_3_axuser_f = wr_req_desc_7_axuser_3_reg[31:0];
   assign wr_req_desc_7_axuser_4_axuser_f = wr_req_desc_7_axuser_4_reg[31:0];
   assign wr_req_desc_7_axuser_5_axuser_f = wr_req_desc_7_axuser_5_reg[31:0];
   assign wr_req_desc_7_axuser_6_axuser_f = wr_req_desc_7_axuser_6_reg[31:0];
   assign wr_req_desc_7_axuser_7_axuser_f = wr_req_desc_7_axuser_7_reg[31:0];
   assign wr_req_desc_7_axuser_8_axuser_f = wr_req_desc_7_axuser_8_reg[31:0];
   assign wr_req_desc_7_axuser_9_axuser_f = wr_req_desc_7_axuser_9_reg[31:0];
   assign wr_req_desc_7_axuser_10_axuser_f = wr_req_desc_7_axuser_10_reg[31:0];
   assign wr_req_desc_7_axuser_11_axuser_f = wr_req_desc_7_axuser_11_reg[31:0];
   assign wr_req_desc_7_axuser_12_axuser_f = wr_req_desc_7_axuser_12_reg[31:0];
   assign wr_req_desc_7_axuser_13_axuser_f = wr_req_desc_7_axuser_13_reg[31:0];
   assign wr_req_desc_7_axuser_14_axuser_f = wr_req_desc_7_axuser_14_reg[31:0];
   assign wr_req_desc_7_axuser_15_axuser_f = wr_req_desc_7_axuser_15_reg[31:0];
   assign wr_req_desc_7_wuser_0_wuser_f = wr_req_desc_7_wuser_0_reg[31:0];
   assign wr_req_desc_7_wuser_1_wuser_f = wr_req_desc_7_wuser_1_reg[31:0];
   assign wr_req_desc_7_wuser_2_wuser_f = wr_req_desc_7_wuser_2_reg[31:0];
   assign wr_req_desc_7_wuser_3_wuser_f = wr_req_desc_7_wuser_3_reg[31:0];
   assign wr_req_desc_7_wuser_4_wuser_f = wr_req_desc_7_wuser_4_reg[31:0];
   assign wr_req_desc_7_wuser_5_wuser_f = wr_req_desc_7_wuser_5_reg[31:0];
   assign wr_req_desc_7_wuser_6_wuser_f = wr_req_desc_7_wuser_6_reg[31:0];
   assign wr_req_desc_7_wuser_7_wuser_f = wr_req_desc_7_wuser_7_reg[31:0];
   assign wr_req_desc_7_wuser_8_wuser_f = wr_req_desc_7_wuser_8_reg[31:0];
   assign wr_req_desc_7_wuser_9_wuser_f = wr_req_desc_7_wuser_9_reg[31:0];
   assign wr_req_desc_7_wuser_10_wuser_f = wr_req_desc_7_wuser_10_reg[31:0];
   assign wr_req_desc_7_wuser_11_wuser_f = wr_req_desc_7_wuser_11_reg[31:0];
   assign wr_req_desc_7_wuser_12_wuser_f = wr_req_desc_7_wuser_12_reg[31:0];
   assign wr_req_desc_7_wuser_13_wuser_f = wr_req_desc_7_wuser_13_reg[31:0];
   assign wr_req_desc_7_wuser_14_wuser_f = wr_req_desc_7_wuser_14_reg[31:0];
   assign wr_req_desc_7_wuser_15_wuser_f = wr_req_desc_7_wuser_15_reg[31:0];
   assign wr_resp_desc_7_resp_resp_f = wr_resp_desc_7_resp_reg[4:0];
   assign wr_resp_desc_7_xid_0_xid_f = wr_resp_desc_7_xid_0_reg[31:0];
   assign wr_resp_desc_7_xid_1_xid_f = wr_resp_desc_7_xid_1_reg[31:0];
   assign wr_resp_desc_7_xid_2_xid_f = wr_resp_desc_7_xid_2_reg[31:0];
   assign wr_resp_desc_7_xid_3_xid_f = wr_resp_desc_7_xid_3_reg[31:0];
   assign wr_resp_desc_7_xuser_0_xuser_f = wr_resp_desc_7_xuser_0_reg[31:0];
   assign wr_resp_desc_7_xuser_1_xuser_f = wr_resp_desc_7_xuser_1_reg[31:0];
   assign wr_resp_desc_7_xuser_2_xuser_f = wr_resp_desc_7_xuser_2_reg[31:0];
   assign wr_resp_desc_7_xuser_3_xuser_f = wr_resp_desc_7_xuser_3_reg[31:0];
   assign wr_resp_desc_7_xuser_4_xuser_f = wr_resp_desc_7_xuser_4_reg[31:0];
   assign wr_resp_desc_7_xuser_5_xuser_f = wr_resp_desc_7_xuser_5_reg[31:0];
   assign wr_resp_desc_7_xuser_6_xuser_f = wr_resp_desc_7_xuser_6_reg[31:0];
   assign wr_resp_desc_7_xuser_7_xuser_f = wr_resp_desc_7_xuser_7_reg[31:0];
   assign wr_resp_desc_7_xuser_8_xuser_f = wr_resp_desc_7_xuser_8_reg[31:0];
   assign wr_resp_desc_7_xuser_9_xuser_f = wr_resp_desc_7_xuser_9_reg[31:0];
   assign wr_resp_desc_7_xuser_10_xuser_f = wr_resp_desc_7_xuser_10_reg[31:0];
   assign wr_resp_desc_7_xuser_11_xuser_f = wr_resp_desc_7_xuser_11_reg[31:0];
   assign wr_resp_desc_7_xuser_12_xuser_f = wr_resp_desc_7_xuser_12_reg[31:0];
   assign wr_resp_desc_7_xuser_13_xuser_f = wr_resp_desc_7_xuser_13_reg[31:0];
   assign wr_resp_desc_7_xuser_14_xuser_f = wr_resp_desc_7_xuser_14_reg[31:0];
   assign wr_resp_desc_7_xuser_15_xuser_f = wr_resp_desc_7_xuser_15_reg[31:0];
   assign sn_req_desc_7_attr_acsnoop_f = sn_req_desc_7_attr_reg[27:24];
   assign sn_req_desc_7_attr_acprot_f = sn_req_desc_7_attr_reg[10:8];
   assign sn_req_desc_7_acaddr_0_addr_f = sn_req_desc_7_acaddr_0_reg[31:0];
   assign sn_req_desc_7_acaddr_1_addr_f = sn_req_desc_7_acaddr_1_reg[31:0];
   assign sn_req_desc_7_acaddr_2_addr_f = sn_req_desc_7_acaddr_2_reg[31:0];
   assign sn_req_desc_7_acaddr_3_addr_f = sn_req_desc_7_acaddr_3_reg[31:0];
   assign sn_resp_desc_7_resp_resp_f = sn_resp_desc_7_resp_reg[4:0];
   assign rd_req_desc_8_size_txn_size_f = rd_req_desc_8_size_reg[31:0];
   assign rd_req_desc_8_axsize_axsize_f = rd_req_desc_8_axsize_reg[2:0];
   assign rd_req_desc_8_attr_axsnoop_f = rd_req_desc_8_attr_reg[27:24];
   assign rd_req_desc_8_attr_axdomain_f = rd_req_desc_8_attr_reg[23:22];
   assign rd_req_desc_8_attr_axbar_f = rd_req_desc_8_attr_reg[21:20];
   assign rd_req_desc_8_attr_axregion_f = rd_req_desc_8_attr_reg[18:15];
   assign rd_req_desc_8_attr_axqos_f = rd_req_desc_8_attr_reg[14:11];
   assign rd_req_desc_8_attr_axprot_f = rd_req_desc_8_attr_reg[10:8];
   assign rd_req_desc_8_attr_axcache_f = rd_req_desc_8_attr_reg[7:4];
   assign rd_req_desc_8_attr_axlock_f = rd_req_desc_8_attr_reg[2];
   assign rd_req_desc_8_attr_axburst_f = rd_req_desc_8_attr_reg[1:0];
   assign rd_req_desc_8_axaddr_0_addr_f = rd_req_desc_8_axaddr_0_reg[31:0];
   assign rd_req_desc_8_axaddr_1_addr_f = rd_req_desc_8_axaddr_1_reg[31:0];
   assign rd_req_desc_8_axaddr_2_addr_f = rd_req_desc_8_axaddr_2_reg[31:0];
   assign rd_req_desc_8_axaddr_3_addr_f = rd_req_desc_8_axaddr_3_reg[31:0];
   assign rd_req_desc_8_axid_0_axid_f = rd_req_desc_8_axid_0_reg[31:0];
   assign rd_req_desc_8_axid_1_axid_f = rd_req_desc_8_axid_1_reg[31:0];
   assign rd_req_desc_8_axid_2_axid_f = rd_req_desc_8_axid_2_reg[31:0];
   assign rd_req_desc_8_axid_3_axid_f = rd_req_desc_8_axid_3_reg[31:0];
   assign rd_req_desc_8_axuser_0_axuser_f = rd_req_desc_8_axuser_0_reg[31:0];
   assign rd_req_desc_8_axuser_1_axuser_f = rd_req_desc_8_axuser_1_reg[31:0];
   assign rd_req_desc_8_axuser_2_axuser_f = rd_req_desc_8_axuser_2_reg[31:0];
   assign rd_req_desc_8_axuser_3_axuser_f = rd_req_desc_8_axuser_3_reg[31:0];
   assign rd_req_desc_8_axuser_4_axuser_f = rd_req_desc_8_axuser_4_reg[31:0];
   assign rd_req_desc_8_axuser_5_axuser_f = rd_req_desc_8_axuser_5_reg[31:0];
   assign rd_req_desc_8_axuser_6_axuser_f = rd_req_desc_8_axuser_6_reg[31:0];
   assign rd_req_desc_8_axuser_7_axuser_f = rd_req_desc_8_axuser_7_reg[31:0];
   assign rd_req_desc_8_axuser_8_axuser_f = rd_req_desc_8_axuser_8_reg[31:0];
   assign rd_req_desc_8_axuser_9_axuser_f = rd_req_desc_8_axuser_9_reg[31:0];
   assign rd_req_desc_8_axuser_10_axuser_f = rd_req_desc_8_axuser_10_reg[31:0];
   assign rd_req_desc_8_axuser_11_axuser_f = rd_req_desc_8_axuser_11_reg[31:0];
   assign rd_req_desc_8_axuser_12_axuser_f = rd_req_desc_8_axuser_12_reg[31:0];
   assign rd_req_desc_8_axuser_13_axuser_f = rd_req_desc_8_axuser_13_reg[31:0];
   assign rd_req_desc_8_axuser_14_axuser_f = rd_req_desc_8_axuser_14_reg[31:0];
   assign rd_req_desc_8_axuser_15_axuser_f = rd_req_desc_8_axuser_15_reg[31:0];
   assign rd_resp_desc_8_data_offset_addr_f = rd_resp_desc_8_data_offset_reg[13:0];
   assign rd_resp_desc_8_data_size_size_f = rd_resp_desc_8_data_size_reg[31:0];
   assign rd_resp_desc_8_data_host_addr_0_addr_f = rd_resp_desc_8_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_8_data_host_addr_1_addr_f = rd_resp_desc_8_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_8_data_host_addr_2_addr_f = rd_resp_desc_8_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_8_data_host_addr_3_addr_f = rd_resp_desc_8_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_8_resp_resp_f = rd_resp_desc_8_resp_reg[4:0];
   assign rd_resp_desc_8_xid_0_xid_f = rd_resp_desc_8_xid_0_reg[31:0];
   assign rd_resp_desc_8_xid_1_xid_f = rd_resp_desc_8_xid_1_reg[31:0];
   assign rd_resp_desc_8_xid_2_xid_f = rd_resp_desc_8_xid_2_reg[31:0];
   assign rd_resp_desc_8_xid_3_xid_f = rd_resp_desc_8_xid_3_reg[31:0];
   assign rd_resp_desc_8_xuser_0_xuser_f = rd_resp_desc_8_xuser_0_reg[31:0];
   assign rd_resp_desc_8_xuser_1_xuser_f = rd_resp_desc_8_xuser_1_reg[31:0];
   assign rd_resp_desc_8_xuser_2_xuser_f = rd_resp_desc_8_xuser_2_reg[31:0];
   assign rd_resp_desc_8_xuser_3_xuser_f = rd_resp_desc_8_xuser_3_reg[31:0];
   assign rd_resp_desc_8_xuser_4_xuser_f = rd_resp_desc_8_xuser_4_reg[31:0];
   assign rd_resp_desc_8_xuser_5_xuser_f = rd_resp_desc_8_xuser_5_reg[31:0];
   assign rd_resp_desc_8_xuser_6_xuser_f = rd_resp_desc_8_xuser_6_reg[31:0];
   assign rd_resp_desc_8_xuser_7_xuser_f = rd_resp_desc_8_xuser_7_reg[31:0];
   assign rd_resp_desc_8_xuser_8_xuser_f = rd_resp_desc_8_xuser_8_reg[31:0];
   assign rd_resp_desc_8_xuser_9_xuser_f = rd_resp_desc_8_xuser_9_reg[31:0];
   assign rd_resp_desc_8_xuser_10_xuser_f = rd_resp_desc_8_xuser_10_reg[31:0];
   assign rd_resp_desc_8_xuser_11_xuser_f = rd_resp_desc_8_xuser_11_reg[31:0];
   assign rd_resp_desc_8_xuser_12_xuser_f = rd_resp_desc_8_xuser_12_reg[31:0];
   assign rd_resp_desc_8_xuser_13_xuser_f = rd_resp_desc_8_xuser_13_reg[31:0];
   assign rd_resp_desc_8_xuser_14_xuser_f = rd_resp_desc_8_xuser_14_reg[31:0];
   assign rd_resp_desc_8_xuser_15_xuser_f = rd_resp_desc_8_xuser_15_reg[31:0];
   assign wr_req_desc_8_txn_type_wr_strb_f = wr_req_desc_8_txn_type_reg[1];
   assign wr_req_desc_8_size_txn_size_f = wr_req_desc_8_size_reg[31:0];
   assign wr_req_desc_8_data_offset_addr_f = wr_req_desc_8_data_offset_reg[13:0];
   assign wr_req_desc_8_data_host_addr_0_addr_f = wr_req_desc_8_data_host_addr_0_reg[31:0];
   assign wr_req_desc_8_data_host_addr_1_addr_f = wr_req_desc_8_data_host_addr_1_reg[31:0];
   assign wr_req_desc_8_data_host_addr_2_addr_f = wr_req_desc_8_data_host_addr_2_reg[31:0];
   assign wr_req_desc_8_data_host_addr_3_addr_f = wr_req_desc_8_data_host_addr_3_reg[31:0];
   assign wr_req_desc_8_wstrb_host_addr_0_addr_f = wr_req_desc_8_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_8_wstrb_host_addr_1_addr_f = wr_req_desc_8_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_8_wstrb_host_addr_2_addr_f = wr_req_desc_8_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_8_wstrb_host_addr_3_addr_f = wr_req_desc_8_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_8_axsize_axsize_f = wr_req_desc_8_axsize_reg[2:0];
   assign wr_req_desc_8_attr_axsnoop_f = wr_req_desc_8_attr_reg[27:24];
   assign wr_req_desc_8_attr_axdomain_f = wr_req_desc_8_attr_reg[23:22];
   assign wr_req_desc_8_attr_axbar_f = wr_req_desc_8_attr_reg[21:20];
   assign wr_req_desc_8_attr_awunique_f = wr_req_desc_8_attr_reg[19];
   assign wr_req_desc_8_attr_axregion_f = wr_req_desc_8_attr_reg[18:15];
   assign wr_req_desc_8_attr_axqos_f = wr_req_desc_8_attr_reg[14:11];
   assign wr_req_desc_8_attr_axprot_f = wr_req_desc_8_attr_reg[10:8];
   assign wr_req_desc_8_attr_axcache_f = wr_req_desc_8_attr_reg[7:4];
   assign wr_req_desc_8_attr_axlock_f = wr_req_desc_8_attr_reg[2];
   assign wr_req_desc_8_attr_axburst_f = wr_req_desc_8_attr_reg[1:0];
   assign wr_req_desc_8_axaddr_0_addr_f = wr_req_desc_8_axaddr_0_reg[31:0];
   assign wr_req_desc_8_axaddr_1_addr_f = wr_req_desc_8_axaddr_1_reg[31:0];
   assign wr_req_desc_8_axaddr_2_addr_f = wr_req_desc_8_axaddr_2_reg[31:0];
   assign wr_req_desc_8_axaddr_3_addr_f = wr_req_desc_8_axaddr_3_reg[31:0];
   assign wr_req_desc_8_axid_0_axid_f = wr_req_desc_8_axid_0_reg[31:0];
   assign wr_req_desc_8_axid_1_axid_f = wr_req_desc_8_axid_1_reg[31:0];
   assign wr_req_desc_8_axid_2_axid_f = wr_req_desc_8_axid_2_reg[31:0];
   assign wr_req_desc_8_axid_3_axid_f = wr_req_desc_8_axid_3_reg[31:0];
   assign wr_req_desc_8_axuser_0_axuser_f = wr_req_desc_8_axuser_0_reg[31:0];
   assign wr_req_desc_8_axuser_1_axuser_f = wr_req_desc_8_axuser_1_reg[31:0];
   assign wr_req_desc_8_axuser_2_axuser_f = wr_req_desc_8_axuser_2_reg[31:0];
   assign wr_req_desc_8_axuser_3_axuser_f = wr_req_desc_8_axuser_3_reg[31:0];
   assign wr_req_desc_8_axuser_4_axuser_f = wr_req_desc_8_axuser_4_reg[31:0];
   assign wr_req_desc_8_axuser_5_axuser_f = wr_req_desc_8_axuser_5_reg[31:0];
   assign wr_req_desc_8_axuser_6_axuser_f = wr_req_desc_8_axuser_6_reg[31:0];
   assign wr_req_desc_8_axuser_7_axuser_f = wr_req_desc_8_axuser_7_reg[31:0];
   assign wr_req_desc_8_axuser_8_axuser_f = wr_req_desc_8_axuser_8_reg[31:0];
   assign wr_req_desc_8_axuser_9_axuser_f = wr_req_desc_8_axuser_9_reg[31:0];
   assign wr_req_desc_8_axuser_10_axuser_f = wr_req_desc_8_axuser_10_reg[31:0];
   assign wr_req_desc_8_axuser_11_axuser_f = wr_req_desc_8_axuser_11_reg[31:0];
   assign wr_req_desc_8_axuser_12_axuser_f = wr_req_desc_8_axuser_12_reg[31:0];
   assign wr_req_desc_8_axuser_13_axuser_f = wr_req_desc_8_axuser_13_reg[31:0];
   assign wr_req_desc_8_axuser_14_axuser_f = wr_req_desc_8_axuser_14_reg[31:0];
   assign wr_req_desc_8_axuser_15_axuser_f = wr_req_desc_8_axuser_15_reg[31:0];
   assign wr_req_desc_8_wuser_0_wuser_f = wr_req_desc_8_wuser_0_reg[31:0];
   assign wr_req_desc_8_wuser_1_wuser_f = wr_req_desc_8_wuser_1_reg[31:0];
   assign wr_req_desc_8_wuser_2_wuser_f = wr_req_desc_8_wuser_2_reg[31:0];
   assign wr_req_desc_8_wuser_3_wuser_f = wr_req_desc_8_wuser_3_reg[31:0];
   assign wr_req_desc_8_wuser_4_wuser_f = wr_req_desc_8_wuser_4_reg[31:0];
   assign wr_req_desc_8_wuser_5_wuser_f = wr_req_desc_8_wuser_5_reg[31:0];
   assign wr_req_desc_8_wuser_6_wuser_f = wr_req_desc_8_wuser_6_reg[31:0];
   assign wr_req_desc_8_wuser_7_wuser_f = wr_req_desc_8_wuser_7_reg[31:0];
   assign wr_req_desc_8_wuser_8_wuser_f = wr_req_desc_8_wuser_8_reg[31:0];
   assign wr_req_desc_8_wuser_9_wuser_f = wr_req_desc_8_wuser_9_reg[31:0];
   assign wr_req_desc_8_wuser_10_wuser_f = wr_req_desc_8_wuser_10_reg[31:0];
   assign wr_req_desc_8_wuser_11_wuser_f = wr_req_desc_8_wuser_11_reg[31:0];
   assign wr_req_desc_8_wuser_12_wuser_f = wr_req_desc_8_wuser_12_reg[31:0];
   assign wr_req_desc_8_wuser_13_wuser_f = wr_req_desc_8_wuser_13_reg[31:0];
   assign wr_req_desc_8_wuser_14_wuser_f = wr_req_desc_8_wuser_14_reg[31:0];
   assign wr_req_desc_8_wuser_15_wuser_f = wr_req_desc_8_wuser_15_reg[31:0];
   assign wr_resp_desc_8_resp_resp_f = wr_resp_desc_8_resp_reg[4:0];
   assign wr_resp_desc_8_xid_0_xid_f = wr_resp_desc_8_xid_0_reg[31:0];
   assign wr_resp_desc_8_xid_1_xid_f = wr_resp_desc_8_xid_1_reg[31:0];
   assign wr_resp_desc_8_xid_2_xid_f = wr_resp_desc_8_xid_2_reg[31:0];
   assign wr_resp_desc_8_xid_3_xid_f = wr_resp_desc_8_xid_3_reg[31:0];
   assign wr_resp_desc_8_xuser_0_xuser_f = wr_resp_desc_8_xuser_0_reg[31:0];
   assign wr_resp_desc_8_xuser_1_xuser_f = wr_resp_desc_8_xuser_1_reg[31:0];
   assign wr_resp_desc_8_xuser_2_xuser_f = wr_resp_desc_8_xuser_2_reg[31:0];
   assign wr_resp_desc_8_xuser_3_xuser_f = wr_resp_desc_8_xuser_3_reg[31:0];
   assign wr_resp_desc_8_xuser_4_xuser_f = wr_resp_desc_8_xuser_4_reg[31:0];
   assign wr_resp_desc_8_xuser_5_xuser_f = wr_resp_desc_8_xuser_5_reg[31:0];
   assign wr_resp_desc_8_xuser_6_xuser_f = wr_resp_desc_8_xuser_6_reg[31:0];
   assign wr_resp_desc_8_xuser_7_xuser_f = wr_resp_desc_8_xuser_7_reg[31:0];
   assign wr_resp_desc_8_xuser_8_xuser_f = wr_resp_desc_8_xuser_8_reg[31:0];
   assign wr_resp_desc_8_xuser_9_xuser_f = wr_resp_desc_8_xuser_9_reg[31:0];
   assign wr_resp_desc_8_xuser_10_xuser_f = wr_resp_desc_8_xuser_10_reg[31:0];
   assign wr_resp_desc_8_xuser_11_xuser_f = wr_resp_desc_8_xuser_11_reg[31:0];
   assign wr_resp_desc_8_xuser_12_xuser_f = wr_resp_desc_8_xuser_12_reg[31:0];
   assign wr_resp_desc_8_xuser_13_xuser_f = wr_resp_desc_8_xuser_13_reg[31:0];
   assign wr_resp_desc_8_xuser_14_xuser_f = wr_resp_desc_8_xuser_14_reg[31:0];
   assign wr_resp_desc_8_xuser_15_xuser_f = wr_resp_desc_8_xuser_15_reg[31:0];
   assign sn_req_desc_8_attr_acsnoop_f = sn_req_desc_8_attr_reg[27:24];
   assign sn_req_desc_8_attr_acprot_f = sn_req_desc_8_attr_reg[10:8];
   assign sn_req_desc_8_acaddr_0_addr_f = sn_req_desc_8_acaddr_0_reg[31:0];
   assign sn_req_desc_8_acaddr_1_addr_f = sn_req_desc_8_acaddr_1_reg[31:0];
   assign sn_req_desc_8_acaddr_2_addr_f = sn_req_desc_8_acaddr_2_reg[31:0];
   assign sn_req_desc_8_acaddr_3_addr_f = sn_req_desc_8_acaddr_3_reg[31:0];
   assign sn_resp_desc_8_resp_resp_f = sn_resp_desc_8_resp_reg[4:0];
   assign rd_req_desc_9_size_txn_size_f = rd_req_desc_9_size_reg[31:0];
   assign rd_req_desc_9_axsize_axsize_f = rd_req_desc_9_axsize_reg[2:0];
   assign rd_req_desc_9_attr_axsnoop_f = rd_req_desc_9_attr_reg[27:24];
   assign rd_req_desc_9_attr_axdomain_f = rd_req_desc_9_attr_reg[23:22];
   assign rd_req_desc_9_attr_axbar_f = rd_req_desc_9_attr_reg[21:20];
   assign rd_req_desc_9_attr_axregion_f = rd_req_desc_9_attr_reg[18:15];
   assign rd_req_desc_9_attr_axqos_f = rd_req_desc_9_attr_reg[14:11];
   assign rd_req_desc_9_attr_axprot_f = rd_req_desc_9_attr_reg[10:8];
   assign rd_req_desc_9_attr_axcache_f = rd_req_desc_9_attr_reg[7:4];
   assign rd_req_desc_9_attr_axlock_f = rd_req_desc_9_attr_reg[2];
   assign rd_req_desc_9_attr_axburst_f = rd_req_desc_9_attr_reg[1:0];
   assign rd_req_desc_9_axaddr_0_addr_f = rd_req_desc_9_axaddr_0_reg[31:0];
   assign rd_req_desc_9_axaddr_1_addr_f = rd_req_desc_9_axaddr_1_reg[31:0];
   assign rd_req_desc_9_axaddr_2_addr_f = rd_req_desc_9_axaddr_2_reg[31:0];
   assign rd_req_desc_9_axaddr_3_addr_f = rd_req_desc_9_axaddr_3_reg[31:0];
   assign rd_req_desc_9_axid_0_axid_f = rd_req_desc_9_axid_0_reg[31:0];
   assign rd_req_desc_9_axid_1_axid_f = rd_req_desc_9_axid_1_reg[31:0];
   assign rd_req_desc_9_axid_2_axid_f = rd_req_desc_9_axid_2_reg[31:0];
   assign rd_req_desc_9_axid_3_axid_f = rd_req_desc_9_axid_3_reg[31:0];
   assign rd_req_desc_9_axuser_0_axuser_f = rd_req_desc_9_axuser_0_reg[31:0];
   assign rd_req_desc_9_axuser_1_axuser_f = rd_req_desc_9_axuser_1_reg[31:0];
   assign rd_req_desc_9_axuser_2_axuser_f = rd_req_desc_9_axuser_2_reg[31:0];
   assign rd_req_desc_9_axuser_3_axuser_f = rd_req_desc_9_axuser_3_reg[31:0];
   assign rd_req_desc_9_axuser_4_axuser_f = rd_req_desc_9_axuser_4_reg[31:0];
   assign rd_req_desc_9_axuser_5_axuser_f = rd_req_desc_9_axuser_5_reg[31:0];
   assign rd_req_desc_9_axuser_6_axuser_f = rd_req_desc_9_axuser_6_reg[31:0];
   assign rd_req_desc_9_axuser_7_axuser_f = rd_req_desc_9_axuser_7_reg[31:0];
   assign rd_req_desc_9_axuser_8_axuser_f = rd_req_desc_9_axuser_8_reg[31:0];
   assign rd_req_desc_9_axuser_9_axuser_f = rd_req_desc_9_axuser_9_reg[31:0];
   assign rd_req_desc_9_axuser_10_axuser_f = rd_req_desc_9_axuser_10_reg[31:0];
   assign rd_req_desc_9_axuser_11_axuser_f = rd_req_desc_9_axuser_11_reg[31:0];
   assign rd_req_desc_9_axuser_12_axuser_f = rd_req_desc_9_axuser_12_reg[31:0];
   assign rd_req_desc_9_axuser_13_axuser_f = rd_req_desc_9_axuser_13_reg[31:0];
   assign rd_req_desc_9_axuser_14_axuser_f = rd_req_desc_9_axuser_14_reg[31:0];
   assign rd_req_desc_9_axuser_15_axuser_f = rd_req_desc_9_axuser_15_reg[31:0];
   assign rd_resp_desc_9_data_offset_addr_f = rd_resp_desc_9_data_offset_reg[13:0];
   assign rd_resp_desc_9_data_size_size_f = rd_resp_desc_9_data_size_reg[31:0];
   assign rd_resp_desc_9_data_host_addr_0_addr_f = rd_resp_desc_9_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_9_data_host_addr_1_addr_f = rd_resp_desc_9_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_9_data_host_addr_2_addr_f = rd_resp_desc_9_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_9_data_host_addr_3_addr_f = rd_resp_desc_9_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_9_resp_resp_f = rd_resp_desc_9_resp_reg[4:0];
   assign rd_resp_desc_9_xid_0_xid_f = rd_resp_desc_9_xid_0_reg[31:0];
   assign rd_resp_desc_9_xid_1_xid_f = rd_resp_desc_9_xid_1_reg[31:0];
   assign rd_resp_desc_9_xid_2_xid_f = rd_resp_desc_9_xid_2_reg[31:0];
   assign rd_resp_desc_9_xid_3_xid_f = rd_resp_desc_9_xid_3_reg[31:0];
   assign rd_resp_desc_9_xuser_0_xuser_f = rd_resp_desc_9_xuser_0_reg[31:0];
   assign rd_resp_desc_9_xuser_1_xuser_f = rd_resp_desc_9_xuser_1_reg[31:0];
   assign rd_resp_desc_9_xuser_2_xuser_f = rd_resp_desc_9_xuser_2_reg[31:0];
   assign rd_resp_desc_9_xuser_3_xuser_f = rd_resp_desc_9_xuser_3_reg[31:0];
   assign rd_resp_desc_9_xuser_4_xuser_f = rd_resp_desc_9_xuser_4_reg[31:0];
   assign rd_resp_desc_9_xuser_5_xuser_f = rd_resp_desc_9_xuser_5_reg[31:0];
   assign rd_resp_desc_9_xuser_6_xuser_f = rd_resp_desc_9_xuser_6_reg[31:0];
   assign rd_resp_desc_9_xuser_7_xuser_f = rd_resp_desc_9_xuser_7_reg[31:0];
   assign rd_resp_desc_9_xuser_8_xuser_f = rd_resp_desc_9_xuser_8_reg[31:0];
   assign rd_resp_desc_9_xuser_9_xuser_f = rd_resp_desc_9_xuser_9_reg[31:0];
   assign rd_resp_desc_9_xuser_10_xuser_f = rd_resp_desc_9_xuser_10_reg[31:0];
   assign rd_resp_desc_9_xuser_11_xuser_f = rd_resp_desc_9_xuser_11_reg[31:0];
   assign rd_resp_desc_9_xuser_12_xuser_f = rd_resp_desc_9_xuser_12_reg[31:0];
   assign rd_resp_desc_9_xuser_13_xuser_f = rd_resp_desc_9_xuser_13_reg[31:0];
   assign rd_resp_desc_9_xuser_14_xuser_f = rd_resp_desc_9_xuser_14_reg[31:0];
   assign rd_resp_desc_9_xuser_15_xuser_f = rd_resp_desc_9_xuser_15_reg[31:0];
   assign wr_req_desc_9_txn_type_wr_strb_f = wr_req_desc_9_txn_type_reg[1];
   assign wr_req_desc_9_size_txn_size_f = wr_req_desc_9_size_reg[31:0];
   assign wr_req_desc_9_data_offset_addr_f = wr_req_desc_9_data_offset_reg[13:0];
   assign wr_req_desc_9_data_host_addr_0_addr_f = wr_req_desc_9_data_host_addr_0_reg[31:0];
   assign wr_req_desc_9_data_host_addr_1_addr_f = wr_req_desc_9_data_host_addr_1_reg[31:0];
   assign wr_req_desc_9_data_host_addr_2_addr_f = wr_req_desc_9_data_host_addr_2_reg[31:0];
   assign wr_req_desc_9_data_host_addr_3_addr_f = wr_req_desc_9_data_host_addr_3_reg[31:0];
   assign wr_req_desc_9_wstrb_host_addr_0_addr_f = wr_req_desc_9_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_9_wstrb_host_addr_1_addr_f = wr_req_desc_9_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_9_wstrb_host_addr_2_addr_f = wr_req_desc_9_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_9_wstrb_host_addr_3_addr_f = wr_req_desc_9_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_9_axsize_axsize_f = wr_req_desc_9_axsize_reg[2:0];
   assign wr_req_desc_9_attr_axsnoop_f = wr_req_desc_9_attr_reg[27:24];
   assign wr_req_desc_9_attr_axdomain_f = wr_req_desc_9_attr_reg[23:22];
   assign wr_req_desc_9_attr_axbar_f = wr_req_desc_9_attr_reg[21:20];
   assign wr_req_desc_9_attr_awunique_f = wr_req_desc_9_attr_reg[19];
   assign wr_req_desc_9_attr_axregion_f = wr_req_desc_9_attr_reg[18:15];
   assign wr_req_desc_9_attr_axqos_f = wr_req_desc_9_attr_reg[14:11];
   assign wr_req_desc_9_attr_axprot_f = wr_req_desc_9_attr_reg[10:8];
   assign wr_req_desc_9_attr_axcache_f = wr_req_desc_9_attr_reg[7:4];
   assign wr_req_desc_9_attr_axlock_f = wr_req_desc_9_attr_reg[2];
   assign wr_req_desc_9_attr_axburst_f = wr_req_desc_9_attr_reg[1:0];
   assign wr_req_desc_9_axaddr_0_addr_f = wr_req_desc_9_axaddr_0_reg[31:0];
   assign wr_req_desc_9_axaddr_1_addr_f = wr_req_desc_9_axaddr_1_reg[31:0];
   assign wr_req_desc_9_axaddr_2_addr_f = wr_req_desc_9_axaddr_2_reg[31:0];
   assign wr_req_desc_9_axaddr_3_addr_f = wr_req_desc_9_axaddr_3_reg[31:0];
   assign wr_req_desc_9_axid_0_axid_f = wr_req_desc_9_axid_0_reg[31:0];
   assign wr_req_desc_9_axid_1_axid_f = wr_req_desc_9_axid_1_reg[31:0];
   assign wr_req_desc_9_axid_2_axid_f = wr_req_desc_9_axid_2_reg[31:0];
   assign wr_req_desc_9_axid_3_axid_f = wr_req_desc_9_axid_3_reg[31:0];
   assign wr_req_desc_9_axuser_0_axuser_f = wr_req_desc_9_axuser_0_reg[31:0];
   assign wr_req_desc_9_axuser_1_axuser_f = wr_req_desc_9_axuser_1_reg[31:0];
   assign wr_req_desc_9_axuser_2_axuser_f = wr_req_desc_9_axuser_2_reg[31:0];
   assign wr_req_desc_9_axuser_3_axuser_f = wr_req_desc_9_axuser_3_reg[31:0];
   assign wr_req_desc_9_axuser_4_axuser_f = wr_req_desc_9_axuser_4_reg[31:0];
   assign wr_req_desc_9_axuser_5_axuser_f = wr_req_desc_9_axuser_5_reg[31:0];
   assign wr_req_desc_9_axuser_6_axuser_f = wr_req_desc_9_axuser_6_reg[31:0];
   assign wr_req_desc_9_axuser_7_axuser_f = wr_req_desc_9_axuser_7_reg[31:0];
   assign wr_req_desc_9_axuser_8_axuser_f = wr_req_desc_9_axuser_8_reg[31:0];
   assign wr_req_desc_9_axuser_9_axuser_f = wr_req_desc_9_axuser_9_reg[31:0];
   assign wr_req_desc_9_axuser_10_axuser_f = wr_req_desc_9_axuser_10_reg[31:0];
   assign wr_req_desc_9_axuser_11_axuser_f = wr_req_desc_9_axuser_11_reg[31:0];
   assign wr_req_desc_9_axuser_12_axuser_f = wr_req_desc_9_axuser_12_reg[31:0];
   assign wr_req_desc_9_axuser_13_axuser_f = wr_req_desc_9_axuser_13_reg[31:0];
   assign wr_req_desc_9_axuser_14_axuser_f = wr_req_desc_9_axuser_14_reg[31:0];
   assign wr_req_desc_9_axuser_15_axuser_f = wr_req_desc_9_axuser_15_reg[31:0];
   assign wr_req_desc_9_wuser_0_wuser_f = wr_req_desc_9_wuser_0_reg[31:0];
   assign wr_req_desc_9_wuser_1_wuser_f = wr_req_desc_9_wuser_1_reg[31:0];
   assign wr_req_desc_9_wuser_2_wuser_f = wr_req_desc_9_wuser_2_reg[31:0];
   assign wr_req_desc_9_wuser_3_wuser_f = wr_req_desc_9_wuser_3_reg[31:0];
   assign wr_req_desc_9_wuser_4_wuser_f = wr_req_desc_9_wuser_4_reg[31:0];
   assign wr_req_desc_9_wuser_5_wuser_f = wr_req_desc_9_wuser_5_reg[31:0];
   assign wr_req_desc_9_wuser_6_wuser_f = wr_req_desc_9_wuser_6_reg[31:0];
   assign wr_req_desc_9_wuser_7_wuser_f = wr_req_desc_9_wuser_7_reg[31:0];
   assign wr_req_desc_9_wuser_8_wuser_f = wr_req_desc_9_wuser_8_reg[31:0];
   assign wr_req_desc_9_wuser_9_wuser_f = wr_req_desc_9_wuser_9_reg[31:0];
   assign wr_req_desc_9_wuser_10_wuser_f = wr_req_desc_9_wuser_10_reg[31:0];
   assign wr_req_desc_9_wuser_11_wuser_f = wr_req_desc_9_wuser_11_reg[31:0];
   assign wr_req_desc_9_wuser_12_wuser_f = wr_req_desc_9_wuser_12_reg[31:0];
   assign wr_req_desc_9_wuser_13_wuser_f = wr_req_desc_9_wuser_13_reg[31:0];
   assign wr_req_desc_9_wuser_14_wuser_f = wr_req_desc_9_wuser_14_reg[31:0];
   assign wr_req_desc_9_wuser_15_wuser_f = wr_req_desc_9_wuser_15_reg[31:0];
   assign wr_resp_desc_9_resp_resp_f = wr_resp_desc_9_resp_reg[4:0];
   assign wr_resp_desc_9_xid_0_xid_f = wr_resp_desc_9_xid_0_reg[31:0];
   assign wr_resp_desc_9_xid_1_xid_f = wr_resp_desc_9_xid_1_reg[31:0];
   assign wr_resp_desc_9_xid_2_xid_f = wr_resp_desc_9_xid_2_reg[31:0];
   assign wr_resp_desc_9_xid_3_xid_f = wr_resp_desc_9_xid_3_reg[31:0];
   assign wr_resp_desc_9_xuser_0_xuser_f = wr_resp_desc_9_xuser_0_reg[31:0];
   assign wr_resp_desc_9_xuser_1_xuser_f = wr_resp_desc_9_xuser_1_reg[31:0];
   assign wr_resp_desc_9_xuser_2_xuser_f = wr_resp_desc_9_xuser_2_reg[31:0];
   assign wr_resp_desc_9_xuser_3_xuser_f = wr_resp_desc_9_xuser_3_reg[31:0];
   assign wr_resp_desc_9_xuser_4_xuser_f = wr_resp_desc_9_xuser_4_reg[31:0];
   assign wr_resp_desc_9_xuser_5_xuser_f = wr_resp_desc_9_xuser_5_reg[31:0];
   assign wr_resp_desc_9_xuser_6_xuser_f = wr_resp_desc_9_xuser_6_reg[31:0];
   assign wr_resp_desc_9_xuser_7_xuser_f = wr_resp_desc_9_xuser_7_reg[31:0];
   assign wr_resp_desc_9_xuser_8_xuser_f = wr_resp_desc_9_xuser_8_reg[31:0];
   assign wr_resp_desc_9_xuser_9_xuser_f = wr_resp_desc_9_xuser_9_reg[31:0];
   assign wr_resp_desc_9_xuser_10_xuser_f = wr_resp_desc_9_xuser_10_reg[31:0];
   assign wr_resp_desc_9_xuser_11_xuser_f = wr_resp_desc_9_xuser_11_reg[31:0];
   assign wr_resp_desc_9_xuser_12_xuser_f = wr_resp_desc_9_xuser_12_reg[31:0];
   assign wr_resp_desc_9_xuser_13_xuser_f = wr_resp_desc_9_xuser_13_reg[31:0];
   assign wr_resp_desc_9_xuser_14_xuser_f = wr_resp_desc_9_xuser_14_reg[31:0];
   assign wr_resp_desc_9_xuser_15_xuser_f = wr_resp_desc_9_xuser_15_reg[31:0];
   assign sn_req_desc_9_attr_acsnoop_f = sn_req_desc_9_attr_reg[27:24];
   assign sn_req_desc_9_attr_acprot_f = sn_req_desc_9_attr_reg[10:8];
   assign sn_req_desc_9_acaddr_0_addr_f = sn_req_desc_9_acaddr_0_reg[31:0];
   assign sn_req_desc_9_acaddr_1_addr_f = sn_req_desc_9_acaddr_1_reg[31:0];
   assign sn_req_desc_9_acaddr_2_addr_f = sn_req_desc_9_acaddr_2_reg[31:0];
   assign sn_req_desc_9_acaddr_3_addr_f = sn_req_desc_9_acaddr_3_reg[31:0];
   assign sn_resp_desc_9_resp_resp_f = sn_resp_desc_9_resp_reg[4:0];
   assign rd_req_desc_a_size_txn_size_f = rd_req_desc_a_size_reg[31:0];
   assign rd_req_desc_a_axsize_axsize_f = rd_req_desc_a_axsize_reg[2:0];
   assign rd_req_desc_a_attr_axsnoop_f = rd_req_desc_a_attr_reg[27:24];
   assign rd_req_desc_a_attr_axdomain_f = rd_req_desc_a_attr_reg[23:22];
   assign rd_req_desc_a_attr_axbar_f = rd_req_desc_a_attr_reg[21:20];
   assign rd_req_desc_a_attr_axregion_f = rd_req_desc_a_attr_reg[18:15];
   assign rd_req_desc_a_attr_axqos_f = rd_req_desc_a_attr_reg[14:11];
   assign rd_req_desc_a_attr_axprot_f = rd_req_desc_a_attr_reg[10:8];
   assign rd_req_desc_a_attr_axcache_f = rd_req_desc_a_attr_reg[7:4];
   assign rd_req_desc_a_attr_axlock_f = rd_req_desc_a_attr_reg[2];
   assign rd_req_desc_a_attr_axburst_f = rd_req_desc_a_attr_reg[1:0];
   assign rd_req_desc_a_axaddr_0_addr_f = rd_req_desc_a_axaddr_0_reg[31:0];
   assign rd_req_desc_a_axaddr_1_addr_f = rd_req_desc_a_axaddr_1_reg[31:0];
   assign rd_req_desc_a_axaddr_2_addr_f = rd_req_desc_a_axaddr_2_reg[31:0];
   assign rd_req_desc_a_axaddr_3_addr_f = rd_req_desc_a_axaddr_3_reg[31:0];
   assign rd_req_desc_a_axid_0_axid_f = rd_req_desc_a_axid_0_reg[31:0];
   assign rd_req_desc_a_axid_1_axid_f = rd_req_desc_a_axid_1_reg[31:0];
   assign rd_req_desc_a_axid_2_axid_f = rd_req_desc_a_axid_2_reg[31:0];
   assign rd_req_desc_a_axid_3_axid_f = rd_req_desc_a_axid_3_reg[31:0];
   assign rd_req_desc_a_axuser_0_axuser_f = rd_req_desc_a_axuser_0_reg[31:0];
   assign rd_req_desc_a_axuser_1_axuser_f = rd_req_desc_a_axuser_1_reg[31:0];
   assign rd_req_desc_a_axuser_2_axuser_f = rd_req_desc_a_axuser_2_reg[31:0];
   assign rd_req_desc_a_axuser_3_axuser_f = rd_req_desc_a_axuser_3_reg[31:0];
   assign rd_req_desc_a_axuser_4_axuser_f = rd_req_desc_a_axuser_4_reg[31:0];
   assign rd_req_desc_a_axuser_5_axuser_f = rd_req_desc_a_axuser_5_reg[31:0];
   assign rd_req_desc_a_axuser_6_axuser_f = rd_req_desc_a_axuser_6_reg[31:0];
   assign rd_req_desc_a_axuser_7_axuser_f = rd_req_desc_a_axuser_7_reg[31:0];
   assign rd_req_desc_a_axuser_8_axuser_f = rd_req_desc_a_axuser_8_reg[31:0];
   assign rd_req_desc_a_axuser_9_axuser_f = rd_req_desc_a_axuser_9_reg[31:0];
   assign rd_req_desc_a_axuser_10_axuser_f = rd_req_desc_a_axuser_10_reg[31:0];
   assign rd_req_desc_a_axuser_11_axuser_f = rd_req_desc_a_axuser_11_reg[31:0];
   assign rd_req_desc_a_axuser_12_axuser_f = rd_req_desc_a_axuser_12_reg[31:0];
   assign rd_req_desc_a_axuser_13_axuser_f = rd_req_desc_a_axuser_13_reg[31:0];
   assign rd_req_desc_a_axuser_14_axuser_f = rd_req_desc_a_axuser_14_reg[31:0];
   assign rd_req_desc_a_axuser_15_axuser_f = rd_req_desc_a_axuser_15_reg[31:0];
   assign rd_resp_desc_a_data_offset_addr_f = rd_resp_desc_a_data_offset_reg[13:0];
   assign rd_resp_desc_a_data_size_size_f = rd_resp_desc_a_data_size_reg[31:0];
   assign rd_resp_desc_a_data_host_addr_0_addr_f = rd_resp_desc_a_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_a_data_host_addr_1_addr_f = rd_resp_desc_a_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_a_data_host_addr_2_addr_f = rd_resp_desc_a_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_a_data_host_addr_3_addr_f = rd_resp_desc_a_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_a_resp_resp_f = rd_resp_desc_a_resp_reg[4:0];
   assign rd_resp_desc_a_xid_0_xid_f = rd_resp_desc_a_xid_0_reg[31:0];
   assign rd_resp_desc_a_xid_1_xid_f = rd_resp_desc_a_xid_1_reg[31:0];
   assign rd_resp_desc_a_xid_2_xid_f = rd_resp_desc_a_xid_2_reg[31:0];
   assign rd_resp_desc_a_xid_3_xid_f = rd_resp_desc_a_xid_3_reg[31:0];
   assign rd_resp_desc_a_xuser_0_xuser_f = rd_resp_desc_a_xuser_0_reg[31:0];
   assign rd_resp_desc_a_xuser_1_xuser_f = rd_resp_desc_a_xuser_1_reg[31:0];
   assign rd_resp_desc_a_xuser_2_xuser_f = rd_resp_desc_a_xuser_2_reg[31:0];
   assign rd_resp_desc_a_xuser_3_xuser_f = rd_resp_desc_a_xuser_3_reg[31:0];
   assign rd_resp_desc_a_xuser_4_xuser_f = rd_resp_desc_a_xuser_4_reg[31:0];
   assign rd_resp_desc_a_xuser_5_xuser_f = rd_resp_desc_a_xuser_5_reg[31:0];
   assign rd_resp_desc_a_xuser_6_xuser_f = rd_resp_desc_a_xuser_6_reg[31:0];
   assign rd_resp_desc_a_xuser_7_xuser_f = rd_resp_desc_a_xuser_7_reg[31:0];
   assign rd_resp_desc_a_xuser_8_xuser_f = rd_resp_desc_a_xuser_8_reg[31:0];
   assign rd_resp_desc_a_xuser_9_xuser_f = rd_resp_desc_a_xuser_9_reg[31:0];
   assign rd_resp_desc_a_xuser_10_xuser_f = rd_resp_desc_a_xuser_10_reg[31:0];
   assign rd_resp_desc_a_xuser_11_xuser_f = rd_resp_desc_a_xuser_11_reg[31:0];
   assign rd_resp_desc_a_xuser_12_xuser_f = rd_resp_desc_a_xuser_12_reg[31:0];
   assign rd_resp_desc_a_xuser_13_xuser_f = rd_resp_desc_a_xuser_13_reg[31:0];
   assign rd_resp_desc_a_xuser_14_xuser_f = rd_resp_desc_a_xuser_14_reg[31:0];
   assign rd_resp_desc_a_xuser_15_xuser_f = rd_resp_desc_a_xuser_15_reg[31:0];
   assign wr_req_desc_a_txn_type_wr_strb_f = wr_req_desc_a_txn_type_reg[1];
   assign wr_req_desc_a_size_txn_size_f = wr_req_desc_a_size_reg[31:0];
   assign wr_req_desc_a_data_offset_addr_f = wr_req_desc_a_data_offset_reg[13:0];
   assign wr_req_desc_a_data_host_addr_0_addr_f = wr_req_desc_a_data_host_addr_0_reg[31:0];
   assign wr_req_desc_a_data_host_addr_1_addr_f = wr_req_desc_a_data_host_addr_1_reg[31:0];
   assign wr_req_desc_a_data_host_addr_2_addr_f = wr_req_desc_a_data_host_addr_2_reg[31:0];
   assign wr_req_desc_a_data_host_addr_3_addr_f = wr_req_desc_a_data_host_addr_3_reg[31:0];
   assign wr_req_desc_a_wstrb_host_addr_0_addr_f = wr_req_desc_a_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_a_wstrb_host_addr_1_addr_f = wr_req_desc_a_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_a_wstrb_host_addr_2_addr_f = wr_req_desc_a_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_a_wstrb_host_addr_3_addr_f = wr_req_desc_a_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_a_axsize_axsize_f = wr_req_desc_a_axsize_reg[2:0];
   assign wr_req_desc_a_attr_axsnoop_f = wr_req_desc_a_attr_reg[27:24];
   assign wr_req_desc_a_attr_axdomain_f = wr_req_desc_a_attr_reg[23:22];
   assign wr_req_desc_a_attr_axbar_f = wr_req_desc_a_attr_reg[21:20];
   assign wr_req_desc_a_attr_awunique_f = wr_req_desc_a_attr_reg[19];
   assign wr_req_desc_a_attr_axregion_f = wr_req_desc_a_attr_reg[18:15];
   assign wr_req_desc_a_attr_axqos_f = wr_req_desc_a_attr_reg[14:11];
   assign wr_req_desc_a_attr_axprot_f = wr_req_desc_a_attr_reg[10:8];
   assign wr_req_desc_a_attr_axcache_f = wr_req_desc_a_attr_reg[7:4];
   assign wr_req_desc_a_attr_axlock_f = wr_req_desc_a_attr_reg[2];
   assign wr_req_desc_a_attr_axburst_f = wr_req_desc_a_attr_reg[1:0];
   assign wr_req_desc_a_axaddr_0_addr_f = wr_req_desc_a_axaddr_0_reg[31:0];
   assign wr_req_desc_a_axaddr_1_addr_f = wr_req_desc_a_axaddr_1_reg[31:0];
   assign wr_req_desc_a_axaddr_2_addr_f = wr_req_desc_a_axaddr_2_reg[31:0];
   assign wr_req_desc_a_axaddr_3_addr_f = wr_req_desc_a_axaddr_3_reg[31:0];
   assign wr_req_desc_a_axid_0_axid_f = wr_req_desc_a_axid_0_reg[31:0];
   assign wr_req_desc_a_axid_1_axid_f = wr_req_desc_a_axid_1_reg[31:0];
   assign wr_req_desc_a_axid_2_axid_f = wr_req_desc_a_axid_2_reg[31:0];
   assign wr_req_desc_a_axid_3_axid_f = wr_req_desc_a_axid_3_reg[31:0];
   assign wr_req_desc_a_axuser_0_axuser_f = wr_req_desc_a_axuser_0_reg[31:0];
   assign wr_req_desc_a_axuser_1_axuser_f = wr_req_desc_a_axuser_1_reg[31:0];
   assign wr_req_desc_a_axuser_2_axuser_f = wr_req_desc_a_axuser_2_reg[31:0];
   assign wr_req_desc_a_axuser_3_axuser_f = wr_req_desc_a_axuser_3_reg[31:0];
   assign wr_req_desc_a_axuser_4_axuser_f = wr_req_desc_a_axuser_4_reg[31:0];
   assign wr_req_desc_a_axuser_5_axuser_f = wr_req_desc_a_axuser_5_reg[31:0];
   assign wr_req_desc_a_axuser_6_axuser_f = wr_req_desc_a_axuser_6_reg[31:0];
   assign wr_req_desc_a_axuser_7_axuser_f = wr_req_desc_a_axuser_7_reg[31:0];
   assign wr_req_desc_a_axuser_8_axuser_f = wr_req_desc_a_axuser_8_reg[31:0];
   assign wr_req_desc_a_axuser_9_axuser_f = wr_req_desc_a_axuser_9_reg[31:0];
   assign wr_req_desc_a_axuser_10_axuser_f = wr_req_desc_a_axuser_10_reg[31:0];
   assign wr_req_desc_a_axuser_11_axuser_f = wr_req_desc_a_axuser_11_reg[31:0];
   assign wr_req_desc_a_axuser_12_axuser_f = wr_req_desc_a_axuser_12_reg[31:0];
   assign wr_req_desc_a_axuser_13_axuser_f = wr_req_desc_a_axuser_13_reg[31:0];
   assign wr_req_desc_a_axuser_14_axuser_f = wr_req_desc_a_axuser_14_reg[31:0];
   assign wr_req_desc_a_axuser_15_axuser_f = wr_req_desc_a_axuser_15_reg[31:0];
   assign wr_req_desc_a_wuser_0_wuser_f = wr_req_desc_a_wuser_0_reg[31:0];
   assign wr_req_desc_a_wuser_1_wuser_f = wr_req_desc_a_wuser_1_reg[31:0];
   assign wr_req_desc_a_wuser_2_wuser_f = wr_req_desc_a_wuser_2_reg[31:0];
   assign wr_req_desc_a_wuser_3_wuser_f = wr_req_desc_a_wuser_3_reg[31:0];
   assign wr_req_desc_a_wuser_4_wuser_f = wr_req_desc_a_wuser_4_reg[31:0];
   assign wr_req_desc_a_wuser_5_wuser_f = wr_req_desc_a_wuser_5_reg[31:0];
   assign wr_req_desc_a_wuser_6_wuser_f = wr_req_desc_a_wuser_6_reg[31:0];
   assign wr_req_desc_a_wuser_7_wuser_f = wr_req_desc_a_wuser_7_reg[31:0];
   assign wr_req_desc_a_wuser_8_wuser_f = wr_req_desc_a_wuser_8_reg[31:0];
   assign wr_req_desc_a_wuser_9_wuser_f = wr_req_desc_a_wuser_9_reg[31:0];
   assign wr_req_desc_a_wuser_10_wuser_f = wr_req_desc_a_wuser_10_reg[31:0];
   assign wr_req_desc_a_wuser_11_wuser_f = wr_req_desc_a_wuser_11_reg[31:0];
   assign wr_req_desc_a_wuser_12_wuser_f = wr_req_desc_a_wuser_12_reg[31:0];
   assign wr_req_desc_a_wuser_13_wuser_f = wr_req_desc_a_wuser_13_reg[31:0];
   assign wr_req_desc_a_wuser_14_wuser_f = wr_req_desc_a_wuser_14_reg[31:0];
   assign wr_req_desc_a_wuser_15_wuser_f = wr_req_desc_a_wuser_15_reg[31:0];
   assign wr_resp_desc_a_resp_resp_f = wr_resp_desc_a_resp_reg[4:0];
   assign wr_resp_desc_a_xid_0_xid_f = wr_resp_desc_a_xid_0_reg[31:0];
   assign wr_resp_desc_a_xid_1_xid_f = wr_resp_desc_a_xid_1_reg[31:0];
   assign wr_resp_desc_a_xid_2_xid_f = wr_resp_desc_a_xid_2_reg[31:0];
   assign wr_resp_desc_a_xid_3_xid_f = wr_resp_desc_a_xid_3_reg[31:0];
   assign wr_resp_desc_a_xuser_0_xuser_f = wr_resp_desc_a_xuser_0_reg[31:0];
   assign wr_resp_desc_a_xuser_1_xuser_f = wr_resp_desc_a_xuser_1_reg[31:0];
   assign wr_resp_desc_a_xuser_2_xuser_f = wr_resp_desc_a_xuser_2_reg[31:0];
   assign wr_resp_desc_a_xuser_3_xuser_f = wr_resp_desc_a_xuser_3_reg[31:0];
   assign wr_resp_desc_a_xuser_4_xuser_f = wr_resp_desc_a_xuser_4_reg[31:0];
   assign wr_resp_desc_a_xuser_5_xuser_f = wr_resp_desc_a_xuser_5_reg[31:0];
   assign wr_resp_desc_a_xuser_6_xuser_f = wr_resp_desc_a_xuser_6_reg[31:0];
   assign wr_resp_desc_a_xuser_7_xuser_f = wr_resp_desc_a_xuser_7_reg[31:0];
   assign wr_resp_desc_a_xuser_8_xuser_f = wr_resp_desc_a_xuser_8_reg[31:0];
   assign wr_resp_desc_a_xuser_9_xuser_f = wr_resp_desc_a_xuser_9_reg[31:0];
   assign wr_resp_desc_a_xuser_10_xuser_f = wr_resp_desc_a_xuser_10_reg[31:0];
   assign wr_resp_desc_a_xuser_11_xuser_f = wr_resp_desc_a_xuser_11_reg[31:0];
   assign wr_resp_desc_a_xuser_12_xuser_f = wr_resp_desc_a_xuser_12_reg[31:0];
   assign wr_resp_desc_a_xuser_13_xuser_f = wr_resp_desc_a_xuser_13_reg[31:0];
   assign wr_resp_desc_a_xuser_14_xuser_f = wr_resp_desc_a_xuser_14_reg[31:0];
   assign wr_resp_desc_a_xuser_15_xuser_f = wr_resp_desc_a_xuser_15_reg[31:0];
   assign sn_req_desc_a_attr_acsnoop_f = sn_req_desc_a_attr_reg[27:24];
   assign sn_req_desc_a_attr_acprot_f = sn_req_desc_a_attr_reg[10:8];
   assign sn_req_desc_a_acaddr_0_addr_f = sn_req_desc_a_acaddr_0_reg[31:0];
   assign sn_req_desc_a_acaddr_1_addr_f = sn_req_desc_a_acaddr_1_reg[31:0];
   assign sn_req_desc_a_acaddr_2_addr_f = sn_req_desc_a_acaddr_2_reg[31:0];
   assign sn_req_desc_a_acaddr_3_addr_f = sn_req_desc_a_acaddr_3_reg[31:0];
   assign sn_resp_desc_a_resp_resp_f = sn_resp_desc_a_resp_reg[4:0];
   assign rd_req_desc_b_size_txn_size_f = rd_req_desc_b_size_reg[31:0];
   assign rd_req_desc_b_axsize_axsize_f = rd_req_desc_b_axsize_reg[2:0];
   assign rd_req_desc_b_attr_axsnoop_f = rd_req_desc_b_attr_reg[27:24];
   assign rd_req_desc_b_attr_axdomain_f = rd_req_desc_b_attr_reg[23:22];
   assign rd_req_desc_b_attr_axbar_f = rd_req_desc_b_attr_reg[21:20];
   assign rd_req_desc_b_attr_axregion_f = rd_req_desc_b_attr_reg[18:15];
   assign rd_req_desc_b_attr_axqos_f = rd_req_desc_b_attr_reg[14:11];
   assign rd_req_desc_b_attr_axprot_f = rd_req_desc_b_attr_reg[10:8];
   assign rd_req_desc_b_attr_axcache_f = rd_req_desc_b_attr_reg[7:4];
   assign rd_req_desc_b_attr_axlock_f = rd_req_desc_b_attr_reg[2];
   assign rd_req_desc_b_attr_axburst_f = rd_req_desc_b_attr_reg[1:0];
   assign rd_req_desc_b_axaddr_0_addr_f = rd_req_desc_b_axaddr_0_reg[31:0];
   assign rd_req_desc_b_axaddr_1_addr_f = rd_req_desc_b_axaddr_1_reg[31:0];
   assign rd_req_desc_b_axaddr_2_addr_f = rd_req_desc_b_axaddr_2_reg[31:0];
   assign rd_req_desc_b_axaddr_3_addr_f = rd_req_desc_b_axaddr_3_reg[31:0];
   assign rd_req_desc_b_axid_0_axid_f = rd_req_desc_b_axid_0_reg[31:0];
   assign rd_req_desc_b_axid_1_axid_f = rd_req_desc_b_axid_1_reg[31:0];
   assign rd_req_desc_b_axid_2_axid_f = rd_req_desc_b_axid_2_reg[31:0];
   assign rd_req_desc_b_axid_3_axid_f = rd_req_desc_b_axid_3_reg[31:0];
   assign rd_req_desc_b_axuser_0_axuser_f = rd_req_desc_b_axuser_0_reg[31:0];
   assign rd_req_desc_b_axuser_1_axuser_f = rd_req_desc_b_axuser_1_reg[31:0];
   assign rd_req_desc_b_axuser_2_axuser_f = rd_req_desc_b_axuser_2_reg[31:0];
   assign rd_req_desc_b_axuser_3_axuser_f = rd_req_desc_b_axuser_3_reg[31:0];
   assign rd_req_desc_b_axuser_4_axuser_f = rd_req_desc_b_axuser_4_reg[31:0];
   assign rd_req_desc_b_axuser_5_axuser_f = rd_req_desc_b_axuser_5_reg[31:0];
   assign rd_req_desc_b_axuser_6_axuser_f = rd_req_desc_b_axuser_6_reg[31:0];
   assign rd_req_desc_b_axuser_7_axuser_f = rd_req_desc_b_axuser_7_reg[31:0];
   assign rd_req_desc_b_axuser_8_axuser_f = rd_req_desc_b_axuser_8_reg[31:0];
   assign rd_req_desc_b_axuser_9_axuser_f = rd_req_desc_b_axuser_9_reg[31:0];
   assign rd_req_desc_b_axuser_10_axuser_f = rd_req_desc_b_axuser_10_reg[31:0];
   assign rd_req_desc_b_axuser_11_axuser_f = rd_req_desc_b_axuser_11_reg[31:0];
   assign rd_req_desc_b_axuser_12_axuser_f = rd_req_desc_b_axuser_12_reg[31:0];
   assign rd_req_desc_b_axuser_13_axuser_f = rd_req_desc_b_axuser_13_reg[31:0];
   assign rd_req_desc_b_axuser_14_axuser_f = rd_req_desc_b_axuser_14_reg[31:0];
   assign rd_req_desc_b_axuser_15_axuser_f = rd_req_desc_b_axuser_15_reg[31:0];
   assign rd_resp_desc_b_data_offset_addr_f = rd_resp_desc_b_data_offset_reg[13:0];
   assign rd_resp_desc_b_data_size_size_f = rd_resp_desc_b_data_size_reg[31:0];
   assign rd_resp_desc_b_data_host_addr_0_addr_f = rd_resp_desc_b_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_b_data_host_addr_1_addr_f = rd_resp_desc_b_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_b_data_host_addr_2_addr_f = rd_resp_desc_b_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_b_data_host_addr_3_addr_f = rd_resp_desc_b_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_b_resp_resp_f = rd_resp_desc_b_resp_reg[4:0];
   assign rd_resp_desc_b_xid_0_xid_f = rd_resp_desc_b_xid_0_reg[31:0];
   assign rd_resp_desc_b_xid_1_xid_f = rd_resp_desc_b_xid_1_reg[31:0];
   assign rd_resp_desc_b_xid_2_xid_f = rd_resp_desc_b_xid_2_reg[31:0];
   assign rd_resp_desc_b_xid_3_xid_f = rd_resp_desc_b_xid_3_reg[31:0];
   assign rd_resp_desc_b_xuser_0_xuser_f = rd_resp_desc_b_xuser_0_reg[31:0];
   assign rd_resp_desc_b_xuser_1_xuser_f = rd_resp_desc_b_xuser_1_reg[31:0];
   assign rd_resp_desc_b_xuser_2_xuser_f = rd_resp_desc_b_xuser_2_reg[31:0];
   assign rd_resp_desc_b_xuser_3_xuser_f = rd_resp_desc_b_xuser_3_reg[31:0];
   assign rd_resp_desc_b_xuser_4_xuser_f = rd_resp_desc_b_xuser_4_reg[31:0];
   assign rd_resp_desc_b_xuser_5_xuser_f = rd_resp_desc_b_xuser_5_reg[31:0];
   assign rd_resp_desc_b_xuser_6_xuser_f = rd_resp_desc_b_xuser_6_reg[31:0];
   assign rd_resp_desc_b_xuser_7_xuser_f = rd_resp_desc_b_xuser_7_reg[31:0];
   assign rd_resp_desc_b_xuser_8_xuser_f = rd_resp_desc_b_xuser_8_reg[31:0];
   assign rd_resp_desc_b_xuser_9_xuser_f = rd_resp_desc_b_xuser_9_reg[31:0];
   assign rd_resp_desc_b_xuser_10_xuser_f = rd_resp_desc_b_xuser_10_reg[31:0];
   assign rd_resp_desc_b_xuser_11_xuser_f = rd_resp_desc_b_xuser_11_reg[31:0];
   assign rd_resp_desc_b_xuser_12_xuser_f = rd_resp_desc_b_xuser_12_reg[31:0];
   assign rd_resp_desc_b_xuser_13_xuser_f = rd_resp_desc_b_xuser_13_reg[31:0];
   assign rd_resp_desc_b_xuser_14_xuser_f = rd_resp_desc_b_xuser_14_reg[31:0];
   assign rd_resp_desc_b_xuser_15_xuser_f = rd_resp_desc_b_xuser_15_reg[31:0];
   assign wr_req_desc_b_txn_type_wr_strb_f = wr_req_desc_b_txn_type_reg[1];
   assign wr_req_desc_b_size_txn_size_f = wr_req_desc_b_size_reg[31:0];
   assign wr_req_desc_b_data_offset_addr_f = wr_req_desc_b_data_offset_reg[13:0];
   assign wr_req_desc_b_data_host_addr_0_addr_f = wr_req_desc_b_data_host_addr_0_reg[31:0];
   assign wr_req_desc_b_data_host_addr_1_addr_f = wr_req_desc_b_data_host_addr_1_reg[31:0];
   assign wr_req_desc_b_data_host_addr_2_addr_f = wr_req_desc_b_data_host_addr_2_reg[31:0];
   assign wr_req_desc_b_data_host_addr_3_addr_f = wr_req_desc_b_data_host_addr_3_reg[31:0];
   assign wr_req_desc_b_wstrb_host_addr_0_addr_f = wr_req_desc_b_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_b_wstrb_host_addr_1_addr_f = wr_req_desc_b_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_b_wstrb_host_addr_2_addr_f = wr_req_desc_b_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_b_wstrb_host_addr_3_addr_f = wr_req_desc_b_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_b_axsize_axsize_f = wr_req_desc_b_axsize_reg[2:0];
   assign wr_req_desc_b_attr_axsnoop_f = wr_req_desc_b_attr_reg[27:24];
   assign wr_req_desc_b_attr_axdomain_f = wr_req_desc_b_attr_reg[23:22];
   assign wr_req_desc_b_attr_axbar_f = wr_req_desc_b_attr_reg[21:20];
   assign wr_req_desc_b_attr_awunique_f = wr_req_desc_b_attr_reg[19];
   assign wr_req_desc_b_attr_axregion_f = wr_req_desc_b_attr_reg[18:15];
   assign wr_req_desc_b_attr_axqos_f = wr_req_desc_b_attr_reg[14:11];
   assign wr_req_desc_b_attr_axprot_f = wr_req_desc_b_attr_reg[10:8];
   assign wr_req_desc_b_attr_axcache_f = wr_req_desc_b_attr_reg[7:4];
   assign wr_req_desc_b_attr_axlock_f = wr_req_desc_b_attr_reg[2];
   assign wr_req_desc_b_attr_axburst_f = wr_req_desc_b_attr_reg[1:0];
   assign wr_req_desc_b_axaddr_0_addr_f = wr_req_desc_b_axaddr_0_reg[31:0];
   assign wr_req_desc_b_axaddr_1_addr_f = wr_req_desc_b_axaddr_1_reg[31:0];
   assign wr_req_desc_b_axaddr_2_addr_f = wr_req_desc_b_axaddr_2_reg[31:0];
   assign wr_req_desc_b_axaddr_3_addr_f = wr_req_desc_b_axaddr_3_reg[31:0];
   assign wr_req_desc_b_axid_0_axid_f = wr_req_desc_b_axid_0_reg[31:0];
   assign wr_req_desc_b_axid_1_axid_f = wr_req_desc_b_axid_1_reg[31:0];
   assign wr_req_desc_b_axid_2_axid_f = wr_req_desc_b_axid_2_reg[31:0];
   assign wr_req_desc_b_axid_3_axid_f = wr_req_desc_b_axid_3_reg[31:0];
   assign wr_req_desc_b_axuser_0_axuser_f = wr_req_desc_b_axuser_0_reg[31:0];
   assign wr_req_desc_b_axuser_1_axuser_f = wr_req_desc_b_axuser_1_reg[31:0];
   assign wr_req_desc_b_axuser_2_axuser_f = wr_req_desc_b_axuser_2_reg[31:0];
   assign wr_req_desc_b_axuser_3_axuser_f = wr_req_desc_b_axuser_3_reg[31:0];
   assign wr_req_desc_b_axuser_4_axuser_f = wr_req_desc_b_axuser_4_reg[31:0];
   assign wr_req_desc_b_axuser_5_axuser_f = wr_req_desc_b_axuser_5_reg[31:0];
   assign wr_req_desc_b_axuser_6_axuser_f = wr_req_desc_b_axuser_6_reg[31:0];
   assign wr_req_desc_b_axuser_7_axuser_f = wr_req_desc_b_axuser_7_reg[31:0];
   assign wr_req_desc_b_axuser_8_axuser_f = wr_req_desc_b_axuser_8_reg[31:0];
   assign wr_req_desc_b_axuser_9_axuser_f = wr_req_desc_b_axuser_9_reg[31:0];
   assign wr_req_desc_b_axuser_10_axuser_f = wr_req_desc_b_axuser_10_reg[31:0];
   assign wr_req_desc_b_axuser_11_axuser_f = wr_req_desc_b_axuser_11_reg[31:0];
   assign wr_req_desc_b_axuser_12_axuser_f = wr_req_desc_b_axuser_12_reg[31:0];
   assign wr_req_desc_b_axuser_13_axuser_f = wr_req_desc_b_axuser_13_reg[31:0];
   assign wr_req_desc_b_axuser_14_axuser_f = wr_req_desc_b_axuser_14_reg[31:0];
   assign wr_req_desc_b_axuser_15_axuser_f = wr_req_desc_b_axuser_15_reg[31:0];
   assign wr_req_desc_b_wuser_0_wuser_f = wr_req_desc_b_wuser_0_reg[31:0];
   assign wr_req_desc_b_wuser_1_wuser_f = wr_req_desc_b_wuser_1_reg[31:0];
   assign wr_req_desc_b_wuser_2_wuser_f = wr_req_desc_b_wuser_2_reg[31:0];
   assign wr_req_desc_b_wuser_3_wuser_f = wr_req_desc_b_wuser_3_reg[31:0];
   assign wr_req_desc_b_wuser_4_wuser_f = wr_req_desc_b_wuser_4_reg[31:0];
   assign wr_req_desc_b_wuser_5_wuser_f = wr_req_desc_b_wuser_5_reg[31:0];
   assign wr_req_desc_b_wuser_6_wuser_f = wr_req_desc_b_wuser_6_reg[31:0];
   assign wr_req_desc_b_wuser_7_wuser_f = wr_req_desc_b_wuser_7_reg[31:0];
   assign wr_req_desc_b_wuser_8_wuser_f = wr_req_desc_b_wuser_8_reg[31:0];
   assign wr_req_desc_b_wuser_9_wuser_f = wr_req_desc_b_wuser_9_reg[31:0];
   assign wr_req_desc_b_wuser_10_wuser_f = wr_req_desc_b_wuser_10_reg[31:0];
   assign wr_req_desc_b_wuser_11_wuser_f = wr_req_desc_b_wuser_11_reg[31:0];
   assign wr_req_desc_b_wuser_12_wuser_f = wr_req_desc_b_wuser_12_reg[31:0];
   assign wr_req_desc_b_wuser_13_wuser_f = wr_req_desc_b_wuser_13_reg[31:0];
   assign wr_req_desc_b_wuser_14_wuser_f = wr_req_desc_b_wuser_14_reg[31:0];
   assign wr_req_desc_b_wuser_15_wuser_f = wr_req_desc_b_wuser_15_reg[31:0];
   assign wr_resp_desc_b_resp_resp_f = wr_resp_desc_b_resp_reg[4:0];
   assign wr_resp_desc_b_xid_0_xid_f = wr_resp_desc_b_xid_0_reg[31:0];
   assign wr_resp_desc_b_xid_1_xid_f = wr_resp_desc_b_xid_1_reg[31:0];
   assign wr_resp_desc_b_xid_2_xid_f = wr_resp_desc_b_xid_2_reg[31:0];
   assign wr_resp_desc_b_xid_3_xid_f = wr_resp_desc_b_xid_3_reg[31:0];
   assign wr_resp_desc_b_xuser_0_xuser_f = wr_resp_desc_b_xuser_0_reg[31:0];
   assign wr_resp_desc_b_xuser_1_xuser_f = wr_resp_desc_b_xuser_1_reg[31:0];
   assign wr_resp_desc_b_xuser_2_xuser_f = wr_resp_desc_b_xuser_2_reg[31:0];
   assign wr_resp_desc_b_xuser_3_xuser_f = wr_resp_desc_b_xuser_3_reg[31:0];
   assign wr_resp_desc_b_xuser_4_xuser_f = wr_resp_desc_b_xuser_4_reg[31:0];
   assign wr_resp_desc_b_xuser_5_xuser_f = wr_resp_desc_b_xuser_5_reg[31:0];
   assign wr_resp_desc_b_xuser_6_xuser_f = wr_resp_desc_b_xuser_6_reg[31:0];
   assign wr_resp_desc_b_xuser_7_xuser_f = wr_resp_desc_b_xuser_7_reg[31:0];
   assign wr_resp_desc_b_xuser_8_xuser_f = wr_resp_desc_b_xuser_8_reg[31:0];
   assign wr_resp_desc_b_xuser_9_xuser_f = wr_resp_desc_b_xuser_9_reg[31:0];
   assign wr_resp_desc_b_xuser_10_xuser_f = wr_resp_desc_b_xuser_10_reg[31:0];
   assign wr_resp_desc_b_xuser_11_xuser_f = wr_resp_desc_b_xuser_11_reg[31:0];
   assign wr_resp_desc_b_xuser_12_xuser_f = wr_resp_desc_b_xuser_12_reg[31:0];
   assign wr_resp_desc_b_xuser_13_xuser_f = wr_resp_desc_b_xuser_13_reg[31:0];
   assign wr_resp_desc_b_xuser_14_xuser_f = wr_resp_desc_b_xuser_14_reg[31:0];
   assign wr_resp_desc_b_xuser_15_xuser_f = wr_resp_desc_b_xuser_15_reg[31:0];
   assign sn_req_desc_b_attr_acsnoop_f = sn_req_desc_b_attr_reg[27:24];
   assign sn_req_desc_b_attr_acprot_f = sn_req_desc_b_attr_reg[10:8];
   assign sn_req_desc_b_acaddr_0_addr_f = sn_req_desc_b_acaddr_0_reg[31:0];
   assign sn_req_desc_b_acaddr_1_addr_f = sn_req_desc_b_acaddr_1_reg[31:0];
   assign sn_req_desc_b_acaddr_2_addr_f = sn_req_desc_b_acaddr_2_reg[31:0];
   assign sn_req_desc_b_acaddr_3_addr_f = sn_req_desc_b_acaddr_3_reg[31:0];
   assign sn_resp_desc_b_resp_resp_f = sn_resp_desc_b_resp_reg[4:0];
   assign rd_req_desc_c_size_txn_size_f = rd_req_desc_c_size_reg[31:0];
   assign rd_req_desc_c_axsize_axsize_f = rd_req_desc_c_axsize_reg[2:0];
   assign rd_req_desc_c_attr_axsnoop_f = rd_req_desc_c_attr_reg[27:24];
   assign rd_req_desc_c_attr_axdomain_f = rd_req_desc_c_attr_reg[23:22];
   assign rd_req_desc_c_attr_axbar_f = rd_req_desc_c_attr_reg[21:20];
   assign rd_req_desc_c_attr_axregion_f = rd_req_desc_c_attr_reg[18:15];
   assign rd_req_desc_c_attr_axqos_f = rd_req_desc_c_attr_reg[14:11];
   assign rd_req_desc_c_attr_axprot_f = rd_req_desc_c_attr_reg[10:8];
   assign rd_req_desc_c_attr_axcache_f = rd_req_desc_c_attr_reg[7:4];
   assign rd_req_desc_c_attr_axlock_f = rd_req_desc_c_attr_reg[2];
   assign rd_req_desc_c_attr_axburst_f = rd_req_desc_c_attr_reg[1:0];
   assign rd_req_desc_c_axaddr_0_addr_f = rd_req_desc_c_axaddr_0_reg[31:0];
   assign rd_req_desc_c_axaddr_1_addr_f = rd_req_desc_c_axaddr_1_reg[31:0];
   assign rd_req_desc_c_axaddr_2_addr_f = rd_req_desc_c_axaddr_2_reg[31:0];
   assign rd_req_desc_c_axaddr_3_addr_f = rd_req_desc_c_axaddr_3_reg[31:0];
   assign rd_req_desc_c_axid_0_axid_f = rd_req_desc_c_axid_0_reg[31:0];
   assign rd_req_desc_c_axid_1_axid_f = rd_req_desc_c_axid_1_reg[31:0];
   assign rd_req_desc_c_axid_2_axid_f = rd_req_desc_c_axid_2_reg[31:0];
   assign rd_req_desc_c_axid_3_axid_f = rd_req_desc_c_axid_3_reg[31:0];
   assign rd_req_desc_c_axuser_0_axuser_f = rd_req_desc_c_axuser_0_reg[31:0];
   assign rd_req_desc_c_axuser_1_axuser_f = rd_req_desc_c_axuser_1_reg[31:0];
   assign rd_req_desc_c_axuser_2_axuser_f = rd_req_desc_c_axuser_2_reg[31:0];
   assign rd_req_desc_c_axuser_3_axuser_f = rd_req_desc_c_axuser_3_reg[31:0];
   assign rd_req_desc_c_axuser_4_axuser_f = rd_req_desc_c_axuser_4_reg[31:0];
   assign rd_req_desc_c_axuser_5_axuser_f = rd_req_desc_c_axuser_5_reg[31:0];
   assign rd_req_desc_c_axuser_6_axuser_f = rd_req_desc_c_axuser_6_reg[31:0];
   assign rd_req_desc_c_axuser_7_axuser_f = rd_req_desc_c_axuser_7_reg[31:0];
   assign rd_req_desc_c_axuser_8_axuser_f = rd_req_desc_c_axuser_8_reg[31:0];
   assign rd_req_desc_c_axuser_9_axuser_f = rd_req_desc_c_axuser_9_reg[31:0];
   assign rd_req_desc_c_axuser_10_axuser_f = rd_req_desc_c_axuser_10_reg[31:0];
   assign rd_req_desc_c_axuser_11_axuser_f = rd_req_desc_c_axuser_11_reg[31:0];
   assign rd_req_desc_c_axuser_12_axuser_f = rd_req_desc_c_axuser_12_reg[31:0];
   assign rd_req_desc_c_axuser_13_axuser_f = rd_req_desc_c_axuser_13_reg[31:0];
   assign rd_req_desc_c_axuser_14_axuser_f = rd_req_desc_c_axuser_14_reg[31:0];
   assign rd_req_desc_c_axuser_15_axuser_f = rd_req_desc_c_axuser_15_reg[31:0];
   assign rd_resp_desc_c_data_offset_addr_f = rd_resp_desc_c_data_offset_reg[13:0];
   assign rd_resp_desc_c_data_size_size_f = rd_resp_desc_c_data_size_reg[31:0];
   assign rd_resp_desc_c_data_host_addr_0_addr_f = rd_resp_desc_c_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_c_data_host_addr_1_addr_f = rd_resp_desc_c_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_c_data_host_addr_2_addr_f = rd_resp_desc_c_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_c_data_host_addr_3_addr_f = rd_resp_desc_c_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_c_resp_resp_f = rd_resp_desc_c_resp_reg[4:0];
   assign rd_resp_desc_c_xid_0_xid_f = rd_resp_desc_c_xid_0_reg[31:0];
   assign rd_resp_desc_c_xid_1_xid_f = rd_resp_desc_c_xid_1_reg[31:0];
   assign rd_resp_desc_c_xid_2_xid_f = rd_resp_desc_c_xid_2_reg[31:0];
   assign rd_resp_desc_c_xid_3_xid_f = rd_resp_desc_c_xid_3_reg[31:0];
   assign rd_resp_desc_c_xuser_0_xuser_f = rd_resp_desc_c_xuser_0_reg[31:0];
   assign rd_resp_desc_c_xuser_1_xuser_f = rd_resp_desc_c_xuser_1_reg[31:0];
   assign rd_resp_desc_c_xuser_2_xuser_f = rd_resp_desc_c_xuser_2_reg[31:0];
   assign rd_resp_desc_c_xuser_3_xuser_f = rd_resp_desc_c_xuser_3_reg[31:0];
   assign rd_resp_desc_c_xuser_4_xuser_f = rd_resp_desc_c_xuser_4_reg[31:0];
   assign rd_resp_desc_c_xuser_5_xuser_f = rd_resp_desc_c_xuser_5_reg[31:0];
   assign rd_resp_desc_c_xuser_6_xuser_f = rd_resp_desc_c_xuser_6_reg[31:0];
   assign rd_resp_desc_c_xuser_7_xuser_f = rd_resp_desc_c_xuser_7_reg[31:0];
   assign rd_resp_desc_c_xuser_8_xuser_f = rd_resp_desc_c_xuser_8_reg[31:0];
   assign rd_resp_desc_c_xuser_9_xuser_f = rd_resp_desc_c_xuser_9_reg[31:0];
   assign rd_resp_desc_c_xuser_10_xuser_f = rd_resp_desc_c_xuser_10_reg[31:0];
   assign rd_resp_desc_c_xuser_11_xuser_f = rd_resp_desc_c_xuser_11_reg[31:0];
   assign rd_resp_desc_c_xuser_12_xuser_f = rd_resp_desc_c_xuser_12_reg[31:0];
   assign rd_resp_desc_c_xuser_13_xuser_f = rd_resp_desc_c_xuser_13_reg[31:0];
   assign rd_resp_desc_c_xuser_14_xuser_f = rd_resp_desc_c_xuser_14_reg[31:0];
   assign rd_resp_desc_c_xuser_15_xuser_f = rd_resp_desc_c_xuser_15_reg[31:0];
   assign wr_req_desc_c_txn_type_wr_strb_f = wr_req_desc_c_txn_type_reg[1];
   assign wr_req_desc_c_size_txn_size_f = wr_req_desc_c_size_reg[31:0];
   assign wr_req_desc_c_data_offset_addr_f = wr_req_desc_c_data_offset_reg[13:0];
   assign wr_req_desc_c_data_host_addr_0_addr_f = wr_req_desc_c_data_host_addr_0_reg[31:0];
   assign wr_req_desc_c_data_host_addr_1_addr_f = wr_req_desc_c_data_host_addr_1_reg[31:0];
   assign wr_req_desc_c_data_host_addr_2_addr_f = wr_req_desc_c_data_host_addr_2_reg[31:0];
   assign wr_req_desc_c_data_host_addr_3_addr_f = wr_req_desc_c_data_host_addr_3_reg[31:0];
   assign wr_req_desc_c_wstrb_host_addr_0_addr_f = wr_req_desc_c_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_c_wstrb_host_addr_1_addr_f = wr_req_desc_c_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_c_wstrb_host_addr_2_addr_f = wr_req_desc_c_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_c_wstrb_host_addr_3_addr_f = wr_req_desc_c_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_c_axsize_axsize_f = wr_req_desc_c_axsize_reg[2:0];
   assign wr_req_desc_c_attr_axsnoop_f = wr_req_desc_c_attr_reg[27:24];
   assign wr_req_desc_c_attr_axdomain_f = wr_req_desc_c_attr_reg[23:22];
   assign wr_req_desc_c_attr_axbar_f = wr_req_desc_c_attr_reg[21:20];
   assign wr_req_desc_c_attr_awunique_f = wr_req_desc_c_attr_reg[19];
   assign wr_req_desc_c_attr_axregion_f = wr_req_desc_c_attr_reg[18:15];
   assign wr_req_desc_c_attr_axqos_f = wr_req_desc_c_attr_reg[14:11];
   assign wr_req_desc_c_attr_axprot_f = wr_req_desc_c_attr_reg[10:8];
   assign wr_req_desc_c_attr_axcache_f = wr_req_desc_c_attr_reg[7:4];
   assign wr_req_desc_c_attr_axlock_f = wr_req_desc_c_attr_reg[2];
   assign wr_req_desc_c_attr_axburst_f = wr_req_desc_c_attr_reg[1:0];
   assign wr_req_desc_c_axaddr_0_addr_f = wr_req_desc_c_axaddr_0_reg[31:0];
   assign wr_req_desc_c_axaddr_1_addr_f = wr_req_desc_c_axaddr_1_reg[31:0];
   assign wr_req_desc_c_axaddr_2_addr_f = wr_req_desc_c_axaddr_2_reg[31:0];
   assign wr_req_desc_c_axaddr_3_addr_f = wr_req_desc_c_axaddr_3_reg[31:0];
   assign wr_req_desc_c_axid_0_axid_f = wr_req_desc_c_axid_0_reg[31:0];
   assign wr_req_desc_c_axid_1_axid_f = wr_req_desc_c_axid_1_reg[31:0];
   assign wr_req_desc_c_axid_2_axid_f = wr_req_desc_c_axid_2_reg[31:0];
   assign wr_req_desc_c_axid_3_axid_f = wr_req_desc_c_axid_3_reg[31:0];
   assign wr_req_desc_c_axuser_0_axuser_f = wr_req_desc_c_axuser_0_reg[31:0];
   assign wr_req_desc_c_axuser_1_axuser_f = wr_req_desc_c_axuser_1_reg[31:0];
   assign wr_req_desc_c_axuser_2_axuser_f = wr_req_desc_c_axuser_2_reg[31:0];
   assign wr_req_desc_c_axuser_3_axuser_f = wr_req_desc_c_axuser_3_reg[31:0];
   assign wr_req_desc_c_axuser_4_axuser_f = wr_req_desc_c_axuser_4_reg[31:0];
   assign wr_req_desc_c_axuser_5_axuser_f = wr_req_desc_c_axuser_5_reg[31:0];
   assign wr_req_desc_c_axuser_6_axuser_f = wr_req_desc_c_axuser_6_reg[31:0];
   assign wr_req_desc_c_axuser_7_axuser_f = wr_req_desc_c_axuser_7_reg[31:0];
   assign wr_req_desc_c_axuser_8_axuser_f = wr_req_desc_c_axuser_8_reg[31:0];
   assign wr_req_desc_c_axuser_9_axuser_f = wr_req_desc_c_axuser_9_reg[31:0];
   assign wr_req_desc_c_axuser_10_axuser_f = wr_req_desc_c_axuser_10_reg[31:0];
   assign wr_req_desc_c_axuser_11_axuser_f = wr_req_desc_c_axuser_11_reg[31:0];
   assign wr_req_desc_c_axuser_12_axuser_f = wr_req_desc_c_axuser_12_reg[31:0];
   assign wr_req_desc_c_axuser_13_axuser_f = wr_req_desc_c_axuser_13_reg[31:0];
   assign wr_req_desc_c_axuser_14_axuser_f = wr_req_desc_c_axuser_14_reg[31:0];
   assign wr_req_desc_c_axuser_15_axuser_f = wr_req_desc_c_axuser_15_reg[31:0];
   assign wr_req_desc_c_wuser_0_wuser_f = wr_req_desc_c_wuser_0_reg[31:0];
   assign wr_req_desc_c_wuser_1_wuser_f = wr_req_desc_c_wuser_1_reg[31:0];
   assign wr_req_desc_c_wuser_2_wuser_f = wr_req_desc_c_wuser_2_reg[31:0];
   assign wr_req_desc_c_wuser_3_wuser_f = wr_req_desc_c_wuser_3_reg[31:0];
   assign wr_req_desc_c_wuser_4_wuser_f = wr_req_desc_c_wuser_4_reg[31:0];
   assign wr_req_desc_c_wuser_5_wuser_f = wr_req_desc_c_wuser_5_reg[31:0];
   assign wr_req_desc_c_wuser_6_wuser_f = wr_req_desc_c_wuser_6_reg[31:0];
   assign wr_req_desc_c_wuser_7_wuser_f = wr_req_desc_c_wuser_7_reg[31:0];
   assign wr_req_desc_c_wuser_8_wuser_f = wr_req_desc_c_wuser_8_reg[31:0];
   assign wr_req_desc_c_wuser_9_wuser_f = wr_req_desc_c_wuser_9_reg[31:0];
   assign wr_req_desc_c_wuser_10_wuser_f = wr_req_desc_c_wuser_10_reg[31:0];
   assign wr_req_desc_c_wuser_11_wuser_f = wr_req_desc_c_wuser_11_reg[31:0];
   assign wr_req_desc_c_wuser_12_wuser_f = wr_req_desc_c_wuser_12_reg[31:0];
   assign wr_req_desc_c_wuser_13_wuser_f = wr_req_desc_c_wuser_13_reg[31:0];
   assign wr_req_desc_c_wuser_14_wuser_f = wr_req_desc_c_wuser_14_reg[31:0];
   assign wr_req_desc_c_wuser_15_wuser_f = wr_req_desc_c_wuser_15_reg[31:0];
   assign wr_resp_desc_c_resp_resp_f = wr_resp_desc_c_resp_reg[4:0];
   assign wr_resp_desc_c_xid_0_xid_f = wr_resp_desc_c_xid_0_reg[31:0];
   assign wr_resp_desc_c_xid_1_xid_f = wr_resp_desc_c_xid_1_reg[31:0];
   assign wr_resp_desc_c_xid_2_xid_f = wr_resp_desc_c_xid_2_reg[31:0];
   assign wr_resp_desc_c_xid_3_xid_f = wr_resp_desc_c_xid_3_reg[31:0];
   assign wr_resp_desc_c_xuser_0_xuser_f = wr_resp_desc_c_xuser_0_reg[31:0];
   assign wr_resp_desc_c_xuser_1_xuser_f = wr_resp_desc_c_xuser_1_reg[31:0];
   assign wr_resp_desc_c_xuser_2_xuser_f = wr_resp_desc_c_xuser_2_reg[31:0];
   assign wr_resp_desc_c_xuser_3_xuser_f = wr_resp_desc_c_xuser_3_reg[31:0];
   assign wr_resp_desc_c_xuser_4_xuser_f = wr_resp_desc_c_xuser_4_reg[31:0];
   assign wr_resp_desc_c_xuser_5_xuser_f = wr_resp_desc_c_xuser_5_reg[31:0];
   assign wr_resp_desc_c_xuser_6_xuser_f = wr_resp_desc_c_xuser_6_reg[31:0];
   assign wr_resp_desc_c_xuser_7_xuser_f = wr_resp_desc_c_xuser_7_reg[31:0];
   assign wr_resp_desc_c_xuser_8_xuser_f = wr_resp_desc_c_xuser_8_reg[31:0];
   assign wr_resp_desc_c_xuser_9_xuser_f = wr_resp_desc_c_xuser_9_reg[31:0];
   assign wr_resp_desc_c_xuser_10_xuser_f = wr_resp_desc_c_xuser_10_reg[31:0];
   assign wr_resp_desc_c_xuser_11_xuser_f = wr_resp_desc_c_xuser_11_reg[31:0];
   assign wr_resp_desc_c_xuser_12_xuser_f = wr_resp_desc_c_xuser_12_reg[31:0];
   assign wr_resp_desc_c_xuser_13_xuser_f = wr_resp_desc_c_xuser_13_reg[31:0];
   assign wr_resp_desc_c_xuser_14_xuser_f = wr_resp_desc_c_xuser_14_reg[31:0];
   assign wr_resp_desc_c_xuser_15_xuser_f = wr_resp_desc_c_xuser_15_reg[31:0];
   assign sn_req_desc_c_attr_acsnoop_f = sn_req_desc_c_attr_reg[27:24];
   assign sn_req_desc_c_attr_acprot_f = sn_req_desc_c_attr_reg[10:8];
   assign sn_req_desc_c_acaddr_0_addr_f = sn_req_desc_c_acaddr_0_reg[31:0];
   assign sn_req_desc_c_acaddr_1_addr_f = sn_req_desc_c_acaddr_1_reg[31:0];
   assign sn_req_desc_c_acaddr_2_addr_f = sn_req_desc_c_acaddr_2_reg[31:0];
   assign sn_req_desc_c_acaddr_3_addr_f = sn_req_desc_c_acaddr_3_reg[31:0];
   assign sn_resp_desc_c_resp_resp_f = sn_resp_desc_c_resp_reg[4:0];
   assign rd_req_desc_d_size_txn_size_f = rd_req_desc_d_size_reg[31:0];
   assign rd_req_desc_d_axsize_axsize_f = rd_req_desc_d_axsize_reg[2:0];
   assign rd_req_desc_d_attr_axsnoop_f = rd_req_desc_d_attr_reg[27:24];
   assign rd_req_desc_d_attr_axdomain_f = rd_req_desc_d_attr_reg[23:22];
   assign rd_req_desc_d_attr_axbar_f = rd_req_desc_d_attr_reg[21:20];
   assign rd_req_desc_d_attr_axregion_f = rd_req_desc_d_attr_reg[18:15];
   assign rd_req_desc_d_attr_axqos_f = rd_req_desc_d_attr_reg[14:11];
   assign rd_req_desc_d_attr_axprot_f = rd_req_desc_d_attr_reg[10:8];
   assign rd_req_desc_d_attr_axcache_f = rd_req_desc_d_attr_reg[7:4];
   assign rd_req_desc_d_attr_axlock_f = rd_req_desc_d_attr_reg[2];
   assign rd_req_desc_d_attr_axburst_f = rd_req_desc_d_attr_reg[1:0];
   assign rd_req_desc_d_axaddr_0_addr_f = rd_req_desc_d_axaddr_0_reg[31:0];
   assign rd_req_desc_d_axaddr_1_addr_f = rd_req_desc_d_axaddr_1_reg[31:0];
   assign rd_req_desc_d_axaddr_2_addr_f = rd_req_desc_d_axaddr_2_reg[31:0];
   assign rd_req_desc_d_axaddr_3_addr_f = rd_req_desc_d_axaddr_3_reg[31:0];
   assign rd_req_desc_d_axid_0_axid_f = rd_req_desc_d_axid_0_reg[31:0];
   assign rd_req_desc_d_axid_1_axid_f = rd_req_desc_d_axid_1_reg[31:0];
   assign rd_req_desc_d_axid_2_axid_f = rd_req_desc_d_axid_2_reg[31:0];
   assign rd_req_desc_d_axid_3_axid_f = rd_req_desc_d_axid_3_reg[31:0];
   assign rd_req_desc_d_axuser_0_axuser_f = rd_req_desc_d_axuser_0_reg[31:0];
   assign rd_req_desc_d_axuser_1_axuser_f = rd_req_desc_d_axuser_1_reg[31:0];
   assign rd_req_desc_d_axuser_2_axuser_f = rd_req_desc_d_axuser_2_reg[31:0];
   assign rd_req_desc_d_axuser_3_axuser_f = rd_req_desc_d_axuser_3_reg[31:0];
   assign rd_req_desc_d_axuser_4_axuser_f = rd_req_desc_d_axuser_4_reg[31:0];
   assign rd_req_desc_d_axuser_5_axuser_f = rd_req_desc_d_axuser_5_reg[31:0];
   assign rd_req_desc_d_axuser_6_axuser_f = rd_req_desc_d_axuser_6_reg[31:0];
   assign rd_req_desc_d_axuser_7_axuser_f = rd_req_desc_d_axuser_7_reg[31:0];
   assign rd_req_desc_d_axuser_8_axuser_f = rd_req_desc_d_axuser_8_reg[31:0];
   assign rd_req_desc_d_axuser_9_axuser_f = rd_req_desc_d_axuser_9_reg[31:0];
   assign rd_req_desc_d_axuser_10_axuser_f = rd_req_desc_d_axuser_10_reg[31:0];
   assign rd_req_desc_d_axuser_11_axuser_f = rd_req_desc_d_axuser_11_reg[31:0];
   assign rd_req_desc_d_axuser_12_axuser_f = rd_req_desc_d_axuser_12_reg[31:0];
   assign rd_req_desc_d_axuser_13_axuser_f = rd_req_desc_d_axuser_13_reg[31:0];
   assign rd_req_desc_d_axuser_14_axuser_f = rd_req_desc_d_axuser_14_reg[31:0];
   assign rd_req_desc_d_axuser_15_axuser_f = rd_req_desc_d_axuser_15_reg[31:0];
   assign rd_resp_desc_d_data_offset_addr_f = rd_resp_desc_d_data_offset_reg[13:0];
   assign rd_resp_desc_d_data_size_size_f = rd_resp_desc_d_data_size_reg[31:0];
   assign rd_resp_desc_d_data_host_addr_0_addr_f = rd_resp_desc_d_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_d_data_host_addr_1_addr_f = rd_resp_desc_d_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_d_data_host_addr_2_addr_f = rd_resp_desc_d_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_d_data_host_addr_3_addr_f = rd_resp_desc_d_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_d_resp_resp_f = rd_resp_desc_d_resp_reg[4:0];
   assign rd_resp_desc_d_xid_0_xid_f = rd_resp_desc_d_xid_0_reg[31:0];
   assign rd_resp_desc_d_xid_1_xid_f = rd_resp_desc_d_xid_1_reg[31:0];
   assign rd_resp_desc_d_xid_2_xid_f = rd_resp_desc_d_xid_2_reg[31:0];
   assign rd_resp_desc_d_xid_3_xid_f = rd_resp_desc_d_xid_3_reg[31:0];
   assign rd_resp_desc_d_xuser_0_xuser_f = rd_resp_desc_d_xuser_0_reg[31:0];
   assign rd_resp_desc_d_xuser_1_xuser_f = rd_resp_desc_d_xuser_1_reg[31:0];
   assign rd_resp_desc_d_xuser_2_xuser_f = rd_resp_desc_d_xuser_2_reg[31:0];
   assign rd_resp_desc_d_xuser_3_xuser_f = rd_resp_desc_d_xuser_3_reg[31:0];
   assign rd_resp_desc_d_xuser_4_xuser_f = rd_resp_desc_d_xuser_4_reg[31:0];
   assign rd_resp_desc_d_xuser_5_xuser_f = rd_resp_desc_d_xuser_5_reg[31:0];
   assign rd_resp_desc_d_xuser_6_xuser_f = rd_resp_desc_d_xuser_6_reg[31:0];
   assign rd_resp_desc_d_xuser_7_xuser_f = rd_resp_desc_d_xuser_7_reg[31:0];
   assign rd_resp_desc_d_xuser_8_xuser_f = rd_resp_desc_d_xuser_8_reg[31:0];
   assign rd_resp_desc_d_xuser_9_xuser_f = rd_resp_desc_d_xuser_9_reg[31:0];
   assign rd_resp_desc_d_xuser_10_xuser_f = rd_resp_desc_d_xuser_10_reg[31:0];
   assign rd_resp_desc_d_xuser_11_xuser_f = rd_resp_desc_d_xuser_11_reg[31:0];
   assign rd_resp_desc_d_xuser_12_xuser_f = rd_resp_desc_d_xuser_12_reg[31:0];
   assign rd_resp_desc_d_xuser_13_xuser_f = rd_resp_desc_d_xuser_13_reg[31:0];
   assign rd_resp_desc_d_xuser_14_xuser_f = rd_resp_desc_d_xuser_14_reg[31:0];
   assign rd_resp_desc_d_xuser_15_xuser_f = rd_resp_desc_d_xuser_15_reg[31:0];
   assign wr_req_desc_d_txn_type_wr_strb_f = wr_req_desc_d_txn_type_reg[1];
   assign wr_req_desc_d_size_txn_size_f = wr_req_desc_d_size_reg[31:0];
   assign wr_req_desc_d_data_offset_addr_f = wr_req_desc_d_data_offset_reg[13:0];
   assign wr_req_desc_d_data_host_addr_0_addr_f = wr_req_desc_d_data_host_addr_0_reg[31:0];
   assign wr_req_desc_d_data_host_addr_1_addr_f = wr_req_desc_d_data_host_addr_1_reg[31:0];
   assign wr_req_desc_d_data_host_addr_2_addr_f = wr_req_desc_d_data_host_addr_2_reg[31:0];
   assign wr_req_desc_d_data_host_addr_3_addr_f = wr_req_desc_d_data_host_addr_3_reg[31:0];
   assign wr_req_desc_d_wstrb_host_addr_0_addr_f = wr_req_desc_d_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_d_wstrb_host_addr_1_addr_f = wr_req_desc_d_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_d_wstrb_host_addr_2_addr_f = wr_req_desc_d_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_d_wstrb_host_addr_3_addr_f = wr_req_desc_d_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_d_axsize_axsize_f = wr_req_desc_d_axsize_reg[2:0];
   assign wr_req_desc_d_attr_axsnoop_f = wr_req_desc_d_attr_reg[27:24];
   assign wr_req_desc_d_attr_axdomain_f = wr_req_desc_d_attr_reg[23:22];
   assign wr_req_desc_d_attr_axbar_f = wr_req_desc_d_attr_reg[21:20];
   assign wr_req_desc_d_attr_awunique_f = wr_req_desc_d_attr_reg[19];
   assign wr_req_desc_d_attr_axregion_f = wr_req_desc_d_attr_reg[18:15];
   assign wr_req_desc_d_attr_axqos_f = wr_req_desc_d_attr_reg[14:11];
   assign wr_req_desc_d_attr_axprot_f = wr_req_desc_d_attr_reg[10:8];
   assign wr_req_desc_d_attr_axcache_f = wr_req_desc_d_attr_reg[7:4];
   assign wr_req_desc_d_attr_axlock_f = wr_req_desc_d_attr_reg[2];
   assign wr_req_desc_d_attr_axburst_f = wr_req_desc_d_attr_reg[1:0];
   assign wr_req_desc_d_axaddr_0_addr_f = wr_req_desc_d_axaddr_0_reg[31:0];
   assign wr_req_desc_d_axaddr_1_addr_f = wr_req_desc_d_axaddr_1_reg[31:0];
   assign wr_req_desc_d_axaddr_2_addr_f = wr_req_desc_d_axaddr_2_reg[31:0];
   assign wr_req_desc_d_axaddr_3_addr_f = wr_req_desc_d_axaddr_3_reg[31:0];
   assign wr_req_desc_d_axid_0_axid_f = wr_req_desc_d_axid_0_reg[31:0];
   assign wr_req_desc_d_axid_1_axid_f = wr_req_desc_d_axid_1_reg[31:0];
   assign wr_req_desc_d_axid_2_axid_f = wr_req_desc_d_axid_2_reg[31:0];
   assign wr_req_desc_d_axid_3_axid_f = wr_req_desc_d_axid_3_reg[31:0];
   assign wr_req_desc_d_axuser_0_axuser_f = wr_req_desc_d_axuser_0_reg[31:0];
   assign wr_req_desc_d_axuser_1_axuser_f = wr_req_desc_d_axuser_1_reg[31:0];
   assign wr_req_desc_d_axuser_2_axuser_f = wr_req_desc_d_axuser_2_reg[31:0];
   assign wr_req_desc_d_axuser_3_axuser_f = wr_req_desc_d_axuser_3_reg[31:0];
   assign wr_req_desc_d_axuser_4_axuser_f = wr_req_desc_d_axuser_4_reg[31:0];
   assign wr_req_desc_d_axuser_5_axuser_f = wr_req_desc_d_axuser_5_reg[31:0];
   assign wr_req_desc_d_axuser_6_axuser_f = wr_req_desc_d_axuser_6_reg[31:0];
   assign wr_req_desc_d_axuser_7_axuser_f = wr_req_desc_d_axuser_7_reg[31:0];
   assign wr_req_desc_d_axuser_8_axuser_f = wr_req_desc_d_axuser_8_reg[31:0];
   assign wr_req_desc_d_axuser_9_axuser_f = wr_req_desc_d_axuser_9_reg[31:0];
   assign wr_req_desc_d_axuser_10_axuser_f = wr_req_desc_d_axuser_10_reg[31:0];
   assign wr_req_desc_d_axuser_11_axuser_f = wr_req_desc_d_axuser_11_reg[31:0];
   assign wr_req_desc_d_axuser_12_axuser_f = wr_req_desc_d_axuser_12_reg[31:0];
   assign wr_req_desc_d_axuser_13_axuser_f = wr_req_desc_d_axuser_13_reg[31:0];
   assign wr_req_desc_d_axuser_14_axuser_f = wr_req_desc_d_axuser_14_reg[31:0];
   assign wr_req_desc_d_axuser_15_axuser_f = wr_req_desc_d_axuser_15_reg[31:0];
   assign wr_req_desc_d_wuser_0_wuser_f = wr_req_desc_d_wuser_0_reg[31:0];
   assign wr_req_desc_d_wuser_1_wuser_f = wr_req_desc_d_wuser_1_reg[31:0];
   assign wr_req_desc_d_wuser_2_wuser_f = wr_req_desc_d_wuser_2_reg[31:0];
   assign wr_req_desc_d_wuser_3_wuser_f = wr_req_desc_d_wuser_3_reg[31:0];
   assign wr_req_desc_d_wuser_4_wuser_f = wr_req_desc_d_wuser_4_reg[31:0];
   assign wr_req_desc_d_wuser_5_wuser_f = wr_req_desc_d_wuser_5_reg[31:0];
   assign wr_req_desc_d_wuser_6_wuser_f = wr_req_desc_d_wuser_6_reg[31:0];
   assign wr_req_desc_d_wuser_7_wuser_f = wr_req_desc_d_wuser_7_reg[31:0];
   assign wr_req_desc_d_wuser_8_wuser_f = wr_req_desc_d_wuser_8_reg[31:0];
   assign wr_req_desc_d_wuser_9_wuser_f = wr_req_desc_d_wuser_9_reg[31:0];
   assign wr_req_desc_d_wuser_10_wuser_f = wr_req_desc_d_wuser_10_reg[31:0];
   assign wr_req_desc_d_wuser_11_wuser_f = wr_req_desc_d_wuser_11_reg[31:0];
   assign wr_req_desc_d_wuser_12_wuser_f = wr_req_desc_d_wuser_12_reg[31:0];
   assign wr_req_desc_d_wuser_13_wuser_f = wr_req_desc_d_wuser_13_reg[31:0];
   assign wr_req_desc_d_wuser_14_wuser_f = wr_req_desc_d_wuser_14_reg[31:0];
   assign wr_req_desc_d_wuser_15_wuser_f = wr_req_desc_d_wuser_15_reg[31:0];
   assign wr_resp_desc_d_resp_resp_f = wr_resp_desc_d_resp_reg[4:0];
   assign wr_resp_desc_d_xid_0_xid_f = wr_resp_desc_d_xid_0_reg[31:0];
   assign wr_resp_desc_d_xid_1_xid_f = wr_resp_desc_d_xid_1_reg[31:0];
   assign wr_resp_desc_d_xid_2_xid_f = wr_resp_desc_d_xid_2_reg[31:0];
   assign wr_resp_desc_d_xid_3_xid_f = wr_resp_desc_d_xid_3_reg[31:0];
   assign wr_resp_desc_d_xuser_0_xuser_f = wr_resp_desc_d_xuser_0_reg[31:0];
   assign wr_resp_desc_d_xuser_1_xuser_f = wr_resp_desc_d_xuser_1_reg[31:0];
   assign wr_resp_desc_d_xuser_2_xuser_f = wr_resp_desc_d_xuser_2_reg[31:0];
   assign wr_resp_desc_d_xuser_3_xuser_f = wr_resp_desc_d_xuser_3_reg[31:0];
   assign wr_resp_desc_d_xuser_4_xuser_f = wr_resp_desc_d_xuser_4_reg[31:0];
   assign wr_resp_desc_d_xuser_5_xuser_f = wr_resp_desc_d_xuser_5_reg[31:0];
   assign wr_resp_desc_d_xuser_6_xuser_f = wr_resp_desc_d_xuser_6_reg[31:0];
   assign wr_resp_desc_d_xuser_7_xuser_f = wr_resp_desc_d_xuser_7_reg[31:0];
   assign wr_resp_desc_d_xuser_8_xuser_f = wr_resp_desc_d_xuser_8_reg[31:0];
   assign wr_resp_desc_d_xuser_9_xuser_f = wr_resp_desc_d_xuser_9_reg[31:0];
   assign wr_resp_desc_d_xuser_10_xuser_f = wr_resp_desc_d_xuser_10_reg[31:0];
   assign wr_resp_desc_d_xuser_11_xuser_f = wr_resp_desc_d_xuser_11_reg[31:0];
   assign wr_resp_desc_d_xuser_12_xuser_f = wr_resp_desc_d_xuser_12_reg[31:0];
   assign wr_resp_desc_d_xuser_13_xuser_f = wr_resp_desc_d_xuser_13_reg[31:0];
   assign wr_resp_desc_d_xuser_14_xuser_f = wr_resp_desc_d_xuser_14_reg[31:0];
   assign wr_resp_desc_d_xuser_15_xuser_f = wr_resp_desc_d_xuser_15_reg[31:0];
   assign sn_req_desc_d_attr_acsnoop_f = sn_req_desc_d_attr_reg[27:24];
   assign sn_req_desc_d_attr_acprot_f = sn_req_desc_d_attr_reg[10:8];
   assign sn_req_desc_d_acaddr_0_addr_f = sn_req_desc_d_acaddr_0_reg[31:0];
   assign sn_req_desc_d_acaddr_1_addr_f = sn_req_desc_d_acaddr_1_reg[31:0];
   assign sn_req_desc_d_acaddr_2_addr_f = sn_req_desc_d_acaddr_2_reg[31:0];
   assign sn_req_desc_d_acaddr_3_addr_f = sn_req_desc_d_acaddr_3_reg[31:0];
   assign sn_resp_desc_d_resp_resp_f = sn_resp_desc_d_resp_reg[4:0];
   assign rd_req_desc_e_size_txn_size_f = rd_req_desc_e_size_reg[31:0];
   assign rd_req_desc_e_axsize_axsize_f = rd_req_desc_e_axsize_reg[2:0];
   assign rd_req_desc_e_attr_axsnoop_f = rd_req_desc_e_attr_reg[27:24];
   assign rd_req_desc_e_attr_axdomain_f = rd_req_desc_e_attr_reg[23:22];
   assign rd_req_desc_e_attr_axbar_f = rd_req_desc_e_attr_reg[21:20];
   assign rd_req_desc_e_attr_axregion_f = rd_req_desc_e_attr_reg[18:15];
   assign rd_req_desc_e_attr_axqos_f = rd_req_desc_e_attr_reg[14:11];
   assign rd_req_desc_e_attr_axprot_f = rd_req_desc_e_attr_reg[10:8];
   assign rd_req_desc_e_attr_axcache_f = rd_req_desc_e_attr_reg[7:4];
   assign rd_req_desc_e_attr_axlock_f = rd_req_desc_e_attr_reg[2];
   assign rd_req_desc_e_attr_axburst_f = rd_req_desc_e_attr_reg[1:0];
   assign rd_req_desc_e_axaddr_0_addr_f = rd_req_desc_e_axaddr_0_reg[31:0];
   assign rd_req_desc_e_axaddr_1_addr_f = rd_req_desc_e_axaddr_1_reg[31:0];
   assign rd_req_desc_e_axaddr_2_addr_f = rd_req_desc_e_axaddr_2_reg[31:0];
   assign rd_req_desc_e_axaddr_3_addr_f = rd_req_desc_e_axaddr_3_reg[31:0];
   assign rd_req_desc_e_axid_0_axid_f = rd_req_desc_e_axid_0_reg[31:0];
   assign rd_req_desc_e_axid_1_axid_f = rd_req_desc_e_axid_1_reg[31:0];
   assign rd_req_desc_e_axid_2_axid_f = rd_req_desc_e_axid_2_reg[31:0];
   assign rd_req_desc_e_axid_3_axid_f = rd_req_desc_e_axid_3_reg[31:0];
   assign rd_req_desc_e_axuser_0_axuser_f = rd_req_desc_e_axuser_0_reg[31:0];
   assign rd_req_desc_e_axuser_1_axuser_f = rd_req_desc_e_axuser_1_reg[31:0];
   assign rd_req_desc_e_axuser_2_axuser_f = rd_req_desc_e_axuser_2_reg[31:0];
   assign rd_req_desc_e_axuser_3_axuser_f = rd_req_desc_e_axuser_3_reg[31:0];
   assign rd_req_desc_e_axuser_4_axuser_f = rd_req_desc_e_axuser_4_reg[31:0];
   assign rd_req_desc_e_axuser_5_axuser_f = rd_req_desc_e_axuser_5_reg[31:0];
   assign rd_req_desc_e_axuser_6_axuser_f = rd_req_desc_e_axuser_6_reg[31:0];
   assign rd_req_desc_e_axuser_7_axuser_f = rd_req_desc_e_axuser_7_reg[31:0];
   assign rd_req_desc_e_axuser_8_axuser_f = rd_req_desc_e_axuser_8_reg[31:0];
   assign rd_req_desc_e_axuser_9_axuser_f = rd_req_desc_e_axuser_9_reg[31:0];
   assign rd_req_desc_e_axuser_10_axuser_f = rd_req_desc_e_axuser_10_reg[31:0];
   assign rd_req_desc_e_axuser_11_axuser_f = rd_req_desc_e_axuser_11_reg[31:0];
   assign rd_req_desc_e_axuser_12_axuser_f = rd_req_desc_e_axuser_12_reg[31:0];
   assign rd_req_desc_e_axuser_13_axuser_f = rd_req_desc_e_axuser_13_reg[31:0];
   assign rd_req_desc_e_axuser_14_axuser_f = rd_req_desc_e_axuser_14_reg[31:0];
   assign rd_req_desc_e_axuser_15_axuser_f = rd_req_desc_e_axuser_15_reg[31:0];
   assign rd_resp_desc_e_data_offset_addr_f = rd_resp_desc_e_data_offset_reg[13:0];
   assign rd_resp_desc_e_data_size_size_f = rd_resp_desc_e_data_size_reg[31:0];
   assign rd_resp_desc_e_data_host_addr_0_addr_f = rd_resp_desc_e_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_e_data_host_addr_1_addr_f = rd_resp_desc_e_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_e_data_host_addr_2_addr_f = rd_resp_desc_e_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_e_data_host_addr_3_addr_f = rd_resp_desc_e_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_e_resp_resp_f = rd_resp_desc_e_resp_reg[4:0];
   assign rd_resp_desc_e_xid_0_xid_f = rd_resp_desc_e_xid_0_reg[31:0];
   assign rd_resp_desc_e_xid_1_xid_f = rd_resp_desc_e_xid_1_reg[31:0];
   assign rd_resp_desc_e_xid_2_xid_f = rd_resp_desc_e_xid_2_reg[31:0];
   assign rd_resp_desc_e_xid_3_xid_f = rd_resp_desc_e_xid_3_reg[31:0];
   assign rd_resp_desc_e_xuser_0_xuser_f = rd_resp_desc_e_xuser_0_reg[31:0];
   assign rd_resp_desc_e_xuser_1_xuser_f = rd_resp_desc_e_xuser_1_reg[31:0];
   assign rd_resp_desc_e_xuser_2_xuser_f = rd_resp_desc_e_xuser_2_reg[31:0];
   assign rd_resp_desc_e_xuser_3_xuser_f = rd_resp_desc_e_xuser_3_reg[31:0];
   assign rd_resp_desc_e_xuser_4_xuser_f = rd_resp_desc_e_xuser_4_reg[31:0];
   assign rd_resp_desc_e_xuser_5_xuser_f = rd_resp_desc_e_xuser_5_reg[31:0];
   assign rd_resp_desc_e_xuser_6_xuser_f = rd_resp_desc_e_xuser_6_reg[31:0];
   assign rd_resp_desc_e_xuser_7_xuser_f = rd_resp_desc_e_xuser_7_reg[31:0];
   assign rd_resp_desc_e_xuser_8_xuser_f = rd_resp_desc_e_xuser_8_reg[31:0];
   assign rd_resp_desc_e_xuser_9_xuser_f = rd_resp_desc_e_xuser_9_reg[31:0];
   assign rd_resp_desc_e_xuser_10_xuser_f = rd_resp_desc_e_xuser_10_reg[31:0];
   assign rd_resp_desc_e_xuser_11_xuser_f = rd_resp_desc_e_xuser_11_reg[31:0];
   assign rd_resp_desc_e_xuser_12_xuser_f = rd_resp_desc_e_xuser_12_reg[31:0];
   assign rd_resp_desc_e_xuser_13_xuser_f = rd_resp_desc_e_xuser_13_reg[31:0];
   assign rd_resp_desc_e_xuser_14_xuser_f = rd_resp_desc_e_xuser_14_reg[31:0];
   assign rd_resp_desc_e_xuser_15_xuser_f = rd_resp_desc_e_xuser_15_reg[31:0];
   assign wr_req_desc_e_txn_type_wr_strb_f = wr_req_desc_e_txn_type_reg[1];
   assign wr_req_desc_e_size_txn_size_f = wr_req_desc_e_size_reg[31:0];
   assign wr_req_desc_e_data_offset_addr_f = wr_req_desc_e_data_offset_reg[13:0];
   assign wr_req_desc_e_data_host_addr_0_addr_f = wr_req_desc_e_data_host_addr_0_reg[31:0];
   assign wr_req_desc_e_data_host_addr_1_addr_f = wr_req_desc_e_data_host_addr_1_reg[31:0];
   assign wr_req_desc_e_data_host_addr_2_addr_f = wr_req_desc_e_data_host_addr_2_reg[31:0];
   assign wr_req_desc_e_data_host_addr_3_addr_f = wr_req_desc_e_data_host_addr_3_reg[31:0];
   assign wr_req_desc_e_wstrb_host_addr_0_addr_f = wr_req_desc_e_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_e_wstrb_host_addr_1_addr_f = wr_req_desc_e_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_e_wstrb_host_addr_2_addr_f = wr_req_desc_e_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_e_wstrb_host_addr_3_addr_f = wr_req_desc_e_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_e_axsize_axsize_f = wr_req_desc_e_axsize_reg[2:0];
   assign wr_req_desc_e_attr_axsnoop_f = wr_req_desc_e_attr_reg[27:24];
   assign wr_req_desc_e_attr_axdomain_f = wr_req_desc_e_attr_reg[23:22];
   assign wr_req_desc_e_attr_axbar_f = wr_req_desc_e_attr_reg[21:20];
   assign wr_req_desc_e_attr_awunique_f = wr_req_desc_e_attr_reg[19];
   assign wr_req_desc_e_attr_axregion_f = wr_req_desc_e_attr_reg[18:15];
   assign wr_req_desc_e_attr_axqos_f = wr_req_desc_e_attr_reg[14:11];
   assign wr_req_desc_e_attr_axprot_f = wr_req_desc_e_attr_reg[10:8];
   assign wr_req_desc_e_attr_axcache_f = wr_req_desc_e_attr_reg[7:4];
   assign wr_req_desc_e_attr_axlock_f = wr_req_desc_e_attr_reg[2];
   assign wr_req_desc_e_attr_axburst_f = wr_req_desc_e_attr_reg[1:0];
   assign wr_req_desc_e_axaddr_0_addr_f = wr_req_desc_e_axaddr_0_reg[31:0];
   assign wr_req_desc_e_axaddr_1_addr_f = wr_req_desc_e_axaddr_1_reg[31:0];
   assign wr_req_desc_e_axaddr_2_addr_f = wr_req_desc_e_axaddr_2_reg[31:0];
   assign wr_req_desc_e_axaddr_3_addr_f = wr_req_desc_e_axaddr_3_reg[31:0];
   assign wr_req_desc_e_axid_0_axid_f = wr_req_desc_e_axid_0_reg[31:0];
   assign wr_req_desc_e_axid_1_axid_f = wr_req_desc_e_axid_1_reg[31:0];
   assign wr_req_desc_e_axid_2_axid_f = wr_req_desc_e_axid_2_reg[31:0];
   assign wr_req_desc_e_axid_3_axid_f = wr_req_desc_e_axid_3_reg[31:0];
   assign wr_req_desc_e_axuser_0_axuser_f = wr_req_desc_e_axuser_0_reg[31:0];
   assign wr_req_desc_e_axuser_1_axuser_f = wr_req_desc_e_axuser_1_reg[31:0];
   assign wr_req_desc_e_axuser_2_axuser_f = wr_req_desc_e_axuser_2_reg[31:0];
   assign wr_req_desc_e_axuser_3_axuser_f = wr_req_desc_e_axuser_3_reg[31:0];
   assign wr_req_desc_e_axuser_4_axuser_f = wr_req_desc_e_axuser_4_reg[31:0];
   assign wr_req_desc_e_axuser_5_axuser_f = wr_req_desc_e_axuser_5_reg[31:0];
   assign wr_req_desc_e_axuser_6_axuser_f = wr_req_desc_e_axuser_6_reg[31:0];
   assign wr_req_desc_e_axuser_7_axuser_f = wr_req_desc_e_axuser_7_reg[31:0];
   assign wr_req_desc_e_axuser_8_axuser_f = wr_req_desc_e_axuser_8_reg[31:0];
   assign wr_req_desc_e_axuser_9_axuser_f = wr_req_desc_e_axuser_9_reg[31:0];
   assign wr_req_desc_e_axuser_10_axuser_f = wr_req_desc_e_axuser_10_reg[31:0];
   assign wr_req_desc_e_axuser_11_axuser_f = wr_req_desc_e_axuser_11_reg[31:0];
   assign wr_req_desc_e_axuser_12_axuser_f = wr_req_desc_e_axuser_12_reg[31:0];
   assign wr_req_desc_e_axuser_13_axuser_f = wr_req_desc_e_axuser_13_reg[31:0];
   assign wr_req_desc_e_axuser_14_axuser_f = wr_req_desc_e_axuser_14_reg[31:0];
   assign wr_req_desc_e_axuser_15_axuser_f = wr_req_desc_e_axuser_15_reg[31:0];
   assign wr_req_desc_e_wuser_0_wuser_f = wr_req_desc_e_wuser_0_reg[31:0];
   assign wr_req_desc_e_wuser_1_wuser_f = wr_req_desc_e_wuser_1_reg[31:0];
   assign wr_req_desc_e_wuser_2_wuser_f = wr_req_desc_e_wuser_2_reg[31:0];
   assign wr_req_desc_e_wuser_3_wuser_f = wr_req_desc_e_wuser_3_reg[31:0];
   assign wr_req_desc_e_wuser_4_wuser_f = wr_req_desc_e_wuser_4_reg[31:0];
   assign wr_req_desc_e_wuser_5_wuser_f = wr_req_desc_e_wuser_5_reg[31:0];
   assign wr_req_desc_e_wuser_6_wuser_f = wr_req_desc_e_wuser_6_reg[31:0];
   assign wr_req_desc_e_wuser_7_wuser_f = wr_req_desc_e_wuser_7_reg[31:0];
   assign wr_req_desc_e_wuser_8_wuser_f = wr_req_desc_e_wuser_8_reg[31:0];
   assign wr_req_desc_e_wuser_9_wuser_f = wr_req_desc_e_wuser_9_reg[31:0];
   assign wr_req_desc_e_wuser_10_wuser_f = wr_req_desc_e_wuser_10_reg[31:0];
   assign wr_req_desc_e_wuser_11_wuser_f = wr_req_desc_e_wuser_11_reg[31:0];
   assign wr_req_desc_e_wuser_12_wuser_f = wr_req_desc_e_wuser_12_reg[31:0];
   assign wr_req_desc_e_wuser_13_wuser_f = wr_req_desc_e_wuser_13_reg[31:0];
   assign wr_req_desc_e_wuser_14_wuser_f = wr_req_desc_e_wuser_14_reg[31:0];
   assign wr_req_desc_e_wuser_15_wuser_f = wr_req_desc_e_wuser_15_reg[31:0];
   assign wr_resp_desc_e_resp_resp_f = wr_resp_desc_e_resp_reg[4:0];
   assign wr_resp_desc_e_xid_0_xid_f = wr_resp_desc_e_xid_0_reg[31:0];
   assign wr_resp_desc_e_xid_1_xid_f = wr_resp_desc_e_xid_1_reg[31:0];
   assign wr_resp_desc_e_xid_2_xid_f = wr_resp_desc_e_xid_2_reg[31:0];
   assign wr_resp_desc_e_xid_3_xid_f = wr_resp_desc_e_xid_3_reg[31:0];
   assign wr_resp_desc_e_xuser_0_xuser_f = wr_resp_desc_e_xuser_0_reg[31:0];
   assign wr_resp_desc_e_xuser_1_xuser_f = wr_resp_desc_e_xuser_1_reg[31:0];
   assign wr_resp_desc_e_xuser_2_xuser_f = wr_resp_desc_e_xuser_2_reg[31:0];
   assign wr_resp_desc_e_xuser_3_xuser_f = wr_resp_desc_e_xuser_3_reg[31:0];
   assign wr_resp_desc_e_xuser_4_xuser_f = wr_resp_desc_e_xuser_4_reg[31:0];
   assign wr_resp_desc_e_xuser_5_xuser_f = wr_resp_desc_e_xuser_5_reg[31:0];
   assign wr_resp_desc_e_xuser_6_xuser_f = wr_resp_desc_e_xuser_6_reg[31:0];
   assign wr_resp_desc_e_xuser_7_xuser_f = wr_resp_desc_e_xuser_7_reg[31:0];
   assign wr_resp_desc_e_xuser_8_xuser_f = wr_resp_desc_e_xuser_8_reg[31:0];
   assign wr_resp_desc_e_xuser_9_xuser_f = wr_resp_desc_e_xuser_9_reg[31:0];
   assign wr_resp_desc_e_xuser_10_xuser_f = wr_resp_desc_e_xuser_10_reg[31:0];
   assign wr_resp_desc_e_xuser_11_xuser_f = wr_resp_desc_e_xuser_11_reg[31:0];
   assign wr_resp_desc_e_xuser_12_xuser_f = wr_resp_desc_e_xuser_12_reg[31:0];
   assign wr_resp_desc_e_xuser_13_xuser_f = wr_resp_desc_e_xuser_13_reg[31:0];
   assign wr_resp_desc_e_xuser_14_xuser_f = wr_resp_desc_e_xuser_14_reg[31:0];
   assign wr_resp_desc_e_xuser_15_xuser_f = wr_resp_desc_e_xuser_15_reg[31:0];
   assign sn_req_desc_e_attr_acsnoop_f = sn_req_desc_e_attr_reg[27:24];
   assign sn_req_desc_e_attr_acprot_f = sn_req_desc_e_attr_reg[10:8];
   assign sn_req_desc_e_acaddr_0_addr_f = sn_req_desc_e_acaddr_0_reg[31:0];
   assign sn_req_desc_e_acaddr_1_addr_f = sn_req_desc_e_acaddr_1_reg[31:0];
   assign sn_req_desc_e_acaddr_2_addr_f = sn_req_desc_e_acaddr_2_reg[31:0];
   assign sn_req_desc_e_acaddr_3_addr_f = sn_req_desc_e_acaddr_3_reg[31:0];
   assign sn_resp_desc_e_resp_resp_f = sn_resp_desc_e_resp_reg[4:0];
   assign rd_req_desc_f_size_txn_size_f = rd_req_desc_f_size_reg[31:0];
   assign rd_req_desc_f_axsize_axsize_f = rd_req_desc_f_axsize_reg[2:0];
   assign rd_req_desc_f_attr_axsnoop_f = rd_req_desc_f_attr_reg[27:24];
   assign rd_req_desc_f_attr_axdomain_f = rd_req_desc_f_attr_reg[23:22];
   assign rd_req_desc_f_attr_axbar_f = rd_req_desc_f_attr_reg[21:20];
   assign rd_req_desc_f_attr_axregion_f = rd_req_desc_f_attr_reg[18:15];
   assign rd_req_desc_f_attr_axqos_f = rd_req_desc_f_attr_reg[14:11];
   assign rd_req_desc_f_attr_axprot_f = rd_req_desc_f_attr_reg[10:8];
   assign rd_req_desc_f_attr_axcache_f = rd_req_desc_f_attr_reg[7:4];
   assign rd_req_desc_f_attr_axlock_f = rd_req_desc_f_attr_reg[2];
   assign rd_req_desc_f_attr_axburst_f = rd_req_desc_f_attr_reg[1:0];
   assign rd_req_desc_f_axaddr_0_addr_f = rd_req_desc_f_axaddr_0_reg[31:0];
   assign rd_req_desc_f_axaddr_1_addr_f = rd_req_desc_f_axaddr_1_reg[31:0];
   assign rd_req_desc_f_axaddr_2_addr_f = rd_req_desc_f_axaddr_2_reg[31:0];
   assign rd_req_desc_f_axaddr_3_addr_f = rd_req_desc_f_axaddr_3_reg[31:0];
   assign rd_req_desc_f_axid_0_axid_f = rd_req_desc_f_axid_0_reg[31:0];
   assign rd_req_desc_f_axid_1_axid_f = rd_req_desc_f_axid_1_reg[31:0];
   assign rd_req_desc_f_axid_2_axid_f = rd_req_desc_f_axid_2_reg[31:0];
   assign rd_req_desc_f_axid_3_axid_f = rd_req_desc_f_axid_3_reg[31:0];
   assign rd_req_desc_f_axuser_0_axuser_f = rd_req_desc_f_axuser_0_reg[31:0];
   assign rd_req_desc_f_axuser_1_axuser_f = rd_req_desc_f_axuser_1_reg[31:0];
   assign rd_req_desc_f_axuser_2_axuser_f = rd_req_desc_f_axuser_2_reg[31:0];
   assign rd_req_desc_f_axuser_3_axuser_f = rd_req_desc_f_axuser_3_reg[31:0];
   assign rd_req_desc_f_axuser_4_axuser_f = rd_req_desc_f_axuser_4_reg[31:0];
   assign rd_req_desc_f_axuser_5_axuser_f = rd_req_desc_f_axuser_5_reg[31:0];
   assign rd_req_desc_f_axuser_6_axuser_f = rd_req_desc_f_axuser_6_reg[31:0];
   assign rd_req_desc_f_axuser_7_axuser_f = rd_req_desc_f_axuser_7_reg[31:0];
   assign rd_req_desc_f_axuser_8_axuser_f = rd_req_desc_f_axuser_8_reg[31:0];
   assign rd_req_desc_f_axuser_9_axuser_f = rd_req_desc_f_axuser_9_reg[31:0];
   assign rd_req_desc_f_axuser_10_axuser_f = rd_req_desc_f_axuser_10_reg[31:0];
   assign rd_req_desc_f_axuser_11_axuser_f = rd_req_desc_f_axuser_11_reg[31:0];
   assign rd_req_desc_f_axuser_12_axuser_f = rd_req_desc_f_axuser_12_reg[31:0];
   assign rd_req_desc_f_axuser_13_axuser_f = rd_req_desc_f_axuser_13_reg[31:0];
   assign rd_req_desc_f_axuser_14_axuser_f = rd_req_desc_f_axuser_14_reg[31:0];
   assign rd_req_desc_f_axuser_15_axuser_f = rd_req_desc_f_axuser_15_reg[31:0];
   assign rd_resp_desc_f_data_offset_addr_f = rd_resp_desc_f_data_offset_reg[13:0];
   assign rd_resp_desc_f_data_size_size_f = rd_resp_desc_f_data_size_reg[31:0];
   assign rd_resp_desc_f_data_host_addr_0_addr_f = rd_resp_desc_f_data_host_addr_0_reg[31:0];
   assign rd_resp_desc_f_data_host_addr_1_addr_f = rd_resp_desc_f_data_host_addr_1_reg[31:0];
   assign rd_resp_desc_f_data_host_addr_2_addr_f = rd_resp_desc_f_data_host_addr_2_reg[31:0];
   assign rd_resp_desc_f_data_host_addr_3_addr_f = rd_resp_desc_f_data_host_addr_3_reg[31:0];
   assign rd_resp_desc_f_resp_resp_f = rd_resp_desc_f_resp_reg[4:0];
   assign rd_resp_desc_f_xid_0_xid_f = rd_resp_desc_f_xid_0_reg[31:0];
   assign rd_resp_desc_f_xid_1_xid_f = rd_resp_desc_f_xid_1_reg[31:0];
   assign rd_resp_desc_f_xid_2_xid_f = rd_resp_desc_f_xid_2_reg[31:0];
   assign rd_resp_desc_f_xid_3_xid_f = rd_resp_desc_f_xid_3_reg[31:0];
   assign rd_resp_desc_f_xuser_0_xuser_f = rd_resp_desc_f_xuser_0_reg[31:0];
   assign rd_resp_desc_f_xuser_1_xuser_f = rd_resp_desc_f_xuser_1_reg[31:0];
   assign rd_resp_desc_f_xuser_2_xuser_f = rd_resp_desc_f_xuser_2_reg[31:0];
   assign rd_resp_desc_f_xuser_3_xuser_f = rd_resp_desc_f_xuser_3_reg[31:0];
   assign rd_resp_desc_f_xuser_4_xuser_f = rd_resp_desc_f_xuser_4_reg[31:0];
   assign rd_resp_desc_f_xuser_5_xuser_f = rd_resp_desc_f_xuser_5_reg[31:0];
   assign rd_resp_desc_f_xuser_6_xuser_f = rd_resp_desc_f_xuser_6_reg[31:0];
   assign rd_resp_desc_f_xuser_7_xuser_f = rd_resp_desc_f_xuser_7_reg[31:0];
   assign rd_resp_desc_f_xuser_8_xuser_f = rd_resp_desc_f_xuser_8_reg[31:0];
   assign rd_resp_desc_f_xuser_9_xuser_f = rd_resp_desc_f_xuser_9_reg[31:0];
   assign rd_resp_desc_f_xuser_10_xuser_f = rd_resp_desc_f_xuser_10_reg[31:0];
   assign rd_resp_desc_f_xuser_11_xuser_f = rd_resp_desc_f_xuser_11_reg[31:0];
   assign rd_resp_desc_f_xuser_12_xuser_f = rd_resp_desc_f_xuser_12_reg[31:0];
   assign rd_resp_desc_f_xuser_13_xuser_f = rd_resp_desc_f_xuser_13_reg[31:0];
   assign rd_resp_desc_f_xuser_14_xuser_f = rd_resp_desc_f_xuser_14_reg[31:0];
   assign rd_resp_desc_f_xuser_15_xuser_f = rd_resp_desc_f_xuser_15_reg[31:0];
   assign wr_req_desc_f_txn_type_wr_strb_f = wr_req_desc_f_txn_type_reg[1];
   assign wr_req_desc_f_size_txn_size_f = wr_req_desc_f_size_reg[31:0];
   assign wr_req_desc_f_data_offset_addr_f = wr_req_desc_f_data_offset_reg[13:0];
   assign wr_req_desc_f_data_host_addr_0_addr_f = wr_req_desc_f_data_host_addr_0_reg[31:0];
   assign wr_req_desc_f_data_host_addr_1_addr_f = wr_req_desc_f_data_host_addr_1_reg[31:0];
   assign wr_req_desc_f_data_host_addr_2_addr_f = wr_req_desc_f_data_host_addr_2_reg[31:0];
   assign wr_req_desc_f_data_host_addr_3_addr_f = wr_req_desc_f_data_host_addr_3_reg[31:0];
   assign wr_req_desc_f_wstrb_host_addr_0_addr_f = wr_req_desc_f_wstrb_host_addr_0_reg[31:0];
   assign wr_req_desc_f_wstrb_host_addr_1_addr_f = wr_req_desc_f_wstrb_host_addr_1_reg[31:0];
   assign wr_req_desc_f_wstrb_host_addr_2_addr_f = wr_req_desc_f_wstrb_host_addr_2_reg[31:0];
   assign wr_req_desc_f_wstrb_host_addr_3_addr_f = wr_req_desc_f_wstrb_host_addr_3_reg[31:0];
   assign wr_req_desc_f_axsize_axsize_f = wr_req_desc_f_axsize_reg[2:0];
   assign wr_req_desc_f_attr_axsnoop_f = wr_req_desc_f_attr_reg[27:24];
   assign wr_req_desc_f_attr_axdomain_f = wr_req_desc_f_attr_reg[23:22];
   assign wr_req_desc_f_attr_axbar_f = wr_req_desc_f_attr_reg[21:20];
   assign wr_req_desc_f_attr_awunique_f = wr_req_desc_f_attr_reg[19];
   assign wr_req_desc_f_attr_axregion_f = wr_req_desc_f_attr_reg[18:15];
   assign wr_req_desc_f_attr_axqos_f = wr_req_desc_f_attr_reg[14:11];
   assign wr_req_desc_f_attr_axprot_f = wr_req_desc_f_attr_reg[10:8];
   assign wr_req_desc_f_attr_axcache_f = wr_req_desc_f_attr_reg[7:4];
   assign wr_req_desc_f_attr_axlock_f = wr_req_desc_f_attr_reg[2];
   assign wr_req_desc_f_attr_axburst_f = wr_req_desc_f_attr_reg[1:0];
   assign wr_req_desc_f_axaddr_0_addr_f = wr_req_desc_f_axaddr_0_reg[31:0];
   assign wr_req_desc_f_axaddr_1_addr_f = wr_req_desc_f_axaddr_1_reg[31:0];
   assign wr_req_desc_f_axaddr_2_addr_f = wr_req_desc_f_axaddr_2_reg[31:0];
   assign wr_req_desc_f_axaddr_3_addr_f = wr_req_desc_f_axaddr_3_reg[31:0];
   assign wr_req_desc_f_axid_0_axid_f = wr_req_desc_f_axid_0_reg[31:0];
   assign wr_req_desc_f_axid_1_axid_f = wr_req_desc_f_axid_1_reg[31:0];
   assign wr_req_desc_f_axid_2_axid_f = wr_req_desc_f_axid_2_reg[31:0];
   assign wr_req_desc_f_axid_3_axid_f = wr_req_desc_f_axid_3_reg[31:0];
   assign wr_req_desc_f_axuser_0_axuser_f = wr_req_desc_f_axuser_0_reg[31:0];
   assign wr_req_desc_f_axuser_1_axuser_f = wr_req_desc_f_axuser_1_reg[31:0];
   assign wr_req_desc_f_axuser_2_axuser_f = wr_req_desc_f_axuser_2_reg[31:0];
   assign wr_req_desc_f_axuser_3_axuser_f = wr_req_desc_f_axuser_3_reg[31:0];
   assign wr_req_desc_f_axuser_4_axuser_f = wr_req_desc_f_axuser_4_reg[31:0];
   assign wr_req_desc_f_axuser_5_axuser_f = wr_req_desc_f_axuser_5_reg[31:0];
   assign wr_req_desc_f_axuser_6_axuser_f = wr_req_desc_f_axuser_6_reg[31:0];
   assign wr_req_desc_f_axuser_7_axuser_f = wr_req_desc_f_axuser_7_reg[31:0];
   assign wr_req_desc_f_axuser_8_axuser_f = wr_req_desc_f_axuser_8_reg[31:0];
   assign wr_req_desc_f_axuser_9_axuser_f = wr_req_desc_f_axuser_9_reg[31:0];
   assign wr_req_desc_f_axuser_10_axuser_f = wr_req_desc_f_axuser_10_reg[31:0];
   assign wr_req_desc_f_axuser_11_axuser_f = wr_req_desc_f_axuser_11_reg[31:0];
   assign wr_req_desc_f_axuser_12_axuser_f = wr_req_desc_f_axuser_12_reg[31:0];
   assign wr_req_desc_f_axuser_13_axuser_f = wr_req_desc_f_axuser_13_reg[31:0];
   assign wr_req_desc_f_axuser_14_axuser_f = wr_req_desc_f_axuser_14_reg[31:0];
   assign wr_req_desc_f_axuser_15_axuser_f = wr_req_desc_f_axuser_15_reg[31:0];
   assign wr_req_desc_f_wuser_0_wuser_f = wr_req_desc_f_wuser_0_reg[31:0];
   assign wr_req_desc_f_wuser_1_wuser_f = wr_req_desc_f_wuser_1_reg[31:0];
   assign wr_req_desc_f_wuser_2_wuser_f = wr_req_desc_f_wuser_2_reg[31:0];
   assign wr_req_desc_f_wuser_3_wuser_f = wr_req_desc_f_wuser_3_reg[31:0];
   assign wr_req_desc_f_wuser_4_wuser_f = wr_req_desc_f_wuser_4_reg[31:0];
   assign wr_req_desc_f_wuser_5_wuser_f = wr_req_desc_f_wuser_5_reg[31:0];
   assign wr_req_desc_f_wuser_6_wuser_f = wr_req_desc_f_wuser_6_reg[31:0];
   assign wr_req_desc_f_wuser_7_wuser_f = wr_req_desc_f_wuser_7_reg[31:0];
   assign wr_req_desc_f_wuser_8_wuser_f = wr_req_desc_f_wuser_8_reg[31:0];
   assign wr_req_desc_f_wuser_9_wuser_f = wr_req_desc_f_wuser_9_reg[31:0];
   assign wr_req_desc_f_wuser_10_wuser_f = wr_req_desc_f_wuser_10_reg[31:0];
   assign wr_req_desc_f_wuser_11_wuser_f = wr_req_desc_f_wuser_11_reg[31:0];
   assign wr_req_desc_f_wuser_12_wuser_f = wr_req_desc_f_wuser_12_reg[31:0];
   assign wr_req_desc_f_wuser_13_wuser_f = wr_req_desc_f_wuser_13_reg[31:0];
   assign wr_req_desc_f_wuser_14_wuser_f = wr_req_desc_f_wuser_14_reg[31:0];
   assign wr_req_desc_f_wuser_15_wuser_f = wr_req_desc_f_wuser_15_reg[31:0];
   assign wr_resp_desc_f_resp_resp_f = wr_resp_desc_f_resp_reg[4:0];
   assign wr_resp_desc_f_xid_0_xid_f = wr_resp_desc_f_xid_0_reg[31:0];
   assign wr_resp_desc_f_xid_1_xid_f = wr_resp_desc_f_xid_1_reg[31:0];
   assign wr_resp_desc_f_xid_2_xid_f = wr_resp_desc_f_xid_2_reg[31:0];
   assign wr_resp_desc_f_xid_3_xid_f = wr_resp_desc_f_xid_3_reg[31:0];
   assign wr_resp_desc_f_xuser_0_xuser_f = wr_resp_desc_f_xuser_0_reg[31:0];
   assign wr_resp_desc_f_xuser_1_xuser_f = wr_resp_desc_f_xuser_1_reg[31:0];
   assign wr_resp_desc_f_xuser_2_xuser_f = wr_resp_desc_f_xuser_2_reg[31:0];
   assign wr_resp_desc_f_xuser_3_xuser_f = wr_resp_desc_f_xuser_3_reg[31:0];
   assign wr_resp_desc_f_xuser_4_xuser_f = wr_resp_desc_f_xuser_4_reg[31:0];
   assign wr_resp_desc_f_xuser_5_xuser_f = wr_resp_desc_f_xuser_5_reg[31:0];
   assign wr_resp_desc_f_xuser_6_xuser_f = wr_resp_desc_f_xuser_6_reg[31:0];
   assign wr_resp_desc_f_xuser_7_xuser_f = wr_resp_desc_f_xuser_7_reg[31:0];
   assign wr_resp_desc_f_xuser_8_xuser_f = wr_resp_desc_f_xuser_8_reg[31:0];
   assign wr_resp_desc_f_xuser_9_xuser_f = wr_resp_desc_f_xuser_9_reg[31:0];
   assign wr_resp_desc_f_xuser_10_xuser_f = wr_resp_desc_f_xuser_10_reg[31:0];
   assign wr_resp_desc_f_xuser_11_xuser_f = wr_resp_desc_f_xuser_11_reg[31:0];
   assign wr_resp_desc_f_xuser_12_xuser_f = wr_resp_desc_f_xuser_12_reg[31:0];
   assign wr_resp_desc_f_xuser_13_xuser_f = wr_resp_desc_f_xuser_13_reg[31:0];
   assign wr_resp_desc_f_xuser_14_xuser_f = wr_resp_desc_f_xuser_14_reg[31:0];
   assign wr_resp_desc_f_xuser_15_xuser_f = wr_resp_desc_f_xuser_15_reg[31:0];
   assign sn_req_desc_f_attr_acsnoop_f = sn_req_desc_f_attr_reg[27:24];
   assign sn_req_desc_f_attr_acprot_f = sn_req_desc_f_attr_reg[10:8];
   assign sn_req_desc_f_acaddr_0_addr_f = sn_req_desc_f_acaddr_0_reg[31:0];
   assign sn_req_desc_f_acaddr_1_addr_f = sn_req_desc_f_acaddr_1_reg[31:0];
   assign sn_req_desc_f_acaddr_2_addr_f = sn_req_desc_f_acaddr_2_reg[31:0];
   assign sn_req_desc_f_acaddr_3_addr_f = sn_req_desc_f_acaddr_3_reg[31:0];
   assign sn_resp_desc_f_resp_resp_f = sn_resp_desc_f_resp_reg[4:0];


   //Assign signals to use in entire slave RTL ( int_<reg>_<field> )

   assign int_bridge_identification_last_bridge = bridge_identification_last_bridge_f;
   assign int_version_major_ver = version_major_ver_f;
   assign int_version_minor_ver = version_minor_ver_f;
   assign int_bridge_type_type = bridge_type_type_f;
   assign int_bridge_config_extend_wstrb = bridge_config_extend_wstrb_f;
   assign int_bridge_config_id_width = bridge_config_id_width_f;
   assign int_bridge_config_data_width = bridge_config_data_width_f;
   assign int_bridge_rd_user_config_ruser_width = bridge_rd_user_config_ruser_width_f;
   assign int_bridge_rd_user_config_aruser_width = bridge_rd_user_config_aruser_width_f;
   assign int_bridge_wr_user_config_buser_width = bridge_wr_user_config_buser_width_f;
   assign int_bridge_wr_user_config_wuser_width = bridge_wr_user_config_wuser_width_f;
   assign int_bridge_wr_user_config_awuser_width = bridge_wr_user_config_awuser_width_f;
   assign int_rd_max_desc_resp_max_desc = rd_max_desc_resp_max_desc_f;
   assign int_rd_max_desc_req_max_desc = rd_max_desc_req_max_desc_f;
   assign int_wr_max_desc_resp_max_desc = wr_max_desc_resp_max_desc_f;
   assign int_wr_max_desc_req_max_desc = wr_max_desc_req_max_desc_f;
   assign int_sn_max_desc_data_max_desc = sn_max_desc_data_max_desc_f;
   assign int_sn_max_desc_resp_max_desc = sn_max_desc_resp_max_desc_f;
   assign int_sn_max_desc_req_max_desc = sn_max_desc_req_max_desc_f;
   assign int_reset_dut_srst_3 = reset_dut_srst_3_f;
   assign int_reset_dut_srst_2 = reset_dut_srst_2_f;
   assign int_reset_dut_srst_1 = reset_dut_srst_1_f;
   assign int_reset_dut_srst_0 = reset_dut_srst_0_f;
   assign int_reset_srst = reset_srst_f;
   assign int_mode_select_mode_0_1 = mode_select_mode_0_1_f;
   assign int_intr_status_sn_data_fifo_nonempty = intr_status_sn_data_fifo_nonempty_f;
   assign int_intr_status_sn_resp_fifo_nonempty = intr_status_sn_resp_fifo_nonempty_f;
   assign int_intr_status_sn_req_comp = intr_status_sn_req_comp_f;
   assign int_intr_status_wr_resp_comp = intr_status_wr_resp_comp_f;
   assign int_intr_status_wr_req_fifo_nonempty = intr_status_wr_req_fifo_nonempty_f;
   assign int_intr_status_rd_resp_comp = intr_status_rd_resp_comp_f;
   assign int_intr_status_rd_req_fifo_nonempty = intr_status_rd_req_fifo_nonempty_f;
   assign int_intr_status_c2h = intr_status_c2h_f;
   assign int_intr_status_error = intr_status_error_f;
   assign int_intr_error_status_err_1 = intr_error_status_err_1_f;
   assign int_intr_error_clear_clr_err_2 = intr_error_clear_clr_err_2_f;
   assign int_intr_error_clear_clr_err_1 = intr_error_clear_clr_err_1_f;
   assign int_intr_error_clear_clr_err_0 = intr_error_clear_clr_err_0_f;
   assign int_intr_error_enable_en_err_2 = intr_error_enable_en_err_2_f;
   assign int_intr_error_enable_en_err_1 = intr_error_enable_en_err_1_f;
   assign int_intr_error_enable_en_err_0 = intr_error_enable_en_err_0_f;
   assign int_rd_req_free_desc_desc = rd_req_free_desc_desc_f;
   assign int_rd_resp_fifo_push_desc_valid = rd_resp_fifo_push_desc_valid_f;
   assign int_rd_resp_fifo_push_desc_desc_index = rd_resp_fifo_push_desc_desc_index_f;
   assign int_rd_resp_intr_comp_clear_clr_comp = rd_resp_intr_comp_clear_clr_comp_f;
   assign int_rd_resp_intr_comp_enable_en_comp = rd_resp_intr_comp_enable_en_comp_f;
   assign int_wr_req_free_desc_desc = wr_req_free_desc_desc_f;
   assign int_wr_resp_fifo_push_desc_valid = wr_resp_fifo_push_desc_valid_f;
   assign int_wr_resp_fifo_push_desc_desc_index = wr_resp_fifo_push_desc_desc_index_f;
   assign int_wr_resp_intr_comp_clear_clr_comp = wr_resp_intr_comp_clear_clr_comp_f;
   assign int_wr_resp_intr_comp_enable_en_comp = wr_resp_intr_comp_enable_en_comp_f;
   assign int_sn_req_fifo_push_desc_valid = sn_req_fifo_push_desc_valid_f;
   assign int_sn_req_fifo_push_desc_desc_index = sn_req_fifo_push_desc_desc_index_f;
   assign int_sn_req_intr_comp_clear_clr_comp = sn_req_intr_comp_clear_clr_comp_f;
   assign int_sn_req_intr_comp_enable_en_comp = sn_req_intr_comp_enable_en_comp_f;
   assign int_sn_resp_free_desc_desc = sn_resp_free_desc_desc_f;
   assign int_sn_data_free_desc_desc = sn_data_free_desc_desc_f;
   assign int_intr_fifo_enable_en_sn_data_fifo_nonempty = intr_fifo_enable_en_sn_data_fifo_nonempty_f;
   assign int_intr_fifo_enable_en_sn_resp_fifo_nonempty = intr_fifo_enable_en_sn_resp_fifo_nonempty_f;
   assign int_intr_fifo_enable_en_wr_req_fifo_nonempty = intr_fifo_enable_en_wr_req_fifo_nonempty_f;
   assign int_intr_fifo_enable_en_rd_req_fifo_nonempty = intr_fifo_enable_en_rd_req_fifo_nonempty_f;
   assign int_h2c_intr_0_h2c_31 = h2c_intr_0_h2c_31_f;
   assign int_h2c_intr_0_h2c_30 = h2c_intr_0_h2c_30_f;
   assign int_h2c_intr_0_h2c_29 = h2c_intr_0_h2c_29_f;
   assign int_h2c_intr_0_h2c_28 = h2c_intr_0_h2c_28_f;
   assign int_h2c_intr_0_h2c_27 = h2c_intr_0_h2c_27_f;
   assign int_h2c_intr_0_h2c_26 = h2c_intr_0_h2c_26_f;
   assign int_h2c_intr_0_h2c_25 = h2c_intr_0_h2c_25_f;
   assign int_h2c_intr_0_h2c_24 = h2c_intr_0_h2c_24_f;
   assign int_h2c_intr_0_h2c_23 = h2c_intr_0_h2c_23_f;
   assign int_h2c_intr_0_h2c_22 = h2c_intr_0_h2c_22_f;
   assign int_h2c_intr_0_h2c_21 = h2c_intr_0_h2c_21_f;
   assign int_h2c_intr_0_h2c_20 = h2c_intr_0_h2c_20_f;
   assign int_h2c_intr_0_h2c_19 = h2c_intr_0_h2c_19_f;
   assign int_h2c_intr_0_h2c_18 = h2c_intr_0_h2c_18_f;
   assign int_h2c_intr_0_h2c_17 = h2c_intr_0_h2c_17_f;
   assign int_h2c_intr_0_h2c_16 = h2c_intr_0_h2c_16_f;
   assign int_h2c_intr_0_h2c_15 = h2c_intr_0_h2c_15_f;
   assign int_h2c_intr_0_h2c_14 = h2c_intr_0_h2c_14_f;
   assign int_h2c_intr_0_h2c_13 = h2c_intr_0_h2c_13_f;
   assign int_h2c_intr_0_h2c_12 = h2c_intr_0_h2c_12_f;
   assign int_h2c_intr_0_h2c_11 = h2c_intr_0_h2c_11_f;
   assign int_h2c_intr_0_h2c_10 = h2c_intr_0_h2c_10_f;
   assign int_h2c_intr_0_h2c_9 = h2c_intr_0_h2c_9_f;
   assign int_h2c_intr_0_h2c_8 = h2c_intr_0_h2c_8_f;
   assign int_h2c_intr_0_h2c_7 = h2c_intr_0_h2c_7_f;
   assign int_h2c_intr_0_h2c_6 = h2c_intr_0_h2c_6_f;
   assign int_h2c_intr_0_h2c_5 = h2c_intr_0_h2c_5_f;
   assign int_h2c_intr_0_h2c_4 = h2c_intr_0_h2c_4_f;
   assign int_h2c_intr_0_h2c_3 = h2c_intr_0_h2c_3_f;
   assign int_h2c_intr_0_h2c_2 = h2c_intr_0_h2c_2_f;
   assign int_h2c_intr_0_h2c_1 = h2c_intr_0_h2c_1_f;
   assign int_h2c_intr_0_h2c_0 = h2c_intr_0_h2c_0_f;
   assign int_h2c_intr_1_h2c_31 = h2c_intr_1_h2c_31_f;
   assign int_h2c_intr_1_h2c_30 = h2c_intr_1_h2c_30_f;
   assign int_h2c_intr_1_h2c_29 = h2c_intr_1_h2c_29_f;
   assign int_h2c_intr_1_h2c_28 = h2c_intr_1_h2c_28_f;
   assign int_h2c_intr_1_h2c_27 = h2c_intr_1_h2c_27_f;
   assign int_h2c_intr_1_h2c_26 = h2c_intr_1_h2c_26_f;
   assign int_h2c_intr_1_h2c_25 = h2c_intr_1_h2c_25_f;
   assign int_h2c_intr_1_h2c_24 = h2c_intr_1_h2c_24_f;
   assign int_h2c_intr_1_h2c_23 = h2c_intr_1_h2c_23_f;
   assign int_h2c_intr_1_h2c_22 = h2c_intr_1_h2c_22_f;
   assign int_h2c_intr_1_h2c_21 = h2c_intr_1_h2c_21_f;
   assign int_h2c_intr_1_h2c_20 = h2c_intr_1_h2c_20_f;
   assign int_h2c_intr_1_h2c_19 = h2c_intr_1_h2c_19_f;
   assign int_h2c_intr_1_h2c_18 = h2c_intr_1_h2c_18_f;
   assign int_h2c_intr_1_h2c_17 = h2c_intr_1_h2c_17_f;
   assign int_h2c_intr_1_h2c_16 = h2c_intr_1_h2c_16_f;
   assign int_h2c_intr_1_h2c_15 = h2c_intr_1_h2c_15_f;
   assign int_h2c_intr_1_h2c_14 = h2c_intr_1_h2c_14_f;
   assign int_h2c_intr_1_h2c_13 = h2c_intr_1_h2c_13_f;
   assign int_h2c_intr_1_h2c_12 = h2c_intr_1_h2c_12_f;
   assign int_h2c_intr_1_h2c_11 = h2c_intr_1_h2c_11_f;
   assign int_h2c_intr_1_h2c_10 = h2c_intr_1_h2c_10_f;
   assign int_h2c_intr_1_h2c_9 = h2c_intr_1_h2c_9_f;
   assign int_h2c_intr_1_h2c_8 = h2c_intr_1_h2c_8_f;
   assign int_h2c_intr_1_h2c_7 = h2c_intr_1_h2c_7_f;
   assign int_h2c_intr_1_h2c_6 = h2c_intr_1_h2c_6_f;
   assign int_h2c_intr_1_h2c_5 = h2c_intr_1_h2c_5_f;
   assign int_h2c_intr_1_h2c_4 = h2c_intr_1_h2c_4_f;
   assign int_h2c_intr_1_h2c_3 = h2c_intr_1_h2c_3_f;
   assign int_h2c_intr_1_h2c_2 = h2c_intr_1_h2c_2_f;
   assign int_h2c_intr_1_h2c_1 = h2c_intr_1_h2c_1_f;
   assign int_h2c_intr_1_h2c_0 = h2c_intr_1_h2c_0_f;
   assign int_h2c_intr_2_h2c_31 = h2c_intr_2_h2c_31_f;
   assign int_h2c_intr_2_h2c_30 = h2c_intr_2_h2c_30_f;
   assign int_h2c_intr_2_h2c_29 = h2c_intr_2_h2c_29_f;
   assign int_h2c_intr_2_h2c_28 = h2c_intr_2_h2c_28_f;
   assign int_h2c_intr_2_h2c_27 = h2c_intr_2_h2c_27_f;
   assign int_h2c_intr_2_h2c_26 = h2c_intr_2_h2c_26_f;
   assign int_h2c_intr_2_h2c_25 = h2c_intr_2_h2c_25_f;
   assign int_h2c_intr_2_h2c_24 = h2c_intr_2_h2c_24_f;
   assign int_h2c_intr_2_h2c_23 = h2c_intr_2_h2c_23_f;
   assign int_h2c_intr_2_h2c_22 = h2c_intr_2_h2c_22_f;
   assign int_h2c_intr_2_h2c_21 = h2c_intr_2_h2c_21_f;
   assign int_h2c_intr_2_h2c_20 = h2c_intr_2_h2c_20_f;
   assign int_h2c_intr_2_h2c_19 = h2c_intr_2_h2c_19_f;
   assign int_h2c_intr_2_h2c_18 = h2c_intr_2_h2c_18_f;
   assign int_h2c_intr_2_h2c_17 = h2c_intr_2_h2c_17_f;
   assign int_h2c_intr_2_h2c_16 = h2c_intr_2_h2c_16_f;
   assign int_h2c_intr_2_h2c_15 = h2c_intr_2_h2c_15_f;
   assign int_h2c_intr_2_h2c_14 = h2c_intr_2_h2c_14_f;
   assign int_h2c_intr_2_h2c_13 = h2c_intr_2_h2c_13_f;
   assign int_h2c_intr_2_h2c_12 = h2c_intr_2_h2c_12_f;
   assign int_h2c_intr_2_h2c_11 = h2c_intr_2_h2c_11_f;
   assign int_h2c_intr_2_h2c_10 = h2c_intr_2_h2c_10_f;
   assign int_h2c_intr_2_h2c_9 = h2c_intr_2_h2c_9_f;
   assign int_h2c_intr_2_h2c_8 = h2c_intr_2_h2c_8_f;
   assign int_h2c_intr_2_h2c_7 = h2c_intr_2_h2c_7_f;
   assign int_h2c_intr_2_h2c_6 = h2c_intr_2_h2c_6_f;
   assign int_h2c_intr_2_h2c_5 = h2c_intr_2_h2c_5_f;
   assign int_h2c_intr_2_h2c_4 = h2c_intr_2_h2c_4_f;
   assign int_h2c_intr_2_h2c_3 = h2c_intr_2_h2c_3_f;
   assign int_h2c_intr_2_h2c_2 = h2c_intr_2_h2c_2_f;
   assign int_h2c_intr_2_h2c_1 = h2c_intr_2_h2c_1_f;
   assign int_h2c_intr_2_h2c_0 = h2c_intr_2_h2c_0_f;
   assign int_h2c_intr_3_h2c_31 = h2c_intr_3_h2c_31_f;
   assign int_h2c_intr_3_h2c_30 = h2c_intr_3_h2c_30_f;
   assign int_h2c_intr_3_h2c_29 = h2c_intr_3_h2c_29_f;
   assign int_h2c_intr_3_h2c_28 = h2c_intr_3_h2c_28_f;
   assign int_h2c_intr_3_h2c_27 = h2c_intr_3_h2c_27_f;
   assign int_h2c_intr_3_h2c_26 = h2c_intr_3_h2c_26_f;
   assign int_h2c_intr_3_h2c_25 = h2c_intr_3_h2c_25_f;
   assign int_h2c_intr_3_h2c_24 = h2c_intr_3_h2c_24_f;
   assign int_h2c_intr_3_h2c_23 = h2c_intr_3_h2c_23_f;
   assign int_h2c_intr_3_h2c_22 = h2c_intr_3_h2c_22_f;
   assign int_h2c_intr_3_h2c_21 = h2c_intr_3_h2c_21_f;
   assign int_h2c_intr_3_h2c_20 = h2c_intr_3_h2c_20_f;
   assign int_h2c_intr_3_h2c_19 = h2c_intr_3_h2c_19_f;
   assign int_h2c_intr_3_h2c_18 = h2c_intr_3_h2c_18_f;
   assign int_h2c_intr_3_h2c_17 = h2c_intr_3_h2c_17_f;
   assign int_h2c_intr_3_h2c_16 = h2c_intr_3_h2c_16_f;
   assign int_h2c_intr_3_h2c_15 = h2c_intr_3_h2c_15_f;
   assign int_h2c_intr_3_h2c_14 = h2c_intr_3_h2c_14_f;
   assign int_h2c_intr_3_h2c_13 = h2c_intr_3_h2c_13_f;
   assign int_h2c_intr_3_h2c_12 = h2c_intr_3_h2c_12_f;
   assign int_h2c_intr_3_h2c_11 = h2c_intr_3_h2c_11_f;
   assign int_h2c_intr_3_h2c_10 = h2c_intr_3_h2c_10_f;
   assign int_h2c_intr_3_h2c_9 = h2c_intr_3_h2c_9_f;
   assign int_h2c_intr_3_h2c_8 = h2c_intr_3_h2c_8_f;
   assign int_h2c_intr_3_h2c_7 = h2c_intr_3_h2c_7_f;
   assign int_h2c_intr_3_h2c_6 = h2c_intr_3_h2c_6_f;
   assign int_h2c_intr_3_h2c_5 = h2c_intr_3_h2c_5_f;
   assign int_h2c_intr_3_h2c_4 = h2c_intr_3_h2c_4_f;
   assign int_h2c_intr_3_h2c_3 = h2c_intr_3_h2c_3_f;
   assign int_h2c_intr_3_h2c_2 = h2c_intr_3_h2c_2_f;
   assign int_h2c_intr_3_h2c_1 = h2c_intr_3_h2c_1_f;
   assign int_h2c_intr_3_h2c_0 = h2c_intr_3_h2c_0_f;
   assign int_c2h_intr_status_0_c2h_31 = c2h_intr_status_0_c2h_31_f;
   assign int_c2h_intr_status_0_c2h_30 = c2h_intr_status_0_c2h_30_f;
   assign int_c2h_intr_status_0_c2h_29 = c2h_intr_status_0_c2h_29_f;
   assign int_c2h_intr_status_0_c2h_28 = c2h_intr_status_0_c2h_28_f;
   assign int_c2h_intr_status_0_c2h_27 = c2h_intr_status_0_c2h_27_f;
   assign int_c2h_intr_status_0_c2h_26 = c2h_intr_status_0_c2h_26_f;
   assign int_c2h_intr_status_0_c2h_25 = c2h_intr_status_0_c2h_25_f;
   assign int_c2h_intr_status_0_c2h_24 = c2h_intr_status_0_c2h_24_f;
   assign int_c2h_intr_status_0_c2h_23 = c2h_intr_status_0_c2h_23_f;
   assign int_c2h_intr_status_0_c2h_22 = c2h_intr_status_0_c2h_22_f;
   assign int_c2h_intr_status_0_c2h_21 = c2h_intr_status_0_c2h_21_f;
   assign int_c2h_intr_status_0_c2h_20 = c2h_intr_status_0_c2h_20_f;
   assign int_c2h_intr_status_0_c2h_19 = c2h_intr_status_0_c2h_19_f;
   assign int_c2h_intr_status_0_c2h_18 = c2h_intr_status_0_c2h_18_f;
   assign int_c2h_intr_status_0_c2h_17 = c2h_intr_status_0_c2h_17_f;
   assign int_c2h_intr_status_0_c2h_16 = c2h_intr_status_0_c2h_16_f;
   assign int_c2h_intr_status_0_c2h_15 = c2h_intr_status_0_c2h_15_f;
   assign int_c2h_intr_status_0_c2h_14 = c2h_intr_status_0_c2h_14_f;
   assign int_c2h_intr_status_0_c2h_13 = c2h_intr_status_0_c2h_13_f;
   assign int_c2h_intr_status_0_c2h_12 = c2h_intr_status_0_c2h_12_f;
   assign int_c2h_intr_status_0_c2h_11 = c2h_intr_status_0_c2h_11_f;
   assign int_c2h_intr_status_0_c2h_10 = c2h_intr_status_0_c2h_10_f;
   assign int_c2h_intr_status_0_c2h_9 = c2h_intr_status_0_c2h_9_f;
   assign int_c2h_intr_status_0_c2h_8 = c2h_intr_status_0_c2h_8_f;
   assign int_c2h_intr_status_0_c2h_7 = c2h_intr_status_0_c2h_7_f;
   assign int_c2h_intr_status_0_c2h_6 = c2h_intr_status_0_c2h_6_f;
   assign int_c2h_intr_status_0_c2h_5 = c2h_intr_status_0_c2h_5_f;
   assign int_c2h_intr_status_0_c2h_4 = c2h_intr_status_0_c2h_4_f;
   assign int_c2h_intr_status_0_c2h_3 = c2h_intr_status_0_c2h_3_f;
   assign int_c2h_intr_status_0_c2h_2 = c2h_intr_status_0_c2h_2_f;
   assign int_c2h_intr_status_0_c2h_1 = c2h_intr_status_0_c2h_1_f;
   assign int_c2h_intr_status_0_c2h_0 = c2h_intr_status_0_c2h_0_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_31 = intr_c2h_toggle_status_0_t_c2h_31_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_30 = intr_c2h_toggle_status_0_t_c2h_30_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_29 = intr_c2h_toggle_status_0_t_c2h_29_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_28 = intr_c2h_toggle_status_0_t_c2h_28_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_27 = intr_c2h_toggle_status_0_t_c2h_27_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_26 = intr_c2h_toggle_status_0_t_c2h_26_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_25 = intr_c2h_toggle_status_0_t_c2h_25_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_24 = intr_c2h_toggle_status_0_t_c2h_24_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_23 = intr_c2h_toggle_status_0_t_c2h_23_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_22 = intr_c2h_toggle_status_0_t_c2h_22_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_21 = intr_c2h_toggle_status_0_t_c2h_21_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_20 = intr_c2h_toggle_status_0_t_c2h_20_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_19 = intr_c2h_toggle_status_0_t_c2h_19_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_18 = intr_c2h_toggle_status_0_t_c2h_18_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_17 = intr_c2h_toggle_status_0_t_c2h_17_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_16 = intr_c2h_toggle_status_0_t_c2h_16_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_15 = intr_c2h_toggle_status_0_t_c2h_15_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_14 = intr_c2h_toggle_status_0_t_c2h_14_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_13 = intr_c2h_toggle_status_0_t_c2h_13_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_12 = intr_c2h_toggle_status_0_t_c2h_12_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_11 = intr_c2h_toggle_status_0_t_c2h_11_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_10 = intr_c2h_toggle_status_0_t_c2h_10_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_9 = intr_c2h_toggle_status_0_t_c2h_9_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_8 = intr_c2h_toggle_status_0_t_c2h_8_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_7 = intr_c2h_toggle_status_0_t_c2h_7_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_6 = intr_c2h_toggle_status_0_t_c2h_6_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_5 = intr_c2h_toggle_status_0_t_c2h_5_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_4 = intr_c2h_toggle_status_0_t_c2h_4_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_3 = intr_c2h_toggle_status_0_t_c2h_3_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_2 = intr_c2h_toggle_status_0_t_c2h_2_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_1 = intr_c2h_toggle_status_0_t_c2h_1_f;
   assign int_intr_c2h_toggle_status_0_t_c2h_0 = intr_c2h_toggle_status_0_t_c2h_0_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_31 = intr_c2h_toggle_clear_0_clr_t_c2h_31_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_30 = intr_c2h_toggle_clear_0_clr_t_c2h_30_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_29 = intr_c2h_toggle_clear_0_clr_t_c2h_29_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_28 = intr_c2h_toggle_clear_0_clr_t_c2h_28_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_27 = intr_c2h_toggle_clear_0_clr_t_c2h_27_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_26 = intr_c2h_toggle_clear_0_clr_t_c2h_26_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_25 = intr_c2h_toggle_clear_0_clr_t_c2h_25_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_24 = intr_c2h_toggle_clear_0_clr_t_c2h_24_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_23 = intr_c2h_toggle_clear_0_clr_t_c2h_23_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_22 = intr_c2h_toggle_clear_0_clr_t_c2h_22_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_21 = intr_c2h_toggle_clear_0_clr_t_c2h_21_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_20 = intr_c2h_toggle_clear_0_clr_t_c2h_20_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_19 = intr_c2h_toggle_clear_0_clr_t_c2h_19_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_18 = intr_c2h_toggle_clear_0_clr_t_c2h_18_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_17 = intr_c2h_toggle_clear_0_clr_t_c2h_17_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_16 = intr_c2h_toggle_clear_0_clr_t_c2h_16_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_15 = intr_c2h_toggle_clear_0_clr_t_c2h_15_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_14 = intr_c2h_toggle_clear_0_clr_t_c2h_14_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_13 = intr_c2h_toggle_clear_0_clr_t_c2h_13_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_12 = intr_c2h_toggle_clear_0_clr_t_c2h_12_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_11 = intr_c2h_toggle_clear_0_clr_t_c2h_11_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_10 = intr_c2h_toggle_clear_0_clr_t_c2h_10_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_9 = intr_c2h_toggle_clear_0_clr_t_c2h_9_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_8 = intr_c2h_toggle_clear_0_clr_t_c2h_8_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_7 = intr_c2h_toggle_clear_0_clr_t_c2h_7_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_6 = intr_c2h_toggle_clear_0_clr_t_c2h_6_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_5 = intr_c2h_toggle_clear_0_clr_t_c2h_5_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_4 = intr_c2h_toggle_clear_0_clr_t_c2h_4_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_3 = intr_c2h_toggle_clear_0_clr_t_c2h_3_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_2 = intr_c2h_toggle_clear_0_clr_t_c2h_2_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_1 = intr_c2h_toggle_clear_0_clr_t_c2h_1_f;
   assign int_intr_c2h_toggle_clear_0_clr_t_c2h_0 = intr_c2h_toggle_clear_0_clr_t_c2h_0_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_31 = intr_c2h_toggle_enable_0_en_t_c2h_31_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_30 = intr_c2h_toggle_enable_0_en_t_c2h_30_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_29 = intr_c2h_toggle_enable_0_en_t_c2h_29_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_28 = intr_c2h_toggle_enable_0_en_t_c2h_28_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_27 = intr_c2h_toggle_enable_0_en_t_c2h_27_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_26 = intr_c2h_toggle_enable_0_en_t_c2h_26_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_25 = intr_c2h_toggle_enable_0_en_t_c2h_25_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_24 = intr_c2h_toggle_enable_0_en_t_c2h_24_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_23 = intr_c2h_toggle_enable_0_en_t_c2h_23_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_22 = intr_c2h_toggle_enable_0_en_t_c2h_22_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_21 = intr_c2h_toggle_enable_0_en_t_c2h_21_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_20 = intr_c2h_toggle_enable_0_en_t_c2h_20_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_19 = intr_c2h_toggle_enable_0_en_t_c2h_19_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_18 = intr_c2h_toggle_enable_0_en_t_c2h_18_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_17 = intr_c2h_toggle_enable_0_en_t_c2h_17_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_16 = intr_c2h_toggle_enable_0_en_t_c2h_16_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_15 = intr_c2h_toggle_enable_0_en_t_c2h_15_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_14 = intr_c2h_toggle_enable_0_en_t_c2h_14_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_13 = intr_c2h_toggle_enable_0_en_t_c2h_13_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_12 = intr_c2h_toggle_enable_0_en_t_c2h_12_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_11 = intr_c2h_toggle_enable_0_en_t_c2h_11_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_10 = intr_c2h_toggle_enable_0_en_t_c2h_10_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_9 = intr_c2h_toggle_enable_0_en_t_c2h_9_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_8 = intr_c2h_toggle_enable_0_en_t_c2h_8_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_7 = intr_c2h_toggle_enable_0_en_t_c2h_7_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_6 = intr_c2h_toggle_enable_0_en_t_c2h_6_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_5 = intr_c2h_toggle_enable_0_en_t_c2h_5_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_4 = intr_c2h_toggle_enable_0_en_t_c2h_4_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_3 = intr_c2h_toggle_enable_0_en_t_c2h_3_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_2 = intr_c2h_toggle_enable_0_en_t_c2h_2_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_1 = intr_c2h_toggle_enable_0_en_t_c2h_1_f;
   assign int_intr_c2h_toggle_enable_0_en_t_c2h_0 = intr_c2h_toggle_enable_0_en_t_c2h_0_f;
   assign int_c2h_intr_status_1_c2h_31 = c2h_intr_status_1_c2h_31_f;
   assign int_c2h_intr_status_1_c2h_30 = c2h_intr_status_1_c2h_30_f;
   assign int_c2h_intr_status_1_c2h_29 = c2h_intr_status_1_c2h_29_f;
   assign int_c2h_intr_status_1_c2h_28 = c2h_intr_status_1_c2h_28_f;
   assign int_c2h_intr_status_1_c2h_27 = c2h_intr_status_1_c2h_27_f;
   assign int_c2h_intr_status_1_c2h_26 = c2h_intr_status_1_c2h_26_f;
   assign int_c2h_intr_status_1_c2h_25 = c2h_intr_status_1_c2h_25_f;
   assign int_c2h_intr_status_1_c2h_24 = c2h_intr_status_1_c2h_24_f;
   assign int_c2h_intr_status_1_c2h_23 = c2h_intr_status_1_c2h_23_f;
   assign int_c2h_intr_status_1_c2h_22 = c2h_intr_status_1_c2h_22_f;
   assign int_c2h_intr_status_1_c2h_21 = c2h_intr_status_1_c2h_21_f;
   assign int_c2h_intr_status_1_c2h_20 = c2h_intr_status_1_c2h_20_f;
   assign int_c2h_intr_status_1_c2h_19 = c2h_intr_status_1_c2h_19_f;
   assign int_c2h_intr_status_1_c2h_18 = c2h_intr_status_1_c2h_18_f;
   assign int_c2h_intr_status_1_c2h_17 = c2h_intr_status_1_c2h_17_f;
   assign int_c2h_intr_status_1_c2h_16 = c2h_intr_status_1_c2h_16_f;
   assign int_c2h_intr_status_1_c2h_15 = c2h_intr_status_1_c2h_15_f;
   assign int_c2h_intr_status_1_c2h_14 = c2h_intr_status_1_c2h_14_f;
   assign int_c2h_intr_status_1_c2h_13 = c2h_intr_status_1_c2h_13_f;
   assign int_c2h_intr_status_1_c2h_12 = c2h_intr_status_1_c2h_12_f;
   assign int_c2h_intr_status_1_c2h_11 = c2h_intr_status_1_c2h_11_f;
   assign int_c2h_intr_status_1_c2h_10 = c2h_intr_status_1_c2h_10_f;
   assign int_c2h_intr_status_1_c2h_9 = c2h_intr_status_1_c2h_9_f;
   assign int_c2h_intr_status_1_c2h_8 = c2h_intr_status_1_c2h_8_f;
   assign int_c2h_intr_status_1_c2h_7 = c2h_intr_status_1_c2h_7_f;
   assign int_c2h_intr_status_1_c2h_6 = c2h_intr_status_1_c2h_6_f;
   assign int_c2h_intr_status_1_c2h_5 = c2h_intr_status_1_c2h_5_f;
   assign int_c2h_intr_status_1_c2h_4 = c2h_intr_status_1_c2h_4_f;
   assign int_c2h_intr_status_1_c2h_3 = c2h_intr_status_1_c2h_3_f;
   assign int_c2h_intr_status_1_c2h_2 = c2h_intr_status_1_c2h_2_f;
   assign int_c2h_intr_status_1_c2h_1 = c2h_intr_status_1_c2h_1_f;
   assign int_c2h_intr_status_1_c2h_0 = c2h_intr_status_1_c2h_0_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_31 = intr_c2h_toggle_status_1_t_c2h_31_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_30 = intr_c2h_toggle_status_1_t_c2h_30_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_29 = intr_c2h_toggle_status_1_t_c2h_29_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_28 = intr_c2h_toggle_status_1_t_c2h_28_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_27 = intr_c2h_toggle_status_1_t_c2h_27_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_26 = intr_c2h_toggle_status_1_t_c2h_26_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_25 = intr_c2h_toggle_status_1_t_c2h_25_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_24 = intr_c2h_toggle_status_1_t_c2h_24_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_23 = intr_c2h_toggle_status_1_t_c2h_23_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_22 = intr_c2h_toggle_status_1_t_c2h_22_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_21 = intr_c2h_toggle_status_1_t_c2h_21_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_20 = intr_c2h_toggle_status_1_t_c2h_20_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_19 = intr_c2h_toggle_status_1_t_c2h_19_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_18 = intr_c2h_toggle_status_1_t_c2h_18_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_17 = intr_c2h_toggle_status_1_t_c2h_17_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_16 = intr_c2h_toggle_status_1_t_c2h_16_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_15 = intr_c2h_toggle_status_1_t_c2h_15_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_14 = intr_c2h_toggle_status_1_t_c2h_14_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_13 = intr_c2h_toggle_status_1_t_c2h_13_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_12 = intr_c2h_toggle_status_1_t_c2h_12_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_11 = intr_c2h_toggle_status_1_t_c2h_11_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_10 = intr_c2h_toggle_status_1_t_c2h_10_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_9 = intr_c2h_toggle_status_1_t_c2h_9_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_8 = intr_c2h_toggle_status_1_t_c2h_8_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_7 = intr_c2h_toggle_status_1_t_c2h_7_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_6 = intr_c2h_toggle_status_1_t_c2h_6_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_5 = intr_c2h_toggle_status_1_t_c2h_5_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_4 = intr_c2h_toggle_status_1_t_c2h_4_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_3 = intr_c2h_toggle_status_1_t_c2h_3_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_2 = intr_c2h_toggle_status_1_t_c2h_2_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_1 = intr_c2h_toggle_status_1_t_c2h_1_f;
   assign int_intr_c2h_toggle_status_1_t_c2h_0 = intr_c2h_toggle_status_1_t_c2h_0_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_31 = intr_c2h_toggle_clear_1_clr_t_c2h_31_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_30 = intr_c2h_toggle_clear_1_clr_t_c2h_30_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_29 = intr_c2h_toggle_clear_1_clr_t_c2h_29_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_28 = intr_c2h_toggle_clear_1_clr_t_c2h_28_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_27 = intr_c2h_toggle_clear_1_clr_t_c2h_27_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_26 = intr_c2h_toggle_clear_1_clr_t_c2h_26_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_25 = intr_c2h_toggle_clear_1_clr_t_c2h_25_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_24 = intr_c2h_toggle_clear_1_clr_t_c2h_24_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_23 = intr_c2h_toggle_clear_1_clr_t_c2h_23_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_22 = intr_c2h_toggle_clear_1_clr_t_c2h_22_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_21 = intr_c2h_toggle_clear_1_clr_t_c2h_21_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_20 = intr_c2h_toggle_clear_1_clr_t_c2h_20_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_19 = intr_c2h_toggle_clear_1_clr_t_c2h_19_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_18 = intr_c2h_toggle_clear_1_clr_t_c2h_18_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_17 = intr_c2h_toggle_clear_1_clr_t_c2h_17_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_16 = intr_c2h_toggle_clear_1_clr_t_c2h_16_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_15 = intr_c2h_toggle_clear_1_clr_t_c2h_15_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_14 = intr_c2h_toggle_clear_1_clr_t_c2h_14_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_13 = intr_c2h_toggle_clear_1_clr_t_c2h_13_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_12 = intr_c2h_toggle_clear_1_clr_t_c2h_12_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_11 = intr_c2h_toggle_clear_1_clr_t_c2h_11_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_10 = intr_c2h_toggle_clear_1_clr_t_c2h_10_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_9 = intr_c2h_toggle_clear_1_clr_t_c2h_9_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_8 = intr_c2h_toggle_clear_1_clr_t_c2h_8_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_7 = intr_c2h_toggle_clear_1_clr_t_c2h_7_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_6 = intr_c2h_toggle_clear_1_clr_t_c2h_6_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_5 = intr_c2h_toggle_clear_1_clr_t_c2h_5_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_4 = intr_c2h_toggle_clear_1_clr_t_c2h_4_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_3 = intr_c2h_toggle_clear_1_clr_t_c2h_3_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_2 = intr_c2h_toggle_clear_1_clr_t_c2h_2_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_1 = intr_c2h_toggle_clear_1_clr_t_c2h_1_f;
   assign int_intr_c2h_toggle_clear_1_clr_t_c2h_0 = intr_c2h_toggle_clear_1_clr_t_c2h_0_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_31 = intr_c2h_toggle_enable_1_en_t_c2h_31_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_30 = intr_c2h_toggle_enable_1_en_t_c2h_30_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_29 = intr_c2h_toggle_enable_1_en_t_c2h_29_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_28 = intr_c2h_toggle_enable_1_en_t_c2h_28_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_27 = intr_c2h_toggle_enable_1_en_t_c2h_27_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_26 = intr_c2h_toggle_enable_1_en_t_c2h_26_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_25 = intr_c2h_toggle_enable_1_en_t_c2h_25_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_24 = intr_c2h_toggle_enable_1_en_t_c2h_24_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_23 = intr_c2h_toggle_enable_1_en_t_c2h_23_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_22 = intr_c2h_toggle_enable_1_en_t_c2h_22_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_21 = intr_c2h_toggle_enable_1_en_t_c2h_21_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_20 = intr_c2h_toggle_enable_1_en_t_c2h_20_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_19 = intr_c2h_toggle_enable_1_en_t_c2h_19_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_18 = intr_c2h_toggle_enable_1_en_t_c2h_18_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_17 = intr_c2h_toggle_enable_1_en_t_c2h_17_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_16 = intr_c2h_toggle_enable_1_en_t_c2h_16_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_15 = intr_c2h_toggle_enable_1_en_t_c2h_15_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_14 = intr_c2h_toggle_enable_1_en_t_c2h_14_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_13 = intr_c2h_toggle_enable_1_en_t_c2h_13_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_12 = intr_c2h_toggle_enable_1_en_t_c2h_12_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_11 = intr_c2h_toggle_enable_1_en_t_c2h_11_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_10 = intr_c2h_toggle_enable_1_en_t_c2h_10_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_9 = intr_c2h_toggle_enable_1_en_t_c2h_9_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_8 = intr_c2h_toggle_enable_1_en_t_c2h_8_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_7 = intr_c2h_toggle_enable_1_en_t_c2h_7_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_6 = intr_c2h_toggle_enable_1_en_t_c2h_6_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_5 = intr_c2h_toggle_enable_1_en_t_c2h_5_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_4 = intr_c2h_toggle_enable_1_en_t_c2h_4_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_3 = intr_c2h_toggle_enable_1_en_t_c2h_3_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_2 = intr_c2h_toggle_enable_1_en_t_c2h_2_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_1 = intr_c2h_toggle_enable_1_en_t_c2h_1_f;
   assign int_intr_c2h_toggle_enable_1_en_t_c2h_0 = intr_c2h_toggle_enable_1_en_t_c2h_0_f;
   assign int_c2h_gpio_0_gpio_31 = c2h_gpio_0_gpio_31_f;
   assign int_c2h_gpio_0_gpio_30 = c2h_gpio_0_gpio_30_f;
   assign int_c2h_gpio_0_gpio_29 = c2h_gpio_0_gpio_29_f;
   assign int_c2h_gpio_0_gpio_28 = c2h_gpio_0_gpio_28_f;
   assign int_c2h_gpio_0_gpio_27 = c2h_gpio_0_gpio_27_f;
   assign int_c2h_gpio_0_gpio_26 = c2h_gpio_0_gpio_26_f;
   assign int_c2h_gpio_0_gpio_25 = c2h_gpio_0_gpio_25_f;
   assign int_c2h_gpio_0_gpio_24 = c2h_gpio_0_gpio_24_f;
   assign int_c2h_gpio_0_gpio_23 = c2h_gpio_0_gpio_23_f;
   assign int_c2h_gpio_0_gpio_22 = c2h_gpio_0_gpio_22_f;
   assign int_c2h_gpio_0_gpio_21 = c2h_gpio_0_gpio_21_f;
   assign int_c2h_gpio_0_gpio_20 = c2h_gpio_0_gpio_20_f;
   assign int_c2h_gpio_0_gpio_19 = c2h_gpio_0_gpio_19_f;
   assign int_c2h_gpio_0_gpio_18 = c2h_gpio_0_gpio_18_f;
   assign int_c2h_gpio_0_gpio_17 = c2h_gpio_0_gpio_17_f;
   assign int_c2h_gpio_0_gpio_16 = c2h_gpio_0_gpio_16_f;
   assign int_c2h_gpio_0_gpio_15 = c2h_gpio_0_gpio_15_f;
   assign int_c2h_gpio_0_gpio_14 = c2h_gpio_0_gpio_14_f;
   assign int_c2h_gpio_0_gpio_13 = c2h_gpio_0_gpio_13_f;
   assign int_c2h_gpio_0_gpio_12 = c2h_gpio_0_gpio_12_f;
   assign int_c2h_gpio_0_gpio_11 = c2h_gpio_0_gpio_11_f;
   assign int_c2h_gpio_0_gpio_10 = c2h_gpio_0_gpio_10_f;
   assign int_c2h_gpio_0_gpio_9 = c2h_gpio_0_gpio_9_f;
   assign int_c2h_gpio_0_gpio_8 = c2h_gpio_0_gpio_8_f;
   assign int_c2h_gpio_0_gpio_7 = c2h_gpio_0_gpio_7_f;
   assign int_c2h_gpio_0_gpio_6 = c2h_gpio_0_gpio_6_f;
   assign int_c2h_gpio_0_gpio_5 = c2h_gpio_0_gpio_5_f;
   assign int_c2h_gpio_0_gpio_4 = c2h_gpio_0_gpio_4_f;
   assign int_c2h_gpio_0_gpio_3 = c2h_gpio_0_gpio_3_f;
   assign int_c2h_gpio_0_gpio_2 = c2h_gpio_0_gpio_2_f;
   assign int_c2h_gpio_0_gpio_1 = c2h_gpio_0_gpio_1_f;
   assign int_c2h_gpio_0_gpio_0 = c2h_gpio_0_gpio_0_f;
   assign int_c2h_gpio_1_gpio_31 = c2h_gpio_1_gpio_31_f;
   assign int_c2h_gpio_1_gpio_30 = c2h_gpio_1_gpio_30_f;
   assign int_c2h_gpio_1_gpio_29 = c2h_gpio_1_gpio_29_f;
   assign int_c2h_gpio_1_gpio_28 = c2h_gpio_1_gpio_28_f;
   assign int_c2h_gpio_1_gpio_27 = c2h_gpio_1_gpio_27_f;
   assign int_c2h_gpio_1_gpio_26 = c2h_gpio_1_gpio_26_f;
   assign int_c2h_gpio_1_gpio_25 = c2h_gpio_1_gpio_25_f;
   assign int_c2h_gpio_1_gpio_24 = c2h_gpio_1_gpio_24_f;
   assign int_c2h_gpio_1_gpio_23 = c2h_gpio_1_gpio_23_f;
   assign int_c2h_gpio_1_gpio_22 = c2h_gpio_1_gpio_22_f;
   assign int_c2h_gpio_1_gpio_21 = c2h_gpio_1_gpio_21_f;
   assign int_c2h_gpio_1_gpio_20 = c2h_gpio_1_gpio_20_f;
   assign int_c2h_gpio_1_gpio_19 = c2h_gpio_1_gpio_19_f;
   assign int_c2h_gpio_1_gpio_18 = c2h_gpio_1_gpio_18_f;
   assign int_c2h_gpio_1_gpio_17 = c2h_gpio_1_gpio_17_f;
   assign int_c2h_gpio_1_gpio_16 = c2h_gpio_1_gpio_16_f;
   assign int_c2h_gpio_1_gpio_15 = c2h_gpio_1_gpio_15_f;
   assign int_c2h_gpio_1_gpio_14 = c2h_gpio_1_gpio_14_f;
   assign int_c2h_gpio_1_gpio_13 = c2h_gpio_1_gpio_13_f;
   assign int_c2h_gpio_1_gpio_12 = c2h_gpio_1_gpio_12_f;
   assign int_c2h_gpio_1_gpio_11 = c2h_gpio_1_gpio_11_f;
   assign int_c2h_gpio_1_gpio_10 = c2h_gpio_1_gpio_10_f;
   assign int_c2h_gpio_1_gpio_9 = c2h_gpio_1_gpio_9_f;
   assign int_c2h_gpio_1_gpio_8 = c2h_gpio_1_gpio_8_f;
   assign int_c2h_gpio_1_gpio_7 = c2h_gpio_1_gpio_7_f;
   assign int_c2h_gpio_1_gpio_6 = c2h_gpio_1_gpio_6_f;
   assign int_c2h_gpio_1_gpio_5 = c2h_gpio_1_gpio_5_f;
   assign int_c2h_gpio_1_gpio_4 = c2h_gpio_1_gpio_4_f;
   assign int_c2h_gpio_1_gpio_3 = c2h_gpio_1_gpio_3_f;
   assign int_c2h_gpio_1_gpio_2 = c2h_gpio_1_gpio_2_f;
   assign int_c2h_gpio_1_gpio_1 = c2h_gpio_1_gpio_1_f;
   assign int_c2h_gpio_1_gpio_0 = c2h_gpio_1_gpio_0_f;
   assign int_c2h_gpio_2_gpio_31 = c2h_gpio_2_gpio_31_f;
   assign int_c2h_gpio_2_gpio_30 = c2h_gpio_2_gpio_30_f;
   assign int_c2h_gpio_2_gpio_29 = c2h_gpio_2_gpio_29_f;
   assign int_c2h_gpio_2_gpio_28 = c2h_gpio_2_gpio_28_f;
   assign int_c2h_gpio_2_gpio_27 = c2h_gpio_2_gpio_27_f;
   assign int_c2h_gpio_2_gpio_26 = c2h_gpio_2_gpio_26_f;
   assign int_c2h_gpio_2_gpio_25 = c2h_gpio_2_gpio_25_f;
   assign int_c2h_gpio_2_gpio_24 = c2h_gpio_2_gpio_24_f;
   assign int_c2h_gpio_2_gpio_23 = c2h_gpio_2_gpio_23_f;
   assign int_c2h_gpio_2_gpio_22 = c2h_gpio_2_gpio_22_f;
   assign int_c2h_gpio_2_gpio_21 = c2h_gpio_2_gpio_21_f;
   assign int_c2h_gpio_2_gpio_20 = c2h_gpio_2_gpio_20_f;
   assign int_c2h_gpio_2_gpio_19 = c2h_gpio_2_gpio_19_f;
   assign int_c2h_gpio_2_gpio_18 = c2h_gpio_2_gpio_18_f;
   assign int_c2h_gpio_2_gpio_17 = c2h_gpio_2_gpio_17_f;
   assign int_c2h_gpio_2_gpio_16 = c2h_gpio_2_gpio_16_f;
   assign int_c2h_gpio_2_gpio_15 = c2h_gpio_2_gpio_15_f;
   assign int_c2h_gpio_2_gpio_14 = c2h_gpio_2_gpio_14_f;
   assign int_c2h_gpio_2_gpio_13 = c2h_gpio_2_gpio_13_f;
   assign int_c2h_gpio_2_gpio_12 = c2h_gpio_2_gpio_12_f;
   assign int_c2h_gpio_2_gpio_11 = c2h_gpio_2_gpio_11_f;
   assign int_c2h_gpio_2_gpio_10 = c2h_gpio_2_gpio_10_f;
   assign int_c2h_gpio_2_gpio_9 = c2h_gpio_2_gpio_9_f;
   assign int_c2h_gpio_2_gpio_8 = c2h_gpio_2_gpio_8_f;
   assign int_c2h_gpio_2_gpio_7 = c2h_gpio_2_gpio_7_f;
   assign int_c2h_gpio_2_gpio_6 = c2h_gpio_2_gpio_6_f;
   assign int_c2h_gpio_2_gpio_5 = c2h_gpio_2_gpio_5_f;
   assign int_c2h_gpio_2_gpio_4 = c2h_gpio_2_gpio_4_f;
   assign int_c2h_gpio_2_gpio_3 = c2h_gpio_2_gpio_3_f;
   assign int_c2h_gpio_2_gpio_2 = c2h_gpio_2_gpio_2_f;
   assign int_c2h_gpio_2_gpio_1 = c2h_gpio_2_gpio_1_f;
   assign int_c2h_gpio_2_gpio_0 = c2h_gpio_2_gpio_0_f;
   assign int_c2h_gpio_3_gpio_31 = c2h_gpio_3_gpio_31_f;
   assign int_c2h_gpio_3_gpio_30 = c2h_gpio_3_gpio_30_f;
   assign int_c2h_gpio_3_gpio_29 = c2h_gpio_3_gpio_29_f;
   assign int_c2h_gpio_3_gpio_28 = c2h_gpio_3_gpio_28_f;
   assign int_c2h_gpio_3_gpio_27 = c2h_gpio_3_gpio_27_f;
   assign int_c2h_gpio_3_gpio_26 = c2h_gpio_3_gpio_26_f;
   assign int_c2h_gpio_3_gpio_25 = c2h_gpio_3_gpio_25_f;
   assign int_c2h_gpio_3_gpio_24 = c2h_gpio_3_gpio_24_f;
   assign int_c2h_gpio_3_gpio_23 = c2h_gpio_3_gpio_23_f;
   assign int_c2h_gpio_3_gpio_22 = c2h_gpio_3_gpio_22_f;
   assign int_c2h_gpio_3_gpio_21 = c2h_gpio_3_gpio_21_f;
   assign int_c2h_gpio_3_gpio_20 = c2h_gpio_3_gpio_20_f;
   assign int_c2h_gpio_3_gpio_19 = c2h_gpio_3_gpio_19_f;
   assign int_c2h_gpio_3_gpio_18 = c2h_gpio_3_gpio_18_f;
   assign int_c2h_gpio_3_gpio_17 = c2h_gpio_3_gpio_17_f;
   assign int_c2h_gpio_3_gpio_16 = c2h_gpio_3_gpio_16_f;
   assign int_c2h_gpio_3_gpio_15 = c2h_gpio_3_gpio_15_f;
   assign int_c2h_gpio_3_gpio_14 = c2h_gpio_3_gpio_14_f;
   assign int_c2h_gpio_3_gpio_13 = c2h_gpio_3_gpio_13_f;
   assign int_c2h_gpio_3_gpio_12 = c2h_gpio_3_gpio_12_f;
   assign int_c2h_gpio_3_gpio_11 = c2h_gpio_3_gpio_11_f;
   assign int_c2h_gpio_3_gpio_10 = c2h_gpio_3_gpio_10_f;
   assign int_c2h_gpio_3_gpio_9 = c2h_gpio_3_gpio_9_f;
   assign int_c2h_gpio_3_gpio_8 = c2h_gpio_3_gpio_8_f;
   assign int_c2h_gpio_3_gpio_7 = c2h_gpio_3_gpio_7_f;
   assign int_c2h_gpio_3_gpio_6 = c2h_gpio_3_gpio_6_f;
   assign int_c2h_gpio_3_gpio_5 = c2h_gpio_3_gpio_5_f;
   assign int_c2h_gpio_3_gpio_4 = c2h_gpio_3_gpio_4_f;
   assign int_c2h_gpio_3_gpio_3 = c2h_gpio_3_gpio_3_f;
   assign int_c2h_gpio_3_gpio_2 = c2h_gpio_3_gpio_2_f;
   assign int_c2h_gpio_3_gpio_1 = c2h_gpio_3_gpio_1_f;
   assign int_c2h_gpio_3_gpio_0 = c2h_gpio_3_gpio_0_f;
   assign int_c2h_gpio_4_gpio_31 = c2h_gpio_4_gpio_31_f;
   assign int_c2h_gpio_4_gpio_30 = c2h_gpio_4_gpio_30_f;
   assign int_c2h_gpio_4_gpio_29 = c2h_gpio_4_gpio_29_f;
   assign int_c2h_gpio_4_gpio_28 = c2h_gpio_4_gpio_28_f;
   assign int_c2h_gpio_4_gpio_27 = c2h_gpio_4_gpio_27_f;
   assign int_c2h_gpio_4_gpio_26 = c2h_gpio_4_gpio_26_f;
   assign int_c2h_gpio_4_gpio_25 = c2h_gpio_4_gpio_25_f;
   assign int_c2h_gpio_4_gpio_24 = c2h_gpio_4_gpio_24_f;
   assign int_c2h_gpio_4_gpio_23 = c2h_gpio_4_gpio_23_f;
   assign int_c2h_gpio_4_gpio_22 = c2h_gpio_4_gpio_22_f;
   assign int_c2h_gpio_4_gpio_21 = c2h_gpio_4_gpio_21_f;
   assign int_c2h_gpio_4_gpio_20 = c2h_gpio_4_gpio_20_f;
   assign int_c2h_gpio_4_gpio_19 = c2h_gpio_4_gpio_19_f;
   assign int_c2h_gpio_4_gpio_18 = c2h_gpio_4_gpio_18_f;
   assign int_c2h_gpio_4_gpio_17 = c2h_gpio_4_gpio_17_f;
   assign int_c2h_gpio_4_gpio_16 = c2h_gpio_4_gpio_16_f;
   assign int_c2h_gpio_4_gpio_15 = c2h_gpio_4_gpio_15_f;
   assign int_c2h_gpio_4_gpio_14 = c2h_gpio_4_gpio_14_f;
   assign int_c2h_gpio_4_gpio_13 = c2h_gpio_4_gpio_13_f;
   assign int_c2h_gpio_4_gpio_12 = c2h_gpio_4_gpio_12_f;
   assign int_c2h_gpio_4_gpio_11 = c2h_gpio_4_gpio_11_f;
   assign int_c2h_gpio_4_gpio_10 = c2h_gpio_4_gpio_10_f;
   assign int_c2h_gpio_4_gpio_9 = c2h_gpio_4_gpio_9_f;
   assign int_c2h_gpio_4_gpio_8 = c2h_gpio_4_gpio_8_f;
   assign int_c2h_gpio_4_gpio_7 = c2h_gpio_4_gpio_7_f;
   assign int_c2h_gpio_4_gpio_6 = c2h_gpio_4_gpio_6_f;
   assign int_c2h_gpio_4_gpio_5 = c2h_gpio_4_gpio_5_f;
   assign int_c2h_gpio_4_gpio_4 = c2h_gpio_4_gpio_4_f;
   assign int_c2h_gpio_4_gpio_3 = c2h_gpio_4_gpio_3_f;
   assign int_c2h_gpio_4_gpio_2 = c2h_gpio_4_gpio_2_f;
   assign int_c2h_gpio_4_gpio_1 = c2h_gpio_4_gpio_1_f;
   assign int_c2h_gpio_4_gpio_0 = c2h_gpio_4_gpio_0_f;
   assign int_c2h_gpio_5_gpio_31 = c2h_gpio_5_gpio_31_f;
   assign int_c2h_gpio_5_gpio_30 = c2h_gpio_5_gpio_30_f;
   assign int_c2h_gpio_5_gpio_29 = c2h_gpio_5_gpio_29_f;
   assign int_c2h_gpio_5_gpio_28 = c2h_gpio_5_gpio_28_f;
   assign int_c2h_gpio_5_gpio_27 = c2h_gpio_5_gpio_27_f;
   assign int_c2h_gpio_5_gpio_26 = c2h_gpio_5_gpio_26_f;
   assign int_c2h_gpio_5_gpio_25 = c2h_gpio_5_gpio_25_f;
   assign int_c2h_gpio_5_gpio_24 = c2h_gpio_5_gpio_24_f;
   assign int_c2h_gpio_5_gpio_23 = c2h_gpio_5_gpio_23_f;
   assign int_c2h_gpio_5_gpio_22 = c2h_gpio_5_gpio_22_f;
   assign int_c2h_gpio_5_gpio_21 = c2h_gpio_5_gpio_21_f;
   assign int_c2h_gpio_5_gpio_20 = c2h_gpio_5_gpio_20_f;
   assign int_c2h_gpio_5_gpio_19 = c2h_gpio_5_gpio_19_f;
   assign int_c2h_gpio_5_gpio_18 = c2h_gpio_5_gpio_18_f;
   assign int_c2h_gpio_5_gpio_17 = c2h_gpio_5_gpio_17_f;
   assign int_c2h_gpio_5_gpio_16 = c2h_gpio_5_gpio_16_f;
   assign int_c2h_gpio_5_gpio_15 = c2h_gpio_5_gpio_15_f;
   assign int_c2h_gpio_5_gpio_14 = c2h_gpio_5_gpio_14_f;
   assign int_c2h_gpio_5_gpio_13 = c2h_gpio_5_gpio_13_f;
   assign int_c2h_gpio_5_gpio_12 = c2h_gpio_5_gpio_12_f;
   assign int_c2h_gpio_5_gpio_11 = c2h_gpio_5_gpio_11_f;
   assign int_c2h_gpio_5_gpio_10 = c2h_gpio_5_gpio_10_f;
   assign int_c2h_gpio_5_gpio_9 = c2h_gpio_5_gpio_9_f;
   assign int_c2h_gpio_5_gpio_8 = c2h_gpio_5_gpio_8_f;
   assign int_c2h_gpio_5_gpio_7 = c2h_gpio_5_gpio_7_f;
   assign int_c2h_gpio_5_gpio_6 = c2h_gpio_5_gpio_6_f;
   assign int_c2h_gpio_5_gpio_5 = c2h_gpio_5_gpio_5_f;
   assign int_c2h_gpio_5_gpio_4 = c2h_gpio_5_gpio_4_f;
   assign int_c2h_gpio_5_gpio_3 = c2h_gpio_5_gpio_3_f;
   assign int_c2h_gpio_5_gpio_2 = c2h_gpio_5_gpio_2_f;
   assign int_c2h_gpio_5_gpio_1 = c2h_gpio_5_gpio_1_f;
   assign int_c2h_gpio_5_gpio_0 = c2h_gpio_5_gpio_0_f;
   assign int_c2h_gpio_6_gpio_31 = c2h_gpio_6_gpio_31_f;
   assign int_c2h_gpio_6_gpio_30 = c2h_gpio_6_gpio_30_f;
   assign int_c2h_gpio_6_gpio_29 = c2h_gpio_6_gpio_29_f;
   assign int_c2h_gpio_6_gpio_28 = c2h_gpio_6_gpio_28_f;
   assign int_c2h_gpio_6_gpio_27 = c2h_gpio_6_gpio_27_f;
   assign int_c2h_gpio_6_gpio_26 = c2h_gpio_6_gpio_26_f;
   assign int_c2h_gpio_6_gpio_25 = c2h_gpio_6_gpio_25_f;
   assign int_c2h_gpio_6_gpio_24 = c2h_gpio_6_gpio_24_f;
   assign int_c2h_gpio_6_gpio_23 = c2h_gpio_6_gpio_23_f;
   assign int_c2h_gpio_6_gpio_22 = c2h_gpio_6_gpio_22_f;
   assign int_c2h_gpio_6_gpio_21 = c2h_gpio_6_gpio_21_f;
   assign int_c2h_gpio_6_gpio_20 = c2h_gpio_6_gpio_20_f;
   assign int_c2h_gpio_6_gpio_19 = c2h_gpio_6_gpio_19_f;
   assign int_c2h_gpio_6_gpio_18 = c2h_gpio_6_gpio_18_f;
   assign int_c2h_gpio_6_gpio_17 = c2h_gpio_6_gpio_17_f;
   assign int_c2h_gpio_6_gpio_16 = c2h_gpio_6_gpio_16_f;
   assign int_c2h_gpio_6_gpio_15 = c2h_gpio_6_gpio_15_f;
   assign int_c2h_gpio_6_gpio_14 = c2h_gpio_6_gpio_14_f;
   assign int_c2h_gpio_6_gpio_13 = c2h_gpio_6_gpio_13_f;
   assign int_c2h_gpio_6_gpio_12 = c2h_gpio_6_gpio_12_f;
   assign int_c2h_gpio_6_gpio_11 = c2h_gpio_6_gpio_11_f;
   assign int_c2h_gpio_6_gpio_10 = c2h_gpio_6_gpio_10_f;
   assign int_c2h_gpio_6_gpio_9 = c2h_gpio_6_gpio_9_f;
   assign int_c2h_gpio_6_gpio_8 = c2h_gpio_6_gpio_8_f;
   assign int_c2h_gpio_6_gpio_7 = c2h_gpio_6_gpio_7_f;
   assign int_c2h_gpio_6_gpio_6 = c2h_gpio_6_gpio_6_f;
   assign int_c2h_gpio_6_gpio_5 = c2h_gpio_6_gpio_5_f;
   assign int_c2h_gpio_6_gpio_4 = c2h_gpio_6_gpio_4_f;
   assign int_c2h_gpio_6_gpio_3 = c2h_gpio_6_gpio_3_f;
   assign int_c2h_gpio_6_gpio_2 = c2h_gpio_6_gpio_2_f;
   assign int_c2h_gpio_6_gpio_1 = c2h_gpio_6_gpio_1_f;
   assign int_c2h_gpio_6_gpio_0 = c2h_gpio_6_gpio_0_f;
   assign int_c2h_gpio_7_gpio_31 = c2h_gpio_7_gpio_31_f;
   assign int_c2h_gpio_7_gpio_30 = c2h_gpio_7_gpio_30_f;
   assign int_c2h_gpio_7_gpio_29 = c2h_gpio_7_gpio_29_f;
   assign int_c2h_gpio_7_gpio_28 = c2h_gpio_7_gpio_28_f;
   assign int_c2h_gpio_7_gpio_27 = c2h_gpio_7_gpio_27_f;
   assign int_c2h_gpio_7_gpio_26 = c2h_gpio_7_gpio_26_f;
   assign int_c2h_gpio_7_gpio_25 = c2h_gpio_7_gpio_25_f;
   assign int_c2h_gpio_7_gpio_24 = c2h_gpio_7_gpio_24_f;
   assign int_c2h_gpio_7_gpio_23 = c2h_gpio_7_gpio_23_f;
   assign int_c2h_gpio_7_gpio_22 = c2h_gpio_7_gpio_22_f;
   assign int_c2h_gpio_7_gpio_21 = c2h_gpio_7_gpio_21_f;
   assign int_c2h_gpio_7_gpio_20 = c2h_gpio_7_gpio_20_f;
   assign int_c2h_gpio_7_gpio_19 = c2h_gpio_7_gpio_19_f;
   assign int_c2h_gpio_7_gpio_18 = c2h_gpio_7_gpio_18_f;
   assign int_c2h_gpio_7_gpio_17 = c2h_gpio_7_gpio_17_f;
   assign int_c2h_gpio_7_gpio_16 = c2h_gpio_7_gpio_16_f;
   assign int_c2h_gpio_7_gpio_15 = c2h_gpio_7_gpio_15_f;
   assign int_c2h_gpio_7_gpio_14 = c2h_gpio_7_gpio_14_f;
   assign int_c2h_gpio_7_gpio_13 = c2h_gpio_7_gpio_13_f;
   assign int_c2h_gpio_7_gpio_12 = c2h_gpio_7_gpio_12_f;
   assign int_c2h_gpio_7_gpio_11 = c2h_gpio_7_gpio_11_f;
   assign int_c2h_gpio_7_gpio_10 = c2h_gpio_7_gpio_10_f;
   assign int_c2h_gpio_7_gpio_9 = c2h_gpio_7_gpio_9_f;
   assign int_c2h_gpio_7_gpio_8 = c2h_gpio_7_gpio_8_f;
   assign int_c2h_gpio_7_gpio_7 = c2h_gpio_7_gpio_7_f;
   assign int_c2h_gpio_7_gpio_6 = c2h_gpio_7_gpio_6_f;
   assign int_c2h_gpio_7_gpio_5 = c2h_gpio_7_gpio_5_f;
   assign int_c2h_gpio_7_gpio_4 = c2h_gpio_7_gpio_4_f;
   assign int_c2h_gpio_7_gpio_3 = c2h_gpio_7_gpio_3_f;
   assign int_c2h_gpio_7_gpio_2 = c2h_gpio_7_gpio_2_f;
   assign int_c2h_gpio_7_gpio_1 = c2h_gpio_7_gpio_1_f;
   assign int_c2h_gpio_7_gpio_0 = c2h_gpio_7_gpio_0_f;
   assign int_c2h_gpio_8_gpio_31 = c2h_gpio_8_gpio_31_f;
   assign int_c2h_gpio_8_gpio_30 = c2h_gpio_8_gpio_30_f;
   assign int_c2h_gpio_8_gpio_29 = c2h_gpio_8_gpio_29_f;
   assign int_c2h_gpio_8_gpio_28 = c2h_gpio_8_gpio_28_f;
   assign int_c2h_gpio_8_gpio_27 = c2h_gpio_8_gpio_27_f;
   assign int_c2h_gpio_8_gpio_26 = c2h_gpio_8_gpio_26_f;
   assign int_c2h_gpio_8_gpio_25 = c2h_gpio_8_gpio_25_f;
   assign int_c2h_gpio_8_gpio_24 = c2h_gpio_8_gpio_24_f;
   assign int_c2h_gpio_8_gpio_23 = c2h_gpio_8_gpio_23_f;
   assign int_c2h_gpio_8_gpio_22 = c2h_gpio_8_gpio_22_f;
   assign int_c2h_gpio_8_gpio_21 = c2h_gpio_8_gpio_21_f;
   assign int_c2h_gpio_8_gpio_20 = c2h_gpio_8_gpio_20_f;
   assign int_c2h_gpio_8_gpio_19 = c2h_gpio_8_gpio_19_f;
   assign int_c2h_gpio_8_gpio_18 = c2h_gpio_8_gpio_18_f;
   assign int_c2h_gpio_8_gpio_17 = c2h_gpio_8_gpio_17_f;
   assign int_c2h_gpio_8_gpio_16 = c2h_gpio_8_gpio_16_f;
   assign int_c2h_gpio_8_gpio_15 = c2h_gpio_8_gpio_15_f;
   assign int_c2h_gpio_8_gpio_14 = c2h_gpio_8_gpio_14_f;
   assign int_c2h_gpio_8_gpio_13 = c2h_gpio_8_gpio_13_f;
   assign int_c2h_gpio_8_gpio_12 = c2h_gpio_8_gpio_12_f;
   assign int_c2h_gpio_8_gpio_11 = c2h_gpio_8_gpio_11_f;
   assign int_c2h_gpio_8_gpio_10 = c2h_gpio_8_gpio_10_f;
   assign int_c2h_gpio_8_gpio_9 = c2h_gpio_8_gpio_9_f;
   assign int_c2h_gpio_8_gpio_8 = c2h_gpio_8_gpio_8_f;
   assign int_c2h_gpio_8_gpio_7 = c2h_gpio_8_gpio_7_f;
   assign int_c2h_gpio_8_gpio_6 = c2h_gpio_8_gpio_6_f;
   assign int_c2h_gpio_8_gpio_5 = c2h_gpio_8_gpio_5_f;
   assign int_c2h_gpio_8_gpio_4 = c2h_gpio_8_gpio_4_f;
   assign int_c2h_gpio_8_gpio_3 = c2h_gpio_8_gpio_3_f;
   assign int_c2h_gpio_8_gpio_2 = c2h_gpio_8_gpio_2_f;
   assign int_c2h_gpio_8_gpio_1 = c2h_gpio_8_gpio_1_f;
   assign int_c2h_gpio_8_gpio_0 = c2h_gpio_8_gpio_0_f;
   assign int_c2h_gpio_9_gpio_31 = c2h_gpio_9_gpio_31_f;
   assign int_c2h_gpio_9_gpio_30 = c2h_gpio_9_gpio_30_f;
   assign int_c2h_gpio_9_gpio_29 = c2h_gpio_9_gpio_29_f;
   assign int_c2h_gpio_9_gpio_28 = c2h_gpio_9_gpio_28_f;
   assign int_c2h_gpio_9_gpio_27 = c2h_gpio_9_gpio_27_f;
   assign int_c2h_gpio_9_gpio_26 = c2h_gpio_9_gpio_26_f;
   assign int_c2h_gpio_9_gpio_25 = c2h_gpio_9_gpio_25_f;
   assign int_c2h_gpio_9_gpio_24 = c2h_gpio_9_gpio_24_f;
   assign int_c2h_gpio_9_gpio_23 = c2h_gpio_9_gpio_23_f;
   assign int_c2h_gpio_9_gpio_22 = c2h_gpio_9_gpio_22_f;
   assign int_c2h_gpio_9_gpio_21 = c2h_gpio_9_gpio_21_f;
   assign int_c2h_gpio_9_gpio_20 = c2h_gpio_9_gpio_20_f;
   assign int_c2h_gpio_9_gpio_19 = c2h_gpio_9_gpio_19_f;
   assign int_c2h_gpio_9_gpio_18 = c2h_gpio_9_gpio_18_f;
   assign int_c2h_gpio_9_gpio_17 = c2h_gpio_9_gpio_17_f;
   assign int_c2h_gpio_9_gpio_16 = c2h_gpio_9_gpio_16_f;
   assign int_c2h_gpio_9_gpio_15 = c2h_gpio_9_gpio_15_f;
   assign int_c2h_gpio_9_gpio_14 = c2h_gpio_9_gpio_14_f;
   assign int_c2h_gpio_9_gpio_13 = c2h_gpio_9_gpio_13_f;
   assign int_c2h_gpio_9_gpio_12 = c2h_gpio_9_gpio_12_f;
   assign int_c2h_gpio_9_gpio_11 = c2h_gpio_9_gpio_11_f;
   assign int_c2h_gpio_9_gpio_10 = c2h_gpio_9_gpio_10_f;
   assign int_c2h_gpio_9_gpio_9 = c2h_gpio_9_gpio_9_f;
   assign int_c2h_gpio_9_gpio_8 = c2h_gpio_9_gpio_8_f;
   assign int_c2h_gpio_9_gpio_7 = c2h_gpio_9_gpio_7_f;
   assign int_c2h_gpio_9_gpio_6 = c2h_gpio_9_gpio_6_f;
   assign int_c2h_gpio_9_gpio_5 = c2h_gpio_9_gpio_5_f;
   assign int_c2h_gpio_9_gpio_4 = c2h_gpio_9_gpio_4_f;
   assign int_c2h_gpio_9_gpio_3 = c2h_gpio_9_gpio_3_f;
   assign int_c2h_gpio_9_gpio_2 = c2h_gpio_9_gpio_2_f;
   assign int_c2h_gpio_9_gpio_1 = c2h_gpio_9_gpio_1_f;
   assign int_c2h_gpio_9_gpio_0 = c2h_gpio_9_gpio_0_f;
   assign int_c2h_gpio_10_gpio_31 = c2h_gpio_10_gpio_31_f;
   assign int_c2h_gpio_10_gpio_30 = c2h_gpio_10_gpio_30_f;
   assign int_c2h_gpio_10_gpio_29 = c2h_gpio_10_gpio_29_f;
   assign int_c2h_gpio_10_gpio_28 = c2h_gpio_10_gpio_28_f;
   assign int_c2h_gpio_10_gpio_27 = c2h_gpio_10_gpio_27_f;
   assign int_c2h_gpio_10_gpio_26 = c2h_gpio_10_gpio_26_f;
   assign int_c2h_gpio_10_gpio_25 = c2h_gpio_10_gpio_25_f;
   assign int_c2h_gpio_10_gpio_24 = c2h_gpio_10_gpio_24_f;
   assign int_c2h_gpio_10_gpio_23 = c2h_gpio_10_gpio_23_f;
   assign int_c2h_gpio_10_gpio_22 = c2h_gpio_10_gpio_22_f;
   assign int_c2h_gpio_10_gpio_21 = c2h_gpio_10_gpio_21_f;
   assign int_c2h_gpio_10_gpio_20 = c2h_gpio_10_gpio_20_f;
   assign int_c2h_gpio_10_gpio_19 = c2h_gpio_10_gpio_19_f;
   assign int_c2h_gpio_10_gpio_18 = c2h_gpio_10_gpio_18_f;
   assign int_c2h_gpio_10_gpio_17 = c2h_gpio_10_gpio_17_f;
   assign int_c2h_gpio_10_gpio_16 = c2h_gpio_10_gpio_16_f;
   assign int_c2h_gpio_10_gpio_15 = c2h_gpio_10_gpio_15_f;
   assign int_c2h_gpio_10_gpio_14 = c2h_gpio_10_gpio_14_f;
   assign int_c2h_gpio_10_gpio_13 = c2h_gpio_10_gpio_13_f;
   assign int_c2h_gpio_10_gpio_12 = c2h_gpio_10_gpio_12_f;
   assign int_c2h_gpio_10_gpio_11 = c2h_gpio_10_gpio_11_f;
   assign int_c2h_gpio_10_gpio_10 = c2h_gpio_10_gpio_10_f;
   assign int_c2h_gpio_10_gpio_9 = c2h_gpio_10_gpio_9_f;
   assign int_c2h_gpio_10_gpio_8 = c2h_gpio_10_gpio_8_f;
   assign int_c2h_gpio_10_gpio_7 = c2h_gpio_10_gpio_7_f;
   assign int_c2h_gpio_10_gpio_6 = c2h_gpio_10_gpio_6_f;
   assign int_c2h_gpio_10_gpio_5 = c2h_gpio_10_gpio_5_f;
   assign int_c2h_gpio_10_gpio_4 = c2h_gpio_10_gpio_4_f;
   assign int_c2h_gpio_10_gpio_3 = c2h_gpio_10_gpio_3_f;
   assign int_c2h_gpio_10_gpio_2 = c2h_gpio_10_gpio_2_f;
   assign int_c2h_gpio_10_gpio_1 = c2h_gpio_10_gpio_1_f;
   assign int_c2h_gpio_10_gpio_0 = c2h_gpio_10_gpio_0_f;
   assign int_c2h_gpio_11_gpio_31 = c2h_gpio_11_gpio_31_f;
   assign int_c2h_gpio_11_gpio_30 = c2h_gpio_11_gpio_30_f;
   assign int_c2h_gpio_11_gpio_29 = c2h_gpio_11_gpio_29_f;
   assign int_c2h_gpio_11_gpio_28 = c2h_gpio_11_gpio_28_f;
   assign int_c2h_gpio_11_gpio_27 = c2h_gpio_11_gpio_27_f;
   assign int_c2h_gpio_11_gpio_26 = c2h_gpio_11_gpio_26_f;
   assign int_c2h_gpio_11_gpio_25 = c2h_gpio_11_gpio_25_f;
   assign int_c2h_gpio_11_gpio_24 = c2h_gpio_11_gpio_24_f;
   assign int_c2h_gpio_11_gpio_23 = c2h_gpio_11_gpio_23_f;
   assign int_c2h_gpio_11_gpio_22 = c2h_gpio_11_gpio_22_f;
   assign int_c2h_gpio_11_gpio_21 = c2h_gpio_11_gpio_21_f;
   assign int_c2h_gpio_11_gpio_20 = c2h_gpio_11_gpio_20_f;
   assign int_c2h_gpio_11_gpio_19 = c2h_gpio_11_gpio_19_f;
   assign int_c2h_gpio_11_gpio_18 = c2h_gpio_11_gpio_18_f;
   assign int_c2h_gpio_11_gpio_17 = c2h_gpio_11_gpio_17_f;
   assign int_c2h_gpio_11_gpio_16 = c2h_gpio_11_gpio_16_f;
   assign int_c2h_gpio_11_gpio_15 = c2h_gpio_11_gpio_15_f;
   assign int_c2h_gpio_11_gpio_14 = c2h_gpio_11_gpio_14_f;
   assign int_c2h_gpio_11_gpio_13 = c2h_gpio_11_gpio_13_f;
   assign int_c2h_gpio_11_gpio_12 = c2h_gpio_11_gpio_12_f;
   assign int_c2h_gpio_11_gpio_11 = c2h_gpio_11_gpio_11_f;
   assign int_c2h_gpio_11_gpio_10 = c2h_gpio_11_gpio_10_f;
   assign int_c2h_gpio_11_gpio_9 = c2h_gpio_11_gpio_9_f;
   assign int_c2h_gpio_11_gpio_8 = c2h_gpio_11_gpio_8_f;
   assign int_c2h_gpio_11_gpio_7 = c2h_gpio_11_gpio_7_f;
   assign int_c2h_gpio_11_gpio_6 = c2h_gpio_11_gpio_6_f;
   assign int_c2h_gpio_11_gpio_5 = c2h_gpio_11_gpio_5_f;
   assign int_c2h_gpio_11_gpio_4 = c2h_gpio_11_gpio_4_f;
   assign int_c2h_gpio_11_gpio_3 = c2h_gpio_11_gpio_3_f;
   assign int_c2h_gpio_11_gpio_2 = c2h_gpio_11_gpio_2_f;
   assign int_c2h_gpio_11_gpio_1 = c2h_gpio_11_gpio_1_f;
   assign int_c2h_gpio_11_gpio_0 = c2h_gpio_11_gpio_0_f;
   assign int_c2h_gpio_12_gpio_31 = c2h_gpio_12_gpio_31_f;
   assign int_c2h_gpio_12_gpio_30 = c2h_gpio_12_gpio_30_f;
   assign int_c2h_gpio_12_gpio_29 = c2h_gpio_12_gpio_29_f;
   assign int_c2h_gpio_12_gpio_28 = c2h_gpio_12_gpio_28_f;
   assign int_c2h_gpio_12_gpio_27 = c2h_gpio_12_gpio_27_f;
   assign int_c2h_gpio_12_gpio_26 = c2h_gpio_12_gpio_26_f;
   assign int_c2h_gpio_12_gpio_25 = c2h_gpio_12_gpio_25_f;
   assign int_c2h_gpio_12_gpio_24 = c2h_gpio_12_gpio_24_f;
   assign int_c2h_gpio_12_gpio_23 = c2h_gpio_12_gpio_23_f;
   assign int_c2h_gpio_12_gpio_22 = c2h_gpio_12_gpio_22_f;
   assign int_c2h_gpio_12_gpio_21 = c2h_gpio_12_gpio_21_f;
   assign int_c2h_gpio_12_gpio_20 = c2h_gpio_12_gpio_20_f;
   assign int_c2h_gpio_12_gpio_19 = c2h_gpio_12_gpio_19_f;
   assign int_c2h_gpio_12_gpio_18 = c2h_gpio_12_gpio_18_f;
   assign int_c2h_gpio_12_gpio_17 = c2h_gpio_12_gpio_17_f;
   assign int_c2h_gpio_12_gpio_16 = c2h_gpio_12_gpio_16_f;
   assign int_c2h_gpio_12_gpio_15 = c2h_gpio_12_gpio_15_f;
   assign int_c2h_gpio_12_gpio_14 = c2h_gpio_12_gpio_14_f;
   assign int_c2h_gpio_12_gpio_13 = c2h_gpio_12_gpio_13_f;
   assign int_c2h_gpio_12_gpio_12 = c2h_gpio_12_gpio_12_f;
   assign int_c2h_gpio_12_gpio_11 = c2h_gpio_12_gpio_11_f;
   assign int_c2h_gpio_12_gpio_10 = c2h_gpio_12_gpio_10_f;
   assign int_c2h_gpio_12_gpio_9 = c2h_gpio_12_gpio_9_f;
   assign int_c2h_gpio_12_gpio_8 = c2h_gpio_12_gpio_8_f;
   assign int_c2h_gpio_12_gpio_7 = c2h_gpio_12_gpio_7_f;
   assign int_c2h_gpio_12_gpio_6 = c2h_gpio_12_gpio_6_f;
   assign int_c2h_gpio_12_gpio_5 = c2h_gpio_12_gpio_5_f;
   assign int_c2h_gpio_12_gpio_4 = c2h_gpio_12_gpio_4_f;
   assign int_c2h_gpio_12_gpio_3 = c2h_gpio_12_gpio_3_f;
   assign int_c2h_gpio_12_gpio_2 = c2h_gpio_12_gpio_2_f;
   assign int_c2h_gpio_12_gpio_1 = c2h_gpio_12_gpio_1_f;
   assign int_c2h_gpio_12_gpio_0 = c2h_gpio_12_gpio_0_f;
   assign int_c2h_gpio_13_gpio_31 = c2h_gpio_13_gpio_31_f;
   assign int_c2h_gpio_13_gpio_30 = c2h_gpio_13_gpio_30_f;
   assign int_c2h_gpio_13_gpio_29 = c2h_gpio_13_gpio_29_f;
   assign int_c2h_gpio_13_gpio_28 = c2h_gpio_13_gpio_28_f;
   assign int_c2h_gpio_13_gpio_27 = c2h_gpio_13_gpio_27_f;
   assign int_c2h_gpio_13_gpio_26 = c2h_gpio_13_gpio_26_f;
   assign int_c2h_gpio_13_gpio_25 = c2h_gpio_13_gpio_25_f;
   assign int_c2h_gpio_13_gpio_24 = c2h_gpio_13_gpio_24_f;
   assign int_c2h_gpio_13_gpio_23 = c2h_gpio_13_gpio_23_f;
   assign int_c2h_gpio_13_gpio_22 = c2h_gpio_13_gpio_22_f;
   assign int_c2h_gpio_13_gpio_21 = c2h_gpio_13_gpio_21_f;
   assign int_c2h_gpio_13_gpio_20 = c2h_gpio_13_gpio_20_f;
   assign int_c2h_gpio_13_gpio_19 = c2h_gpio_13_gpio_19_f;
   assign int_c2h_gpio_13_gpio_18 = c2h_gpio_13_gpio_18_f;
   assign int_c2h_gpio_13_gpio_17 = c2h_gpio_13_gpio_17_f;
   assign int_c2h_gpio_13_gpio_16 = c2h_gpio_13_gpio_16_f;
   assign int_c2h_gpio_13_gpio_15 = c2h_gpio_13_gpio_15_f;
   assign int_c2h_gpio_13_gpio_14 = c2h_gpio_13_gpio_14_f;
   assign int_c2h_gpio_13_gpio_13 = c2h_gpio_13_gpio_13_f;
   assign int_c2h_gpio_13_gpio_12 = c2h_gpio_13_gpio_12_f;
   assign int_c2h_gpio_13_gpio_11 = c2h_gpio_13_gpio_11_f;
   assign int_c2h_gpio_13_gpio_10 = c2h_gpio_13_gpio_10_f;
   assign int_c2h_gpio_13_gpio_9 = c2h_gpio_13_gpio_9_f;
   assign int_c2h_gpio_13_gpio_8 = c2h_gpio_13_gpio_8_f;
   assign int_c2h_gpio_13_gpio_7 = c2h_gpio_13_gpio_7_f;
   assign int_c2h_gpio_13_gpio_6 = c2h_gpio_13_gpio_6_f;
   assign int_c2h_gpio_13_gpio_5 = c2h_gpio_13_gpio_5_f;
   assign int_c2h_gpio_13_gpio_4 = c2h_gpio_13_gpio_4_f;
   assign int_c2h_gpio_13_gpio_3 = c2h_gpio_13_gpio_3_f;
   assign int_c2h_gpio_13_gpio_2 = c2h_gpio_13_gpio_2_f;
   assign int_c2h_gpio_13_gpio_1 = c2h_gpio_13_gpio_1_f;
   assign int_c2h_gpio_13_gpio_0 = c2h_gpio_13_gpio_0_f;
   assign int_c2h_gpio_14_gpio_31 = c2h_gpio_14_gpio_31_f;
   assign int_c2h_gpio_14_gpio_30 = c2h_gpio_14_gpio_30_f;
   assign int_c2h_gpio_14_gpio_29 = c2h_gpio_14_gpio_29_f;
   assign int_c2h_gpio_14_gpio_28 = c2h_gpio_14_gpio_28_f;
   assign int_c2h_gpio_14_gpio_27 = c2h_gpio_14_gpio_27_f;
   assign int_c2h_gpio_14_gpio_26 = c2h_gpio_14_gpio_26_f;
   assign int_c2h_gpio_14_gpio_25 = c2h_gpio_14_gpio_25_f;
   assign int_c2h_gpio_14_gpio_24 = c2h_gpio_14_gpio_24_f;
   assign int_c2h_gpio_14_gpio_23 = c2h_gpio_14_gpio_23_f;
   assign int_c2h_gpio_14_gpio_22 = c2h_gpio_14_gpio_22_f;
   assign int_c2h_gpio_14_gpio_21 = c2h_gpio_14_gpio_21_f;
   assign int_c2h_gpio_14_gpio_20 = c2h_gpio_14_gpio_20_f;
   assign int_c2h_gpio_14_gpio_19 = c2h_gpio_14_gpio_19_f;
   assign int_c2h_gpio_14_gpio_18 = c2h_gpio_14_gpio_18_f;
   assign int_c2h_gpio_14_gpio_17 = c2h_gpio_14_gpio_17_f;
   assign int_c2h_gpio_14_gpio_16 = c2h_gpio_14_gpio_16_f;
   assign int_c2h_gpio_14_gpio_15 = c2h_gpio_14_gpio_15_f;
   assign int_c2h_gpio_14_gpio_14 = c2h_gpio_14_gpio_14_f;
   assign int_c2h_gpio_14_gpio_13 = c2h_gpio_14_gpio_13_f;
   assign int_c2h_gpio_14_gpio_12 = c2h_gpio_14_gpio_12_f;
   assign int_c2h_gpio_14_gpio_11 = c2h_gpio_14_gpio_11_f;
   assign int_c2h_gpio_14_gpio_10 = c2h_gpio_14_gpio_10_f;
   assign int_c2h_gpio_14_gpio_9 = c2h_gpio_14_gpio_9_f;
   assign int_c2h_gpio_14_gpio_8 = c2h_gpio_14_gpio_8_f;
   assign int_c2h_gpio_14_gpio_7 = c2h_gpio_14_gpio_7_f;
   assign int_c2h_gpio_14_gpio_6 = c2h_gpio_14_gpio_6_f;
   assign int_c2h_gpio_14_gpio_5 = c2h_gpio_14_gpio_5_f;
   assign int_c2h_gpio_14_gpio_4 = c2h_gpio_14_gpio_4_f;
   assign int_c2h_gpio_14_gpio_3 = c2h_gpio_14_gpio_3_f;
   assign int_c2h_gpio_14_gpio_2 = c2h_gpio_14_gpio_2_f;
   assign int_c2h_gpio_14_gpio_1 = c2h_gpio_14_gpio_1_f;
   assign int_c2h_gpio_14_gpio_0 = c2h_gpio_14_gpio_0_f;
   assign int_c2h_gpio_15_gpio_31 = c2h_gpio_15_gpio_31_f;
   assign int_c2h_gpio_15_gpio_30 = c2h_gpio_15_gpio_30_f;
   assign int_c2h_gpio_15_gpio_29 = c2h_gpio_15_gpio_29_f;
   assign int_c2h_gpio_15_gpio_28 = c2h_gpio_15_gpio_28_f;
   assign int_c2h_gpio_15_gpio_27 = c2h_gpio_15_gpio_27_f;
   assign int_c2h_gpio_15_gpio_26 = c2h_gpio_15_gpio_26_f;
   assign int_c2h_gpio_15_gpio_25 = c2h_gpio_15_gpio_25_f;
   assign int_c2h_gpio_15_gpio_24 = c2h_gpio_15_gpio_24_f;
   assign int_c2h_gpio_15_gpio_23 = c2h_gpio_15_gpio_23_f;
   assign int_c2h_gpio_15_gpio_22 = c2h_gpio_15_gpio_22_f;
   assign int_c2h_gpio_15_gpio_21 = c2h_gpio_15_gpio_21_f;
   assign int_c2h_gpio_15_gpio_20 = c2h_gpio_15_gpio_20_f;
   assign int_c2h_gpio_15_gpio_19 = c2h_gpio_15_gpio_19_f;
   assign int_c2h_gpio_15_gpio_18 = c2h_gpio_15_gpio_18_f;
   assign int_c2h_gpio_15_gpio_17 = c2h_gpio_15_gpio_17_f;
   assign int_c2h_gpio_15_gpio_16 = c2h_gpio_15_gpio_16_f;
   assign int_c2h_gpio_15_gpio_15 = c2h_gpio_15_gpio_15_f;
   assign int_c2h_gpio_15_gpio_14 = c2h_gpio_15_gpio_14_f;
   assign int_c2h_gpio_15_gpio_13 = c2h_gpio_15_gpio_13_f;
   assign int_c2h_gpio_15_gpio_12 = c2h_gpio_15_gpio_12_f;
   assign int_c2h_gpio_15_gpio_11 = c2h_gpio_15_gpio_11_f;
   assign int_c2h_gpio_15_gpio_10 = c2h_gpio_15_gpio_10_f;
   assign int_c2h_gpio_15_gpio_9 = c2h_gpio_15_gpio_9_f;
   assign int_c2h_gpio_15_gpio_8 = c2h_gpio_15_gpio_8_f;
   assign int_c2h_gpio_15_gpio_7 = c2h_gpio_15_gpio_7_f;
   assign int_c2h_gpio_15_gpio_6 = c2h_gpio_15_gpio_6_f;
   assign int_c2h_gpio_15_gpio_5 = c2h_gpio_15_gpio_5_f;
   assign int_c2h_gpio_15_gpio_4 = c2h_gpio_15_gpio_4_f;
   assign int_c2h_gpio_15_gpio_3 = c2h_gpio_15_gpio_3_f;
   assign int_c2h_gpio_15_gpio_2 = c2h_gpio_15_gpio_2_f;
   assign int_c2h_gpio_15_gpio_1 = c2h_gpio_15_gpio_1_f;
   assign int_c2h_gpio_15_gpio_0 = c2h_gpio_15_gpio_0_f;
   assign int_h2c_gpio_0_gpio_31 = h2c_gpio_0_gpio_31_f;
   assign int_h2c_gpio_0_gpio_30 = h2c_gpio_0_gpio_30_f;
   assign int_h2c_gpio_0_gpio_29 = h2c_gpio_0_gpio_29_f;
   assign int_h2c_gpio_0_gpio_28 = h2c_gpio_0_gpio_28_f;
   assign int_h2c_gpio_0_gpio_27 = h2c_gpio_0_gpio_27_f;
   assign int_h2c_gpio_0_gpio_26 = h2c_gpio_0_gpio_26_f;
   assign int_h2c_gpio_0_gpio_25 = h2c_gpio_0_gpio_25_f;
   assign int_h2c_gpio_0_gpio_24 = h2c_gpio_0_gpio_24_f;
   assign int_h2c_gpio_0_gpio_23 = h2c_gpio_0_gpio_23_f;
   assign int_h2c_gpio_0_gpio_22 = h2c_gpio_0_gpio_22_f;
   assign int_h2c_gpio_0_gpio_21 = h2c_gpio_0_gpio_21_f;
   assign int_h2c_gpio_0_gpio_20 = h2c_gpio_0_gpio_20_f;
   assign int_h2c_gpio_0_gpio_19 = h2c_gpio_0_gpio_19_f;
   assign int_h2c_gpio_0_gpio_18 = h2c_gpio_0_gpio_18_f;
   assign int_h2c_gpio_0_gpio_17 = h2c_gpio_0_gpio_17_f;
   assign int_h2c_gpio_0_gpio_16 = h2c_gpio_0_gpio_16_f;
   assign int_h2c_gpio_0_gpio_15 = h2c_gpio_0_gpio_15_f;
   assign int_h2c_gpio_0_gpio_14 = h2c_gpio_0_gpio_14_f;
   assign int_h2c_gpio_0_gpio_13 = h2c_gpio_0_gpio_13_f;
   assign int_h2c_gpio_0_gpio_12 = h2c_gpio_0_gpio_12_f;
   assign int_h2c_gpio_0_gpio_11 = h2c_gpio_0_gpio_11_f;
   assign int_h2c_gpio_0_gpio_10 = h2c_gpio_0_gpio_10_f;
   assign int_h2c_gpio_0_gpio_9 = h2c_gpio_0_gpio_9_f;
   assign int_h2c_gpio_0_gpio_8 = h2c_gpio_0_gpio_8_f;
   assign int_h2c_gpio_0_gpio_7 = h2c_gpio_0_gpio_7_f;
   assign int_h2c_gpio_0_gpio_6 = h2c_gpio_0_gpio_6_f;
   assign int_h2c_gpio_0_gpio_5 = h2c_gpio_0_gpio_5_f;
   assign int_h2c_gpio_0_gpio_4 = h2c_gpio_0_gpio_4_f;
   assign int_h2c_gpio_0_gpio_3 = h2c_gpio_0_gpio_3_f;
   assign int_h2c_gpio_0_gpio_2 = h2c_gpio_0_gpio_2_f;
   assign int_h2c_gpio_0_gpio_1 = h2c_gpio_0_gpio_1_f;
   assign int_h2c_gpio_0_gpio_0 = h2c_gpio_0_gpio_0_f;
   assign int_h2c_gpio_1_gpio_31 = h2c_gpio_1_gpio_31_f;
   assign int_h2c_gpio_1_gpio_30 = h2c_gpio_1_gpio_30_f;
   assign int_h2c_gpio_1_gpio_29 = h2c_gpio_1_gpio_29_f;
   assign int_h2c_gpio_1_gpio_28 = h2c_gpio_1_gpio_28_f;
   assign int_h2c_gpio_1_gpio_27 = h2c_gpio_1_gpio_27_f;
   assign int_h2c_gpio_1_gpio_26 = h2c_gpio_1_gpio_26_f;
   assign int_h2c_gpio_1_gpio_25 = h2c_gpio_1_gpio_25_f;
   assign int_h2c_gpio_1_gpio_24 = h2c_gpio_1_gpio_24_f;
   assign int_h2c_gpio_1_gpio_23 = h2c_gpio_1_gpio_23_f;
   assign int_h2c_gpio_1_gpio_22 = h2c_gpio_1_gpio_22_f;
   assign int_h2c_gpio_1_gpio_21 = h2c_gpio_1_gpio_21_f;
   assign int_h2c_gpio_1_gpio_20 = h2c_gpio_1_gpio_20_f;
   assign int_h2c_gpio_1_gpio_19 = h2c_gpio_1_gpio_19_f;
   assign int_h2c_gpio_1_gpio_18 = h2c_gpio_1_gpio_18_f;
   assign int_h2c_gpio_1_gpio_17 = h2c_gpio_1_gpio_17_f;
   assign int_h2c_gpio_1_gpio_16 = h2c_gpio_1_gpio_16_f;
   assign int_h2c_gpio_1_gpio_15 = h2c_gpio_1_gpio_15_f;
   assign int_h2c_gpio_1_gpio_14 = h2c_gpio_1_gpio_14_f;
   assign int_h2c_gpio_1_gpio_13 = h2c_gpio_1_gpio_13_f;
   assign int_h2c_gpio_1_gpio_12 = h2c_gpio_1_gpio_12_f;
   assign int_h2c_gpio_1_gpio_11 = h2c_gpio_1_gpio_11_f;
   assign int_h2c_gpio_1_gpio_10 = h2c_gpio_1_gpio_10_f;
   assign int_h2c_gpio_1_gpio_9 = h2c_gpio_1_gpio_9_f;
   assign int_h2c_gpio_1_gpio_8 = h2c_gpio_1_gpio_8_f;
   assign int_h2c_gpio_1_gpio_7 = h2c_gpio_1_gpio_7_f;
   assign int_h2c_gpio_1_gpio_6 = h2c_gpio_1_gpio_6_f;
   assign int_h2c_gpio_1_gpio_5 = h2c_gpio_1_gpio_5_f;
   assign int_h2c_gpio_1_gpio_4 = h2c_gpio_1_gpio_4_f;
   assign int_h2c_gpio_1_gpio_3 = h2c_gpio_1_gpio_3_f;
   assign int_h2c_gpio_1_gpio_2 = h2c_gpio_1_gpio_2_f;
   assign int_h2c_gpio_1_gpio_1 = h2c_gpio_1_gpio_1_f;
   assign int_h2c_gpio_1_gpio_0 = h2c_gpio_1_gpio_0_f;
   assign int_h2c_gpio_2_gpio_31 = h2c_gpio_2_gpio_31_f;
   assign int_h2c_gpio_2_gpio_30 = h2c_gpio_2_gpio_30_f;
   assign int_h2c_gpio_2_gpio_29 = h2c_gpio_2_gpio_29_f;
   assign int_h2c_gpio_2_gpio_28 = h2c_gpio_2_gpio_28_f;
   assign int_h2c_gpio_2_gpio_27 = h2c_gpio_2_gpio_27_f;
   assign int_h2c_gpio_2_gpio_26 = h2c_gpio_2_gpio_26_f;
   assign int_h2c_gpio_2_gpio_25 = h2c_gpio_2_gpio_25_f;
   assign int_h2c_gpio_2_gpio_24 = h2c_gpio_2_gpio_24_f;
   assign int_h2c_gpio_2_gpio_23 = h2c_gpio_2_gpio_23_f;
   assign int_h2c_gpio_2_gpio_22 = h2c_gpio_2_gpio_22_f;
   assign int_h2c_gpio_2_gpio_21 = h2c_gpio_2_gpio_21_f;
   assign int_h2c_gpio_2_gpio_20 = h2c_gpio_2_gpio_20_f;
   assign int_h2c_gpio_2_gpio_19 = h2c_gpio_2_gpio_19_f;
   assign int_h2c_gpio_2_gpio_18 = h2c_gpio_2_gpio_18_f;
   assign int_h2c_gpio_2_gpio_17 = h2c_gpio_2_gpio_17_f;
   assign int_h2c_gpio_2_gpio_16 = h2c_gpio_2_gpio_16_f;
   assign int_h2c_gpio_2_gpio_15 = h2c_gpio_2_gpio_15_f;
   assign int_h2c_gpio_2_gpio_14 = h2c_gpio_2_gpio_14_f;
   assign int_h2c_gpio_2_gpio_13 = h2c_gpio_2_gpio_13_f;
   assign int_h2c_gpio_2_gpio_12 = h2c_gpio_2_gpio_12_f;
   assign int_h2c_gpio_2_gpio_11 = h2c_gpio_2_gpio_11_f;
   assign int_h2c_gpio_2_gpio_10 = h2c_gpio_2_gpio_10_f;
   assign int_h2c_gpio_2_gpio_9 = h2c_gpio_2_gpio_9_f;
   assign int_h2c_gpio_2_gpio_8 = h2c_gpio_2_gpio_8_f;
   assign int_h2c_gpio_2_gpio_7 = h2c_gpio_2_gpio_7_f;
   assign int_h2c_gpio_2_gpio_6 = h2c_gpio_2_gpio_6_f;
   assign int_h2c_gpio_2_gpio_5 = h2c_gpio_2_gpio_5_f;
   assign int_h2c_gpio_2_gpio_4 = h2c_gpio_2_gpio_4_f;
   assign int_h2c_gpio_2_gpio_3 = h2c_gpio_2_gpio_3_f;
   assign int_h2c_gpio_2_gpio_2 = h2c_gpio_2_gpio_2_f;
   assign int_h2c_gpio_2_gpio_1 = h2c_gpio_2_gpio_1_f;
   assign int_h2c_gpio_2_gpio_0 = h2c_gpio_2_gpio_0_f;
   assign int_h2c_gpio_3_gpio_31 = h2c_gpio_3_gpio_31_f;
   assign int_h2c_gpio_3_gpio_30 = h2c_gpio_3_gpio_30_f;
   assign int_h2c_gpio_3_gpio_29 = h2c_gpio_3_gpio_29_f;
   assign int_h2c_gpio_3_gpio_28 = h2c_gpio_3_gpio_28_f;
   assign int_h2c_gpio_3_gpio_27 = h2c_gpio_3_gpio_27_f;
   assign int_h2c_gpio_3_gpio_26 = h2c_gpio_3_gpio_26_f;
   assign int_h2c_gpio_3_gpio_25 = h2c_gpio_3_gpio_25_f;
   assign int_h2c_gpio_3_gpio_24 = h2c_gpio_3_gpio_24_f;
   assign int_h2c_gpio_3_gpio_23 = h2c_gpio_3_gpio_23_f;
   assign int_h2c_gpio_3_gpio_22 = h2c_gpio_3_gpio_22_f;
   assign int_h2c_gpio_3_gpio_21 = h2c_gpio_3_gpio_21_f;
   assign int_h2c_gpio_3_gpio_20 = h2c_gpio_3_gpio_20_f;
   assign int_h2c_gpio_3_gpio_19 = h2c_gpio_3_gpio_19_f;
   assign int_h2c_gpio_3_gpio_18 = h2c_gpio_3_gpio_18_f;
   assign int_h2c_gpio_3_gpio_17 = h2c_gpio_3_gpio_17_f;
   assign int_h2c_gpio_3_gpio_16 = h2c_gpio_3_gpio_16_f;
   assign int_h2c_gpio_3_gpio_15 = h2c_gpio_3_gpio_15_f;
   assign int_h2c_gpio_3_gpio_14 = h2c_gpio_3_gpio_14_f;
   assign int_h2c_gpio_3_gpio_13 = h2c_gpio_3_gpio_13_f;
   assign int_h2c_gpio_3_gpio_12 = h2c_gpio_3_gpio_12_f;
   assign int_h2c_gpio_3_gpio_11 = h2c_gpio_3_gpio_11_f;
   assign int_h2c_gpio_3_gpio_10 = h2c_gpio_3_gpio_10_f;
   assign int_h2c_gpio_3_gpio_9 = h2c_gpio_3_gpio_9_f;
   assign int_h2c_gpio_3_gpio_8 = h2c_gpio_3_gpio_8_f;
   assign int_h2c_gpio_3_gpio_7 = h2c_gpio_3_gpio_7_f;
   assign int_h2c_gpio_3_gpio_6 = h2c_gpio_3_gpio_6_f;
   assign int_h2c_gpio_3_gpio_5 = h2c_gpio_3_gpio_5_f;
   assign int_h2c_gpio_3_gpio_4 = h2c_gpio_3_gpio_4_f;
   assign int_h2c_gpio_3_gpio_3 = h2c_gpio_3_gpio_3_f;
   assign int_h2c_gpio_3_gpio_2 = h2c_gpio_3_gpio_2_f;
   assign int_h2c_gpio_3_gpio_1 = h2c_gpio_3_gpio_1_f;
   assign int_h2c_gpio_3_gpio_0 = h2c_gpio_3_gpio_0_f;
   assign int_h2c_gpio_4_gpio_31 = h2c_gpio_4_gpio_31_f;
   assign int_h2c_gpio_4_gpio_30 = h2c_gpio_4_gpio_30_f;
   assign int_h2c_gpio_4_gpio_29 = h2c_gpio_4_gpio_29_f;
   assign int_h2c_gpio_4_gpio_28 = h2c_gpio_4_gpio_28_f;
   assign int_h2c_gpio_4_gpio_27 = h2c_gpio_4_gpio_27_f;
   assign int_h2c_gpio_4_gpio_26 = h2c_gpio_4_gpio_26_f;
   assign int_h2c_gpio_4_gpio_25 = h2c_gpio_4_gpio_25_f;
   assign int_h2c_gpio_4_gpio_24 = h2c_gpio_4_gpio_24_f;
   assign int_h2c_gpio_4_gpio_23 = h2c_gpio_4_gpio_23_f;
   assign int_h2c_gpio_4_gpio_22 = h2c_gpio_4_gpio_22_f;
   assign int_h2c_gpio_4_gpio_21 = h2c_gpio_4_gpio_21_f;
   assign int_h2c_gpio_4_gpio_20 = h2c_gpio_4_gpio_20_f;
   assign int_h2c_gpio_4_gpio_19 = h2c_gpio_4_gpio_19_f;
   assign int_h2c_gpio_4_gpio_18 = h2c_gpio_4_gpio_18_f;
   assign int_h2c_gpio_4_gpio_17 = h2c_gpio_4_gpio_17_f;
   assign int_h2c_gpio_4_gpio_16 = h2c_gpio_4_gpio_16_f;
   assign int_h2c_gpio_4_gpio_15 = h2c_gpio_4_gpio_15_f;
   assign int_h2c_gpio_4_gpio_14 = h2c_gpio_4_gpio_14_f;
   assign int_h2c_gpio_4_gpio_13 = h2c_gpio_4_gpio_13_f;
   assign int_h2c_gpio_4_gpio_12 = h2c_gpio_4_gpio_12_f;
   assign int_h2c_gpio_4_gpio_11 = h2c_gpio_4_gpio_11_f;
   assign int_h2c_gpio_4_gpio_10 = h2c_gpio_4_gpio_10_f;
   assign int_h2c_gpio_4_gpio_9 = h2c_gpio_4_gpio_9_f;
   assign int_h2c_gpio_4_gpio_8 = h2c_gpio_4_gpio_8_f;
   assign int_h2c_gpio_4_gpio_7 = h2c_gpio_4_gpio_7_f;
   assign int_h2c_gpio_4_gpio_6 = h2c_gpio_4_gpio_6_f;
   assign int_h2c_gpio_4_gpio_5 = h2c_gpio_4_gpio_5_f;
   assign int_h2c_gpio_4_gpio_4 = h2c_gpio_4_gpio_4_f;
   assign int_h2c_gpio_4_gpio_3 = h2c_gpio_4_gpio_3_f;
   assign int_h2c_gpio_4_gpio_2 = h2c_gpio_4_gpio_2_f;
   assign int_h2c_gpio_4_gpio_1 = h2c_gpio_4_gpio_1_f;
   assign int_h2c_gpio_4_gpio_0 = h2c_gpio_4_gpio_0_f;
   assign int_h2c_gpio_5_gpio_31 = h2c_gpio_5_gpio_31_f;
   assign int_h2c_gpio_5_gpio_30 = h2c_gpio_5_gpio_30_f;
   assign int_h2c_gpio_5_gpio_29 = h2c_gpio_5_gpio_29_f;
   assign int_h2c_gpio_5_gpio_28 = h2c_gpio_5_gpio_28_f;
   assign int_h2c_gpio_5_gpio_27 = h2c_gpio_5_gpio_27_f;
   assign int_h2c_gpio_5_gpio_26 = h2c_gpio_5_gpio_26_f;
   assign int_h2c_gpio_5_gpio_25 = h2c_gpio_5_gpio_25_f;
   assign int_h2c_gpio_5_gpio_24 = h2c_gpio_5_gpio_24_f;
   assign int_h2c_gpio_5_gpio_23 = h2c_gpio_5_gpio_23_f;
   assign int_h2c_gpio_5_gpio_22 = h2c_gpio_5_gpio_22_f;
   assign int_h2c_gpio_5_gpio_21 = h2c_gpio_5_gpio_21_f;
   assign int_h2c_gpio_5_gpio_20 = h2c_gpio_5_gpio_20_f;
   assign int_h2c_gpio_5_gpio_19 = h2c_gpio_5_gpio_19_f;
   assign int_h2c_gpio_5_gpio_18 = h2c_gpio_5_gpio_18_f;
   assign int_h2c_gpio_5_gpio_17 = h2c_gpio_5_gpio_17_f;
   assign int_h2c_gpio_5_gpio_16 = h2c_gpio_5_gpio_16_f;
   assign int_h2c_gpio_5_gpio_15 = h2c_gpio_5_gpio_15_f;
   assign int_h2c_gpio_5_gpio_14 = h2c_gpio_5_gpio_14_f;
   assign int_h2c_gpio_5_gpio_13 = h2c_gpio_5_gpio_13_f;
   assign int_h2c_gpio_5_gpio_12 = h2c_gpio_5_gpio_12_f;
   assign int_h2c_gpio_5_gpio_11 = h2c_gpio_5_gpio_11_f;
   assign int_h2c_gpio_5_gpio_10 = h2c_gpio_5_gpio_10_f;
   assign int_h2c_gpio_5_gpio_9 = h2c_gpio_5_gpio_9_f;
   assign int_h2c_gpio_5_gpio_8 = h2c_gpio_5_gpio_8_f;
   assign int_h2c_gpio_5_gpio_7 = h2c_gpio_5_gpio_7_f;
   assign int_h2c_gpio_5_gpio_6 = h2c_gpio_5_gpio_6_f;
   assign int_h2c_gpio_5_gpio_5 = h2c_gpio_5_gpio_5_f;
   assign int_h2c_gpio_5_gpio_4 = h2c_gpio_5_gpio_4_f;
   assign int_h2c_gpio_5_gpio_3 = h2c_gpio_5_gpio_3_f;
   assign int_h2c_gpio_5_gpio_2 = h2c_gpio_5_gpio_2_f;
   assign int_h2c_gpio_5_gpio_1 = h2c_gpio_5_gpio_1_f;
   assign int_h2c_gpio_5_gpio_0 = h2c_gpio_5_gpio_0_f;
   assign int_h2c_gpio_6_gpio_31 = h2c_gpio_6_gpio_31_f;
   assign int_h2c_gpio_6_gpio_30 = h2c_gpio_6_gpio_30_f;
   assign int_h2c_gpio_6_gpio_29 = h2c_gpio_6_gpio_29_f;
   assign int_h2c_gpio_6_gpio_28 = h2c_gpio_6_gpio_28_f;
   assign int_h2c_gpio_6_gpio_27 = h2c_gpio_6_gpio_27_f;
   assign int_h2c_gpio_6_gpio_26 = h2c_gpio_6_gpio_26_f;
   assign int_h2c_gpio_6_gpio_25 = h2c_gpio_6_gpio_25_f;
   assign int_h2c_gpio_6_gpio_24 = h2c_gpio_6_gpio_24_f;
   assign int_h2c_gpio_6_gpio_23 = h2c_gpio_6_gpio_23_f;
   assign int_h2c_gpio_6_gpio_22 = h2c_gpio_6_gpio_22_f;
   assign int_h2c_gpio_6_gpio_21 = h2c_gpio_6_gpio_21_f;
   assign int_h2c_gpio_6_gpio_20 = h2c_gpio_6_gpio_20_f;
   assign int_h2c_gpio_6_gpio_19 = h2c_gpio_6_gpio_19_f;
   assign int_h2c_gpio_6_gpio_18 = h2c_gpio_6_gpio_18_f;
   assign int_h2c_gpio_6_gpio_17 = h2c_gpio_6_gpio_17_f;
   assign int_h2c_gpio_6_gpio_16 = h2c_gpio_6_gpio_16_f;
   assign int_h2c_gpio_6_gpio_15 = h2c_gpio_6_gpio_15_f;
   assign int_h2c_gpio_6_gpio_14 = h2c_gpio_6_gpio_14_f;
   assign int_h2c_gpio_6_gpio_13 = h2c_gpio_6_gpio_13_f;
   assign int_h2c_gpio_6_gpio_12 = h2c_gpio_6_gpio_12_f;
   assign int_h2c_gpio_6_gpio_11 = h2c_gpio_6_gpio_11_f;
   assign int_h2c_gpio_6_gpio_10 = h2c_gpio_6_gpio_10_f;
   assign int_h2c_gpio_6_gpio_9 = h2c_gpio_6_gpio_9_f;
   assign int_h2c_gpio_6_gpio_8 = h2c_gpio_6_gpio_8_f;
   assign int_h2c_gpio_6_gpio_7 = h2c_gpio_6_gpio_7_f;
   assign int_h2c_gpio_6_gpio_6 = h2c_gpio_6_gpio_6_f;
   assign int_h2c_gpio_6_gpio_5 = h2c_gpio_6_gpio_5_f;
   assign int_h2c_gpio_6_gpio_4 = h2c_gpio_6_gpio_4_f;
   assign int_h2c_gpio_6_gpio_3 = h2c_gpio_6_gpio_3_f;
   assign int_h2c_gpio_6_gpio_2 = h2c_gpio_6_gpio_2_f;
   assign int_h2c_gpio_6_gpio_1 = h2c_gpio_6_gpio_1_f;
   assign int_h2c_gpio_6_gpio_0 = h2c_gpio_6_gpio_0_f;
   assign int_h2c_gpio_7_gpio_31 = h2c_gpio_7_gpio_31_f;
   assign int_h2c_gpio_7_gpio_30 = h2c_gpio_7_gpio_30_f;
   assign int_h2c_gpio_7_gpio_29 = h2c_gpio_7_gpio_29_f;
   assign int_h2c_gpio_7_gpio_28 = h2c_gpio_7_gpio_28_f;
   assign int_h2c_gpio_7_gpio_27 = h2c_gpio_7_gpio_27_f;
   assign int_h2c_gpio_7_gpio_26 = h2c_gpio_7_gpio_26_f;
   assign int_h2c_gpio_7_gpio_25 = h2c_gpio_7_gpio_25_f;
   assign int_h2c_gpio_7_gpio_24 = h2c_gpio_7_gpio_24_f;
   assign int_h2c_gpio_7_gpio_23 = h2c_gpio_7_gpio_23_f;
   assign int_h2c_gpio_7_gpio_22 = h2c_gpio_7_gpio_22_f;
   assign int_h2c_gpio_7_gpio_21 = h2c_gpio_7_gpio_21_f;
   assign int_h2c_gpio_7_gpio_20 = h2c_gpio_7_gpio_20_f;
   assign int_h2c_gpio_7_gpio_19 = h2c_gpio_7_gpio_19_f;
   assign int_h2c_gpio_7_gpio_18 = h2c_gpio_7_gpio_18_f;
   assign int_h2c_gpio_7_gpio_17 = h2c_gpio_7_gpio_17_f;
   assign int_h2c_gpio_7_gpio_16 = h2c_gpio_7_gpio_16_f;
   assign int_h2c_gpio_7_gpio_15 = h2c_gpio_7_gpio_15_f;
   assign int_h2c_gpio_7_gpio_14 = h2c_gpio_7_gpio_14_f;
   assign int_h2c_gpio_7_gpio_13 = h2c_gpio_7_gpio_13_f;
   assign int_h2c_gpio_7_gpio_12 = h2c_gpio_7_gpio_12_f;
   assign int_h2c_gpio_7_gpio_11 = h2c_gpio_7_gpio_11_f;
   assign int_h2c_gpio_7_gpio_10 = h2c_gpio_7_gpio_10_f;
   assign int_h2c_gpio_7_gpio_9 = h2c_gpio_7_gpio_9_f;
   assign int_h2c_gpio_7_gpio_8 = h2c_gpio_7_gpio_8_f;
   assign int_h2c_gpio_7_gpio_7 = h2c_gpio_7_gpio_7_f;
   assign int_h2c_gpio_7_gpio_6 = h2c_gpio_7_gpio_6_f;
   assign int_h2c_gpio_7_gpio_5 = h2c_gpio_7_gpio_5_f;
   assign int_h2c_gpio_7_gpio_4 = h2c_gpio_7_gpio_4_f;
   assign int_h2c_gpio_7_gpio_3 = h2c_gpio_7_gpio_3_f;
   assign int_h2c_gpio_7_gpio_2 = h2c_gpio_7_gpio_2_f;
   assign int_h2c_gpio_7_gpio_1 = h2c_gpio_7_gpio_1_f;
   assign int_h2c_gpio_7_gpio_0 = h2c_gpio_7_gpio_0_f;
   assign int_h2c_gpio_8_gpio_31 = h2c_gpio_8_gpio_31_f;
   assign int_h2c_gpio_8_gpio_30 = h2c_gpio_8_gpio_30_f;
   assign int_h2c_gpio_8_gpio_29 = h2c_gpio_8_gpio_29_f;
   assign int_h2c_gpio_8_gpio_28 = h2c_gpio_8_gpio_28_f;
   assign int_h2c_gpio_8_gpio_27 = h2c_gpio_8_gpio_27_f;
   assign int_h2c_gpio_8_gpio_26 = h2c_gpio_8_gpio_26_f;
   assign int_h2c_gpio_8_gpio_25 = h2c_gpio_8_gpio_25_f;
   assign int_h2c_gpio_8_gpio_24 = h2c_gpio_8_gpio_24_f;
   assign int_h2c_gpio_8_gpio_23 = h2c_gpio_8_gpio_23_f;
   assign int_h2c_gpio_8_gpio_22 = h2c_gpio_8_gpio_22_f;
   assign int_h2c_gpio_8_gpio_21 = h2c_gpio_8_gpio_21_f;
   assign int_h2c_gpio_8_gpio_20 = h2c_gpio_8_gpio_20_f;
   assign int_h2c_gpio_8_gpio_19 = h2c_gpio_8_gpio_19_f;
   assign int_h2c_gpio_8_gpio_18 = h2c_gpio_8_gpio_18_f;
   assign int_h2c_gpio_8_gpio_17 = h2c_gpio_8_gpio_17_f;
   assign int_h2c_gpio_8_gpio_16 = h2c_gpio_8_gpio_16_f;
   assign int_h2c_gpio_8_gpio_15 = h2c_gpio_8_gpio_15_f;
   assign int_h2c_gpio_8_gpio_14 = h2c_gpio_8_gpio_14_f;
   assign int_h2c_gpio_8_gpio_13 = h2c_gpio_8_gpio_13_f;
   assign int_h2c_gpio_8_gpio_12 = h2c_gpio_8_gpio_12_f;
   assign int_h2c_gpio_8_gpio_11 = h2c_gpio_8_gpio_11_f;
   assign int_h2c_gpio_8_gpio_10 = h2c_gpio_8_gpio_10_f;
   assign int_h2c_gpio_8_gpio_9 = h2c_gpio_8_gpio_9_f;
   assign int_h2c_gpio_8_gpio_8 = h2c_gpio_8_gpio_8_f;
   assign int_h2c_gpio_8_gpio_7 = h2c_gpio_8_gpio_7_f;
   assign int_h2c_gpio_8_gpio_6 = h2c_gpio_8_gpio_6_f;
   assign int_h2c_gpio_8_gpio_5 = h2c_gpio_8_gpio_5_f;
   assign int_h2c_gpio_8_gpio_4 = h2c_gpio_8_gpio_4_f;
   assign int_h2c_gpio_8_gpio_3 = h2c_gpio_8_gpio_3_f;
   assign int_h2c_gpio_8_gpio_2 = h2c_gpio_8_gpio_2_f;
   assign int_h2c_gpio_8_gpio_1 = h2c_gpio_8_gpio_1_f;
   assign int_h2c_gpio_8_gpio_0 = h2c_gpio_8_gpio_0_f;
   assign int_h2c_gpio_9_gpio_31 = h2c_gpio_9_gpio_31_f;
   assign int_h2c_gpio_9_gpio_30 = h2c_gpio_9_gpio_30_f;
   assign int_h2c_gpio_9_gpio_29 = h2c_gpio_9_gpio_29_f;
   assign int_h2c_gpio_9_gpio_28 = h2c_gpio_9_gpio_28_f;
   assign int_h2c_gpio_9_gpio_27 = h2c_gpio_9_gpio_27_f;
   assign int_h2c_gpio_9_gpio_26 = h2c_gpio_9_gpio_26_f;
   assign int_h2c_gpio_9_gpio_25 = h2c_gpio_9_gpio_25_f;
   assign int_h2c_gpio_9_gpio_24 = h2c_gpio_9_gpio_24_f;
   assign int_h2c_gpio_9_gpio_23 = h2c_gpio_9_gpio_23_f;
   assign int_h2c_gpio_9_gpio_22 = h2c_gpio_9_gpio_22_f;
   assign int_h2c_gpio_9_gpio_21 = h2c_gpio_9_gpio_21_f;
   assign int_h2c_gpio_9_gpio_20 = h2c_gpio_9_gpio_20_f;
   assign int_h2c_gpio_9_gpio_19 = h2c_gpio_9_gpio_19_f;
   assign int_h2c_gpio_9_gpio_18 = h2c_gpio_9_gpio_18_f;
   assign int_h2c_gpio_9_gpio_17 = h2c_gpio_9_gpio_17_f;
   assign int_h2c_gpio_9_gpio_16 = h2c_gpio_9_gpio_16_f;
   assign int_h2c_gpio_9_gpio_15 = h2c_gpio_9_gpio_15_f;
   assign int_h2c_gpio_9_gpio_14 = h2c_gpio_9_gpio_14_f;
   assign int_h2c_gpio_9_gpio_13 = h2c_gpio_9_gpio_13_f;
   assign int_h2c_gpio_9_gpio_12 = h2c_gpio_9_gpio_12_f;
   assign int_h2c_gpio_9_gpio_11 = h2c_gpio_9_gpio_11_f;
   assign int_h2c_gpio_9_gpio_10 = h2c_gpio_9_gpio_10_f;
   assign int_h2c_gpio_9_gpio_9 = h2c_gpio_9_gpio_9_f;
   assign int_h2c_gpio_9_gpio_8 = h2c_gpio_9_gpio_8_f;
   assign int_h2c_gpio_9_gpio_7 = h2c_gpio_9_gpio_7_f;
   assign int_h2c_gpio_9_gpio_6 = h2c_gpio_9_gpio_6_f;
   assign int_h2c_gpio_9_gpio_5 = h2c_gpio_9_gpio_5_f;
   assign int_h2c_gpio_9_gpio_4 = h2c_gpio_9_gpio_4_f;
   assign int_h2c_gpio_9_gpio_3 = h2c_gpio_9_gpio_3_f;
   assign int_h2c_gpio_9_gpio_2 = h2c_gpio_9_gpio_2_f;
   assign int_h2c_gpio_9_gpio_1 = h2c_gpio_9_gpio_1_f;
   assign int_h2c_gpio_9_gpio_0 = h2c_gpio_9_gpio_0_f;
   assign int_h2c_gpio_10_gpio_31 = h2c_gpio_10_gpio_31_f;
   assign int_h2c_gpio_10_gpio_30 = h2c_gpio_10_gpio_30_f;
   assign int_h2c_gpio_10_gpio_29 = h2c_gpio_10_gpio_29_f;
   assign int_h2c_gpio_10_gpio_28 = h2c_gpio_10_gpio_28_f;
   assign int_h2c_gpio_10_gpio_27 = h2c_gpio_10_gpio_27_f;
   assign int_h2c_gpio_10_gpio_26 = h2c_gpio_10_gpio_26_f;
   assign int_h2c_gpio_10_gpio_25 = h2c_gpio_10_gpio_25_f;
   assign int_h2c_gpio_10_gpio_24 = h2c_gpio_10_gpio_24_f;
   assign int_h2c_gpio_10_gpio_23 = h2c_gpio_10_gpio_23_f;
   assign int_h2c_gpio_10_gpio_22 = h2c_gpio_10_gpio_22_f;
   assign int_h2c_gpio_10_gpio_21 = h2c_gpio_10_gpio_21_f;
   assign int_h2c_gpio_10_gpio_20 = h2c_gpio_10_gpio_20_f;
   assign int_h2c_gpio_10_gpio_19 = h2c_gpio_10_gpio_19_f;
   assign int_h2c_gpio_10_gpio_18 = h2c_gpio_10_gpio_18_f;
   assign int_h2c_gpio_10_gpio_17 = h2c_gpio_10_gpio_17_f;
   assign int_h2c_gpio_10_gpio_16 = h2c_gpio_10_gpio_16_f;
   assign int_h2c_gpio_10_gpio_15 = h2c_gpio_10_gpio_15_f;
   assign int_h2c_gpio_10_gpio_14 = h2c_gpio_10_gpio_14_f;
   assign int_h2c_gpio_10_gpio_13 = h2c_gpio_10_gpio_13_f;
   assign int_h2c_gpio_10_gpio_12 = h2c_gpio_10_gpio_12_f;
   assign int_h2c_gpio_10_gpio_11 = h2c_gpio_10_gpio_11_f;
   assign int_h2c_gpio_10_gpio_10 = h2c_gpio_10_gpio_10_f;
   assign int_h2c_gpio_10_gpio_9 = h2c_gpio_10_gpio_9_f;
   assign int_h2c_gpio_10_gpio_8 = h2c_gpio_10_gpio_8_f;
   assign int_h2c_gpio_10_gpio_7 = h2c_gpio_10_gpio_7_f;
   assign int_h2c_gpio_10_gpio_6 = h2c_gpio_10_gpio_6_f;
   assign int_h2c_gpio_10_gpio_5 = h2c_gpio_10_gpio_5_f;
   assign int_h2c_gpio_10_gpio_4 = h2c_gpio_10_gpio_4_f;
   assign int_h2c_gpio_10_gpio_3 = h2c_gpio_10_gpio_3_f;
   assign int_h2c_gpio_10_gpio_2 = h2c_gpio_10_gpio_2_f;
   assign int_h2c_gpio_10_gpio_1 = h2c_gpio_10_gpio_1_f;
   assign int_h2c_gpio_10_gpio_0 = h2c_gpio_10_gpio_0_f;
   assign int_h2c_gpio_11_gpio_31 = h2c_gpio_11_gpio_31_f;
   assign int_h2c_gpio_11_gpio_30 = h2c_gpio_11_gpio_30_f;
   assign int_h2c_gpio_11_gpio_29 = h2c_gpio_11_gpio_29_f;
   assign int_h2c_gpio_11_gpio_28 = h2c_gpio_11_gpio_28_f;
   assign int_h2c_gpio_11_gpio_27 = h2c_gpio_11_gpio_27_f;
   assign int_h2c_gpio_11_gpio_26 = h2c_gpio_11_gpio_26_f;
   assign int_h2c_gpio_11_gpio_25 = h2c_gpio_11_gpio_25_f;
   assign int_h2c_gpio_11_gpio_24 = h2c_gpio_11_gpio_24_f;
   assign int_h2c_gpio_11_gpio_23 = h2c_gpio_11_gpio_23_f;
   assign int_h2c_gpio_11_gpio_22 = h2c_gpio_11_gpio_22_f;
   assign int_h2c_gpio_11_gpio_21 = h2c_gpio_11_gpio_21_f;
   assign int_h2c_gpio_11_gpio_20 = h2c_gpio_11_gpio_20_f;
   assign int_h2c_gpio_11_gpio_19 = h2c_gpio_11_gpio_19_f;
   assign int_h2c_gpio_11_gpio_18 = h2c_gpio_11_gpio_18_f;
   assign int_h2c_gpio_11_gpio_17 = h2c_gpio_11_gpio_17_f;
   assign int_h2c_gpio_11_gpio_16 = h2c_gpio_11_gpio_16_f;
   assign int_h2c_gpio_11_gpio_15 = h2c_gpio_11_gpio_15_f;
   assign int_h2c_gpio_11_gpio_14 = h2c_gpio_11_gpio_14_f;
   assign int_h2c_gpio_11_gpio_13 = h2c_gpio_11_gpio_13_f;
   assign int_h2c_gpio_11_gpio_12 = h2c_gpio_11_gpio_12_f;
   assign int_h2c_gpio_11_gpio_11 = h2c_gpio_11_gpio_11_f;
   assign int_h2c_gpio_11_gpio_10 = h2c_gpio_11_gpio_10_f;
   assign int_h2c_gpio_11_gpio_9 = h2c_gpio_11_gpio_9_f;
   assign int_h2c_gpio_11_gpio_8 = h2c_gpio_11_gpio_8_f;
   assign int_h2c_gpio_11_gpio_7 = h2c_gpio_11_gpio_7_f;
   assign int_h2c_gpio_11_gpio_6 = h2c_gpio_11_gpio_6_f;
   assign int_h2c_gpio_11_gpio_5 = h2c_gpio_11_gpio_5_f;
   assign int_h2c_gpio_11_gpio_4 = h2c_gpio_11_gpio_4_f;
   assign int_h2c_gpio_11_gpio_3 = h2c_gpio_11_gpio_3_f;
   assign int_h2c_gpio_11_gpio_2 = h2c_gpio_11_gpio_2_f;
   assign int_h2c_gpio_11_gpio_1 = h2c_gpio_11_gpio_1_f;
   assign int_h2c_gpio_11_gpio_0 = h2c_gpio_11_gpio_0_f;
   assign int_h2c_gpio_12_gpio_31 = h2c_gpio_12_gpio_31_f;
   assign int_h2c_gpio_12_gpio_30 = h2c_gpio_12_gpio_30_f;
   assign int_h2c_gpio_12_gpio_29 = h2c_gpio_12_gpio_29_f;
   assign int_h2c_gpio_12_gpio_28 = h2c_gpio_12_gpio_28_f;
   assign int_h2c_gpio_12_gpio_27 = h2c_gpio_12_gpio_27_f;
   assign int_h2c_gpio_12_gpio_26 = h2c_gpio_12_gpio_26_f;
   assign int_h2c_gpio_12_gpio_25 = h2c_gpio_12_gpio_25_f;
   assign int_h2c_gpio_12_gpio_24 = h2c_gpio_12_gpio_24_f;
   assign int_h2c_gpio_12_gpio_23 = h2c_gpio_12_gpio_23_f;
   assign int_h2c_gpio_12_gpio_22 = h2c_gpio_12_gpio_22_f;
   assign int_h2c_gpio_12_gpio_21 = h2c_gpio_12_gpio_21_f;
   assign int_h2c_gpio_12_gpio_20 = h2c_gpio_12_gpio_20_f;
   assign int_h2c_gpio_12_gpio_19 = h2c_gpio_12_gpio_19_f;
   assign int_h2c_gpio_12_gpio_18 = h2c_gpio_12_gpio_18_f;
   assign int_h2c_gpio_12_gpio_17 = h2c_gpio_12_gpio_17_f;
   assign int_h2c_gpio_12_gpio_16 = h2c_gpio_12_gpio_16_f;
   assign int_h2c_gpio_12_gpio_15 = h2c_gpio_12_gpio_15_f;
   assign int_h2c_gpio_12_gpio_14 = h2c_gpio_12_gpio_14_f;
   assign int_h2c_gpio_12_gpio_13 = h2c_gpio_12_gpio_13_f;
   assign int_h2c_gpio_12_gpio_12 = h2c_gpio_12_gpio_12_f;
   assign int_h2c_gpio_12_gpio_11 = h2c_gpio_12_gpio_11_f;
   assign int_h2c_gpio_12_gpio_10 = h2c_gpio_12_gpio_10_f;
   assign int_h2c_gpio_12_gpio_9 = h2c_gpio_12_gpio_9_f;
   assign int_h2c_gpio_12_gpio_8 = h2c_gpio_12_gpio_8_f;
   assign int_h2c_gpio_12_gpio_7 = h2c_gpio_12_gpio_7_f;
   assign int_h2c_gpio_12_gpio_6 = h2c_gpio_12_gpio_6_f;
   assign int_h2c_gpio_12_gpio_5 = h2c_gpio_12_gpio_5_f;
   assign int_h2c_gpio_12_gpio_4 = h2c_gpio_12_gpio_4_f;
   assign int_h2c_gpio_12_gpio_3 = h2c_gpio_12_gpio_3_f;
   assign int_h2c_gpio_12_gpio_2 = h2c_gpio_12_gpio_2_f;
   assign int_h2c_gpio_12_gpio_1 = h2c_gpio_12_gpio_1_f;
   assign int_h2c_gpio_12_gpio_0 = h2c_gpio_12_gpio_0_f;
   assign int_h2c_gpio_13_gpio_31 = h2c_gpio_13_gpio_31_f;
   assign int_h2c_gpio_13_gpio_30 = h2c_gpio_13_gpio_30_f;
   assign int_h2c_gpio_13_gpio_29 = h2c_gpio_13_gpio_29_f;
   assign int_h2c_gpio_13_gpio_28 = h2c_gpio_13_gpio_28_f;
   assign int_h2c_gpio_13_gpio_27 = h2c_gpio_13_gpio_27_f;
   assign int_h2c_gpio_13_gpio_26 = h2c_gpio_13_gpio_26_f;
   assign int_h2c_gpio_13_gpio_25 = h2c_gpio_13_gpio_25_f;
   assign int_h2c_gpio_13_gpio_24 = h2c_gpio_13_gpio_24_f;
   assign int_h2c_gpio_13_gpio_23 = h2c_gpio_13_gpio_23_f;
   assign int_h2c_gpio_13_gpio_22 = h2c_gpio_13_gpio_22_f;
   assign int_h2c_gpio_13_gpio_21 = h2c_gpio_13_gpio_21_f;
   assign int_h2c_gpio_13_gpio_20 = h2c_gpio_13_gpio_20_f;
   assign int_h2c_gpio_13_gpio_19 = h2c_gpio_13_gpio_19_f;
   assign int_h2c_gpio_13_gpio_18 = h2c_gpio_13_gpio_18_f;
   assign int_h2c_gpio_13_gpio_17 = h2c_gpio_13_gpio_17_f;
   assign int_h2c_gpio_13_gpio_16 = h2c_gpio_13_gpio_16_f;
   assign int_h2c_gpio_13_gpio_15 = h2c_gpio_13_gpio_15_f;
   assign int_h2c_gpio_13_gpio_14 = h2c_gpio_13_gpio_14_f;
   assign int_h2c_gpio_13_gpio_13 = h2c_gpio_13_gpio_13_f;
   assign int_h2c_gpio_13_gpio_12 = h2c_gpio_13_gpio_12_f;
   assign int_h2c_gpio_13_gpio_11 = h2c_gpio_13_gpio_11_f;
   assign int_h2c_gpio_13_gpio_10 = h2c_gpio_13_gpio_10_f;
   assign int_h2c_gpio_13_gpio_9 = h2c_gpio_13_gpio_9_f;
   assign int_h2c_gpio_13_gpio_8 = h2c_gpio_13_gpio_8_f;
   assign int_h2c_gpio_13_gpio_7 = h2c_gpio_13_gpio_7_f;
   assign int_h2c_gpio_13_gpio_6 = h2c_gpio_13_gpio_6_f;
   assign int_h2c_gpio_13_gpio_5 = h2c_gpio_13_gpio_5_f;
   assign int_h2c_gpio_13_gpio_4 = h2c_gpio_13_gpio_4_f;
   assign int_h2c_gpio_13_gpio_3 = h2c_gpio_13_gpio_3_f;
   assign int_h2c_gpio_13_gpio_2 = h2c_gpio_13_gpio_2_f;
   assign int_h2c_gpio_13_gpio_1 = h2c_gpio_13_gpio_1_f;
   assign int_h2c_gpio_13_gpio_0 = h2c_gpio_13_gpio_0_f;
   assign int_h2c_gpio_14_gpio_31 = h2c_gpio_14_gpio_31_f;
   assign int_h2c_gpio_14_gpio_30 = h2c_gpio_14_gpio_30_f;
   assign int_h2c_gpio_14_gpio_29 = h2c_gpio_14_gpio_29_f;
   assign int_h2c_gpio_14_gpio_28 = h2c_gpio_14_gpio_28_f;
   assign int_h2c_gpio_14_gpio_27 = h2c_gpio_14_gpio_27_f;
   assign int_h2c_gpio_14_gpio_26 = h2c_gpio_14_gpio_26_f;
   assign int_h2c_gpio_14_gpio_25 = h2c_gpio_14_gpio_25_f;
   assign int_h2c_gpio_14_gpio_24 = h2c_gpio_14_gpio_24_f;
   assign int_h2c_gpio_14_gpio_23 = h2c_gpio_14_gpio_23_f;
   assign int_h2c_gpio_14_gpio_22 = h2c_gpio_14_gpio_22_f;
   assign int_h2c_gpio_14_gpio_21 = h2c_gpio_14_gpio_21_f;
   assign int_h2c_gpio_14_gpio_20 = h2c_gpio_14_gpio_20_f;
   assign int_h2c_gpio_14_gpio_19 = h2c_gpio_14_gpio_19_f;
   assign int_h2c_gpio_14_gpio_18 = h2c_gpio_14_gpio_18_f;
   assign int_h2c_gpio_14_gpio_17 = h2c_gpio_14_gpio_17_f;
   assign int_h2c_gpio_14_gpio_16 = h2c_gpio_14_gpio_16_f;
   assign int_h2c_gpio_14_gpio_15 = h2c_gpio_14_gpio_15_f;
   assign int_h2c_gpio_14_gpio_14 = h2c_gpio_14_gpio_14_f;
   assign int_h2c_gpio_14_gpio_13 = h2c_gpio_14_gpio_13_f;
   assign int_h2c_gpio_14_gpio_12 = h2c_gpio_14_gpio_12_f;
   assign int_h2c_gpio_14_gpio_11 = h2c_gpio_14_gpio_11_f;
   assign int_h2c_gpio_14_gpio_10 = h2c_gpio_14_gpio_10_f;
   assign int_h2c_gpio_14_gpio_9 = h2c_gpio_14_gpio_9_f;
   assign int_h2c_gpio_14_gpio_8 = h2c_gpio_14_gpio_8_f;
   assign int_h2c_gpio_14_gpio_7 = h2c_gpio_14_gpio_7_f;
   assign int_h2c_gpio_14_gpio_6 = h2c_gpio_14_gpio_6_f;
   assign int_h2c_gpio_14_gpio_5 = h2c_gpio_14_gpio_5_f;
   assign int_h2c_gpio_14_gpio_4 = h2c_gpio_14_gpio_4_f;
   assign int_h2c_gpio_14_gpio_3 = h2c_gpio_14_gpio_3_f;
   assign int_h2c_gpio_14_gpio_2 = h2c_gpio_14_gpio_2_f;
   assign int_h2c_gpio_14_gpio_1 = h2c_gpio_14_gpio_1_f;
   assign int_h2c_gpio_14_gpio_0 = h2c_gpio_14_gpio_0_f;
   assign int_h2c_gpio_15_gpio_31 = h2c_gpio_15_gpio_31_f;
   assign int_h2c_gpio_15_gpio_30 = h2c_gpio_15_gpio_30_f;
   assign int_h2c_gpio_15_gpio_29 = h2c_gpio_15_gpio_29_f;
   assign int_h2c_gpio_15_gpio_28 = h2c_gpio_15_gpio_28_f;
   assign int_h2c_gpio_15_gpio_27 = h2c_gpio_15_gpio_27_f;
   assign int_h2c_gpio_15_gpio_26 = h2c_gpio_15_gpio_26_f;
   assign int_h2c_gpio_15_gpio_25 = h2c_gpio_15_gpio_25_f;
   assign int_h2c_gpio_15_gpio_24 = h2c_gpio_15_gpio_24_f;
   assign int_h2c_gpio_15_gpio_23 = h2c_gpio_15_gpio_23_f;
   assign int_h2c_gpio_15_gpio_22 = h2c_gpio_15_gpio_22_f;
   assign int_h2c_gpio_15_gpio_21 = h2c_gpio_15_gpio_21_f;
   assign int_h2c_gpio_15_gpio_20 = h2c_gpio_15_gpio_20_f;
   assign int_h2c_gpio_15_gpio_19 = h2c_gpio_15_gpio_19_f;
   assign int_h2c_gpio_15_gpio_18 = h2c_gpio_15_gpio_18_f;
   assign int_h2c_gpio_15_gpio_17 = h2c_gpio_15_gpio_17_f;
   assign int_h2c_gpio_15_gpio_16 = h2c_gpio_15_gpio_16_f;
   assign int_h2c_gpio_15_gpio_15 = h2c_gpio_15_gpio_15_f;
   assign int_h2c_gpio_15_gpio_14 = h2c_gpio_15_gpio_14_f;
   assign int_h2c_gpio_15_gpio_13 = h2c_gpio_15_gpio_13_f;
   assign int_h2c_gpio_15_gpio_12 = h2c_gpio_15_gpio_12_f;
   assign int_h2c_gpio_15_gpio_11 = h2c_gpio_15_gpio_11_f;
   assign int_h2c_gpio_15_gpio_10 = h2c_gpio_15_gpio_10_f;
   assign int_h2c_gpio_15_gpio_9 = h2c_gpio_15_gpio_9_f;
   assign int_h2c_gpio_15_gpio_8 = h2c_gpio_15_gpio_8_f;
   assign int_h2c_gpio_15_gpio_7 = h2c_gpio_15_gpio_7_f;
   assign int_h2c_gpio_15_gpio_6 = h2c_gpio_15_gpio_6_f;
   assign int_h2c_gpio_15_gpio_5 = h2c_gpio_15_gpio_5_f;
   assign int_h2c_gpio_15_gpio_4 = h2c_gpio_15_gpio_4_f;
   assign int_h2c_gpio_15_gpio_3 = h2c_gpio_15_gpio_3_f;
   assign int_h2c_gpio_15_gpio_2 = h2c_gpio_15_gpio_2_f;
   assign int_h2c_gpio_15_gpio_1 = h2c_gpio_15_gpio_1_f;
   assign int_h2c_gpio_15_gpio_0 = h2c_gpio_15_gpio_0_f;
   assign int_rd_resp_desc_0_data_offset_addr = rd_resp_desc_0_data_offset_addr_f;
   assign int_rd_resp_desc_0_data_size_size = rd_resp_desc_0_data_size_size_f;
   assign int_rd_resp_desc_0_data_host_addr_0_addr = rd_resp_desc_0_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_0_data_host_addr_1_addr = rd_resp_desc_0_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_0_data_host_addr_2_addr = rd_resp_desc_0_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_0_data_host_addr_3_addr = rd_resp_desc_0_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_0_resp_resp = rd_resp_desc_0_resp_resp_f;
   assign int_rd_resp_desc_0_xid_0_xid = rd_resp_desc_0_xid_0_xid_f;
   assign int_rd_resp_desc_0_xid_1_xid = rd_resp_desc_0_xid_1_xid_f;
   assign int_rd_resp_desc_0_xid_2_xid = rd_resp_desc_0_xid_2_xid_f;
   assign int_rd_resp_desc_0_xid_3_xid = rd_resp_desc_0_xid_3_xid_f;
   assign int_rd_resp_desc_0_xuser_0_xuser = rd_resp_desc_0_xuser_0_xuser_f;
   assign int_rd_resp_desc_0_xuser_1_xuser = rd_resp_desc_0_xuser_1_xuser_f;
   assign int_rd_resp_desc_0_xuser_2_xuser = rd_resp_desc_0_xuser_2_xuser_f;
   assign int_rd_resp_desc_0_xuser_3_xuser = rd_resp_desc_0_xuser_3_xuser_f;
   assign int_rd_resp_desc_0_xuser_4_xuser = rd_resp_desc_0_xuser_4_xuser_f;
   assign int_rd_resp_desc_0_xuser_5_xuser = rd_resp_desc_0_xuser_5_xuser_f;
   assign int_rd_resp_desc_0_xuser_6_xuser = rd_resp_desc_0_xuser_6_xuser_f;
   assign int_rd_resp_desc_0_xuser_7_xuser = rd_resp_desc_0_xuser_7_xuser_f;
   assign int_rd_resp_desc_0_xuser_8_xuser = rd_resp_desc_0_xuser_8_xuser_f;
   assign int_rd_resp_desc_0_xuser_9_xuser = rd_resp_desc_0_xuser_9_xuser_f;
   assign int_rd_resp_desc_0_xuser_10_xuser = rd_resp_desc_0_xuser_10_xuser_f;
   assign int_rd_resp_desc_0_xuser_11_xuser = rd_resp_desc_0_xuser_11_xuser_f;
   assign int_rd_resp_desc_0_xuser_12_xuser = rd_resp_desc_0_xuser_12_xuser_f;
   assign int_rd_resp_desc_0_xuser_13_xuser = rd_resp_desc_0_xuser_13_xuser_f;
   assign int_rd_resp_desc_0_xuser_14_xuser = rd_resp_desc_0_xuser_14_xuser_f;
   assign int_rd_resp_desc_0_xuser_15_xuser = rd_resp_desc_0_xuser_15_xuser_f;
   assign int_wr_req_desc_0_data_host_addr_0_addr = wr_req_desc_0_data_host_addr_0_addr_f;
   assign int_wr_req_desc_0_data_host_addr_1_addr = wr_req_desc_0_data_host_addr_1_addr_f;
   assign int_wr_req_desc_0_data_host_addr_2_addr = wr_req_desc_0_data_host_addr_2_addr_f;
   assign int_wr_req_desc_0_data_host_addr_3_addr = wr_req_desc_0_data_host_addr_3_addr_f;
   assign int_wr_req_desc_0_wstrb_host_addr_0_addr = wr_req_desc_0_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_0_wstrb_host_addr_1_addr = wr_req_desc_0_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_0_wstrb_host_addr_2_addr = wr_req_desc_0_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_0_wstrb_host_addr_3_addr = wr_req_desc_0_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_0_resp_resp = wr_resp_desc_0_resp_resp_f;
   assign int_wr_resp_desc_0_xid_0_xid = wr_resp_desc_0_xid_0_xid_f;
   assign int_wr_resp_desc_0_xid_1_xid = wr_resp_desc_0_xid_1_xid_f;
   assign int_wr_resp_desc_0_xid_2_xid = wr_resp_desc_0_xid_2_xid_f;
   assign int_wr_resp_desc_0_xid_3_xid = wr_resp_desc_0_xid_3_xid_f;
   assign int_wr_resp_desc_0_xuser_0_xuser = wr_resp_desc_0_xuser_0_xuser_f;
   assign int_wr_resp_desc_0_xuser_1_xuser = wr_resp_desc_0_xuser_1_xuser_f;
   assign int_wr_resp_desc_0_xuser_2_xuser = wr_resp_desc_0_xuser_2_xuser_f;
   assign int_wr_resp_desc_0_xuser_3_xuser = wr_resp_desc_0_xuser_3_xuser_f;
   assign int_wr_resp_desc_0_xuser_4_xuser = wr_resp_desc_0_xuser_4_xuser_f;
   assign int_wr_resp_desc_0_xuser_5_xuser = wr_resp_desc_0_xuser_5_xuser_f;
   assign int_wr_resp_desc_0_xuser_6_xuser = wr_resp_desc_0_xuser_6_xuser_f;
   assign int_wr_resp_desc_0_xuser_7_xuser = wr_resp_desc_0_xuser_7_xuser_f;
   assign int_wr_resp_desc_0_xuser_8_xuser = wr_resp_desc_0_xuser_8_xuser_f;
   assign int_wr_resp_desc_0_xuser_9_xuser = wr_resp_desc_0_xuser_9_xuser_f;
   assign int_wr_resp_desc_0_xuser_10_xuser = wr_resp_desc_0_xuser_10_xuser_f;
   assign int_wr_resp_desc_0_xuser_11_xuser = wr_resp_desc_0_xuser_11_xuser_f;
   assign int_wr_resp_desc_0_xuser_12_xuser = wr_resp_desc_0_xuser_12_xuser_f;
   assign int_wr_resp_desc_0_xuser_13_xuser = wr_resp_desc_0_xuser_13_xuser_f;
   assign int_wr_resp_desc_0_xuser_14_xuser = wr_resp_desc_0_xuser_14_xuser_f;
   assign int_wr_resp_desc_0_xuser_15_xuser = wr_resp_desc_0_xuser_15_xuser_f;
   assign int_sn_req_desc_0_attr_acsnoop = sn_req_desc_0_attr_acsnoop_f;
   assign int_sn_req_desc_0_attr_acprot = sn_req_desc_0_attr_acprot_f;
   assign int_sn_req_desc_0_acaddr_0_addr = sn_req_desc_0_acaddr_0_addr_f;
   assign int_sn_req_desc_0_acaddr_1_addr = sn_req_desc_0_acaddr_1_addr_f;
   assign int_sn_req_desc_0_acaddr_2_addr = sn_req_desc_0_acaddr_2_addr_f;
   assign int_sn_req_desc_0_acaddr_3_addr = sn_req_desc_0_acaddr_3_addr_f;
   assign int_rd_resp_desc_1_data_offset_addr = rd_resp_desc_1_data_offset_addr_f;
   assign int_rd_resp_desc_1_data_size_size = rd_resp_desc_1_data_size_size_f;
   assign int_rd_resp_desc_1_data_host_addr_0_addr = rd_resp_desc_1_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_1_data_host_addr_1_addr = rd_resp_desc_1_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_1_data_host_addr_2_addr = rd_resp_desc_1_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_1_data_host_addr_3_addr = rd_resp_desc_1_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_1_resp_resp = rd_resp_desc_1_resp_resp_f;
   assign int_rd_resp_desc_1_xid_0_xid = rd_resp_desc_1_xid_0_xid_f;
   assign int_rd_resp_desc_1_xid_1_xid = rd_resp_desc_1_xid_1_xid_f;
   assign int_rd_resp_desc_1_xid_2_xid = rd_resp_desc_1_xid_2_xid_f;
   assign int_rd_resp_desc_1_xid_3_xid = rd_resp_desc_1_xid_3_xid_f;
   assign int_rd_resp_desc_1_xuser_0_xuser = rd_resp_desc_1_xuser_0_xuser_f;
   assign int_rd_resp_desc_1_xuser_1_xuser = rd_resp_desc_1_xuser_1_xuser_f;
   assign int_rd_resp_desc_1_xuser_2_xuser = rd_resp_desc_1_xuser_2_xuser_f;
   assign int_rd_resp_desc_1_xuser_3_xuser = rd_resp_desc_1_xuser_3_xuser_f;
   assign int_rd_resp_desc_1_xuser_4_xuser = rd_resp_desc_1_xuser_4_xuser_f;
   assign int_rd_resp_desc_1_xuser_5_xuser = rd_resp_desc_1_xuser_5_xuser_f;
   assign int_rd_resp_desc_1_xuser_6_xuser = rd_resp_desc_1_xuser_6_xuser_f;
   assign int_rd_resp_desc_1_xuser_7_xuser = rd_resp_desc_1_xuser_7_xuser_f;
   assign int_rd_resp_desc_1_xuser_8_xuser = rd_resp_desc_1_xuser_8_xuser_f;
   assign int_rd_resp_desc_1_xuser_9_xuser = rd_resp_desc_1_xuser_9_xuser_f;
   assign int_rd_resp_desc_1_xuser_10_xuser = rd_resp_desc_1_xuser_10_xuser_f;
   assign int_rd_resp_desc_1_xuser_11_xuser = rd_resp_desc_1_xuser_11_xuser_f;
   assign int_rd_resp_desc_1_xuser_12_xuser = rd_resp_desc_1_xuser_12_xuser_f;
   assign int_rd_resp_desc_1_xuser_13_xuser = rd_resp_desc_1_xuser_13_xuser_f;
   assign int_rd_resp_desc_1_xuser_14_xuser = rd_resp_desc_1_xuser_14_xuser_f;
   assign int_rd_resp_desc_1_xuser_15_xuser = rd_resp_desc_1_xuser_15_xuser_f;
   assign int_wr_req_desc_1_data_host_addr_0_addr = wr_req_desc_1_data_host_addr_0_addr_f;
   assign int_wr_req_desc_1_data_host_addr_1_addr = wr_req_desc_1_data_host_addr_1_addr_f;
   assign int_wr_req_desc_1_data_host_addr_2_addr = wr_req_desc_1_data_host_addr_2_addr_f;
   assign int_wr_req_desc_1_data_host_addr_3_addr = wr_req_desc_1_data_host_addr_3_addr_f;
   assign int_wr_req_desc_1_wstrb_host_addr_0_addr = wr_req_desc_1_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_1_wstrb_host_addr_1_addr = wr_req_desc_1_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_1_wstrb_host_addr_2_addr = wr_req_desc_1_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_1_wstrb_host_addr_3_addr = wr_req_desc_1_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_1_resp_resp = wr_resp_desc_1_resp_resp_f;
   assign int_wr_resp_desc_1_xid_0_xid = wr_resp_desc_1_xid_0_xid_f;
   assign int_wr_resp_desc_1_xid_1_xid = wr_resp_desc_1_xid_1_xid_f;
   assign int_wr_resp_desc_1_xid_2_xid = wr_resp_desc_1_xid_2_xid_f;
   assign int_wr_resp_desc_1_xid_3_xid = wr_resp_desc_1_xid_3_xid_f;
   assign int_wr_resp_desc_1_xuser_0_xuser = wr_resp_desc_1_xuser_0_xuser_f;
   assign int_wr_resp_desc_1_xuser_1_xuser = wr_resp_desc_1_xuser_1_xuser_f;
   assign int_wr_resp_desc_1_xuser_2_xuser = wr_resp_desc_1_xuser_2_xuser_f;
   assign int_wr_resp_desc_1_xuser_3_xuser = wr_resp_desc_1_xuser_3_xuser_f;
   assign int_wr_resp_desc_1_xuser_4_xuser = wr_resp_desc_1_xuser_4_xuser_f;
   assign int_wr_resp_desc_1_xuser_5_xuser = wr_resp_desc_1_xuser_5_xuser_f;
   assign int_wr_resp_desc_1_xuser_6_xuser = wr_resp_desc_1_xuser_6_xuser_f;
   assign int_wr_resp_desc_1_xuser_7_xuser = wr_resp_desc_1_xuser_7_xuser_f;
   assign int_wr_resp_desc_1_xuser_8_xuser = wr_resp_desc_1_xuser_8_xuser_f;
   assign int_wr_resp_desc_1_xuser_9_xuser = wr_resp_desc_1_xuser_9_xuser_f;
   assign int_wr_resp_desc_1_xuser_10_xuser = wr_resp_desc_1_xuser_10_xuser_f;
   assign int_wr_resp_desc_1_xuser_11_xuser = wr_resp_desc_1_xuser_11_xuser_f;
   assign int_wr_resp_desc_1_xuser_12_xuser = wr_resp_desc_1_xuser_12_xuser_f;
   assign int_wr_resp_desc_1_xuser_13_xuser = wr_resp_desc_1_xuser_13_xuser_f;
   assign int_wr_resp_desc_1_xuser_14_xuser = wr_resp_desc_1_xuser_14_xuser_f;
   assign int_wr_resp_desc_1_xuser_15_xuser = wr_resp_desc_1_xuser_15_xuser_f;
   assign int_sn_req_desc_1_attr_acsnoop = sn_req_desc_1_attr_acsnoop_f;
   assign int_sn_req_desc_1_attr_acprot = sn_req_desc_1_attr_acprot_f;
   assign int_sn_req_desc_1_acaddr_0_addr = sn_req_desc_1_acaddr_0_addr_f;
   assign int_sn_req_desc_1_acaddr_1_addr = sn_req_desc_1_acaddr_1_addr_f;
   assign int_sn_req_desc_1_acaddr_2_addr = sn_req_desc_1_acaddr_2_addr_f;
   assign int_sn_req_desc_1_acaddr_3_addr = sn_req_desc_1_acaddr_3_addr_f;
   assign int_rd_resp_desc_2_data_offset_addr = rd_resp_desc_2_data_offset_addr_f;
   assign int_rd_resp_desc_2_data_size_size = rd_resp_desc_2_data_size_size_f;
   assign int_rd_resp_desc_2_data_host_addr_0_addr = rd_resp_desc_2_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_2_data_host_addr_1_addr = rd_resp_desc_2_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_2_data_host_addr_2_addr = rd_resp_desc_2_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_2_data_host_addr_3_addr = rd_resp_desc_2_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_2_resp_resp = rd_resp_desc_2_resp_resp_f;
   assign int_rd_resp_desc_2_xid_0_xid = rd_resp_desc_2_xid_0_xid_f;
   assign int_rd_resp_desc_2_xid_1_xid = rd_resp_desc_2_xid_1_xid_f;
   assign int_rd_resp_desc_2_xid_2_xid = rd_resp_desc_2_xid_2_xid_f;
   assign int_rd_resp_desc_2_xid_3_xid = rd_resp_desc_2_xid_3_xid_f;
   assign int_rd_resp_desc_2_xuser_0_xuser = rd_resp_desc_2_xuser_0_xuser_f;
   assign int_rd_resp_desc_2_xuser_1_xuser = rd_resp_desc_2_xuser_1_xuser_f;
   assign int_rd_resp_desc_2_xuser_2_xuser = rd_resp_desc_2_xuser_2_xuser_f;
   assign int_rd_resp_desc_2_xuser_3_xuser = rd_resp_desc_2_xuser_3_xuser_f;
   assign int_rd_resp_desc_2_xuser_4_xuser = rd_resp_desc_2_xuser_4_xuser_f;
   assign int_rd_resp_desc_2_xuser_5_xuser = rd_resp_desc_2_xuser_5_xuser_f;
   assign int_rd_resp_desc_2_xuser_6_xuser = rd_resp_desc_2_xuser_6_xuser_f;
   assign int_rd_resp_desc_2_xuser_7_xuser = rd_resp_desc_2_xuser_7_xuser_f;
   assign int_rd_resp_desc_2_xuser_8_xuser = rd_resp_desc_2_xuser_8_xuser_f;
   assign int_rd_resp_desc_2_xuser_9_xuser = rd_resp_desc_2_xuser_9_xuser_f;
   assign int_rd_resp_desc_2_xuser_10_xuser = rd_resp_desc_2_xuser_10_xuser_f;
   assign int_rd_resp_desc_2_xuser_11_xuser = rd_resp_desc_2_xuser_11_xuser_f;
   assign int_rd_resp_desc_2_xuser_12_xuser = rd_resp_desc_2_xuser_12_xuser_f;
   assign int_rd_resp_desc_2_xuser_13_xuser = rd_resp_desc_2_xuser_13_xuser_f;
   assign int_rd_resp_desc_2_xuser_14_xuser = rd_resp_desc_2_xuser_14_xuser_f;
   assign int_rd_resp_desc_2_xuser_15_xuser = rd_resp_desc_2_xuser_15_xuser_f;
   assign int_wr_req_desc_2_data_host_addr_0_addr = wr_req_desc_2_data_host_addr_0_addr_f;
   assign int_wr_req_desc_2_data_host_addr_1_addr = wr_req_desc_2_data_host_addr_1_addr_f;
   assign int_wr_req_desc_2_data_host_addr_2_addr = wr_req_desc_2_data_host_addr_2_addr_f;
   assign int_wr_req_desc_2_data_host_addr_3_addr = wr_req_desc_2_data_host_addr_3_addr_f;
   assign int_wr_req_desc_2_wstrb_host_addr_0_addr = wr_req_desc_2_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_2_wstrb_host_addr_1_addr = wr_req_desc_2_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_2_wstrb_host_addr_2_addr = wr_req_desc_2_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_2_wstrb_host_addr_3_addr = wr_req_desc_2_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_2_resp_resp = wr_resp_desc_2_resp_resp_f;
   assign int_wr_resp_desc_2_xid_0_xid = wr_resp_desc_2_xid_0_xid_f;
   assign int_wr_resp_desc_2_xid_1_xid = wr_resp_desc_2_xid_1_xid_f;
   assign int_wr_resp_desc_2_xid_2_xid = wr_resp_desc_2_xid_2_xid_f;
   assign int_wr_resp_desc_2_xid_3_xid = wr_resp_desc_2_xid_3_xid_f;
   assign int_wr_resp_desc_2_xuser_0_xuser = wr_resp_desc_2_xuser_0_xuser_f;
   assign int_wr_resp_desc_2_xuser_1_xuser = wr_resp_desc_2_xuser_1_xuser_f;
   assign int_wr_resp_desc_2_xuser_2_xuser = wr_resp_desc_2_xuser_2_xuser_f;
   assign int_wr_resp_desc_2_xuser_3_xuser = wr_resp_desc_2_xuser_3_xuser_f;
   assign int_wr_resp_desc_2_xuser_4_xuser = wr_resp_desc_2_xuser_4_xuser_f;
   assign int_wr_resp_desc_2_xuser_5_xuser = wr_resp_desc_2_xuser_5_xuser_f;
   assign int_wr_resp_desc_2_xuser_6_xuser = wr_resp_desc_2_xuser_6_xuser_f;
   assign int_wr_resp_desc_2_xuser_7_xuser = wr_resp_desc_2_xuser_7_xuser_f;
   assign int_wr_resp_desc_2_xuser_8_xuser = wr_resp_desc_2_xuser_8_xuser_f;
   assign int_wr_resp_desc_2_xuser_9_xuser = wr_resp_desc_2_xuser_9_xuser_f;
   assign int_wr_resp_desc_2_xuser_10_xuser = wr_resp_desc_2_xuser_10_xuser_f;
   assign int_wr_resp_desc_2_xuser_11_xuser = wr_resp_desc_2_xuser_11_xuser_f;
   assign int_wr_resp_desc_2_xuser_12_xuser = wr_resp_desc_2_xuser_12_xuser_f;
   assign int_wr_resp_desc_2_xuser_13_xuser = wr_resp_desc_2_xuser_13_xuser_f;
   assign int_wr_resp_desc_2_xuser_14_xuser = wr_resp_desc_2_xuser_14_xuser_f;
   assign int_wr_resp_desc_2_xuser_15_xuser = wr_resp_desc_2_xuser_15_xuser_f;
   assign int_sn_req_desc_2_attr_acsnoop = sn_req_desc_2_attr_acsnoop_f;
   assign int_sn_req_desc_2_attr_acprot = sn_req_desc_2_attr_acprot_f;
   assign int_sn_req_desc_2_acaddr_0_addr = sn_req_desc_2_acaddr_0_addr_f;
   assign int_sn_req_desc_2_acaddr_1_addr = sn_req_desc_2_acaddr_1_addr_f;
   assign int_sn_req_desc_2_acaddr_2_addr = sn_req_desc_2_acaddr_2_addr_f;
   assign int_sn_req_desc_2_acaddr_3_addr = sn_req_desc_2_acaddr_3_addr_f;
   assign int_rd_resp_desc_3_data_offset_addr = rd_resp_desc_3_data_offset_addr_f;
   assign int_rd_resp_desc_3_data_size_size = rd_resp_desc_3_data_size_size_f;
   assign int_rd_resp_desc_3_data_host_addr_0_addr = rd_resp_desc_3_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_3_data_host_addr_1_addr = rd_resp_desc_3_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_3_data_host_addr_2_addr = rd_resp_desc_3_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_3_data_host_addr_3_addr = rd_resp_desc_3_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_3_resp_resp = rd_resp_desc_3_resp_resp_f;
   assign int_rd_resp_desc_3_xid_0_xid = rd_resp_desc_3_xid_0_xid_f;
   assign int_rd_resp_desc_3_xid_1_xid = rd_resp_desc_3_xid_1_xid_f;
   assign int_rd_resp_desc_3_xid_2_xid = rd_resp_desc_3_xid_2_xid_f;
   assign int_rd_resp_desc_3_xid_3_xid = rd_resp_desc_3_xid_3_xid_f;
   assign int_rd_resp_desc_3_xuser_0_xuser = rd_resp_desc_3_xuser_0_xuser_f;
   assign int_rd_resp_desc_3_xuser_1_xuser = rd_resp_desc_3_xuser_1_xuser_f;
   assign int_rd_resp_desc_3_xuser_2_xuser = rd_resp_desc_3_xuser_2_xuser_f;
   assign int_rd_resp_desc_3_xuser_3_xuser = rd_resp_desc_3_xuser_3_xuser_f;
   assign int_rd_resp_desc_3_xuser_4_xuser = rd_resp_desc_3_xuser_4_xuser_f;
   assign int_rd_resp_desc_3_xuser_5_xuser = rd_resp_desc_3_xuser_5_xuser_f;
   assign int_rd_resp_desc_3_xuser_6_xuser = rd_resp_desc_3_xuser_6_xuser_f;
   assign int_rd_resp_desc_3_xuser_7_xuser = rd_resp_desc_3_xuser_7_xuser_f;
   assign int_rd_resp_desc_3_xuser_8_xuser = rd_resp_desc_3_xuser_8_xuser_f;
   assign int_rd_resp_desc_3_xuser_9_xuser = rd_resp_desc_3_xuser_9_xuser_f;
   assign int_rd_resp_desc_3_xuser_10_xuser = rd_resp_desc_3_xuser_10_xuser_f;
   assign int_rd_resp_desc_3_xuser_11_xuser = rd_resp_desc_3_xuser_11_xuser_f;
   assign int_rd_resp_desc_3_xuser_12_xuser = rd_resp_desc_3_xuser_12_xuser_f;
   assign int_rd_resp_desc_3_xuser_13_xuser = rd_resp_desc_3_xuser_13_xuser_f;
   assign int_rd_resp_desc_3_xuser_14_xuser = rd_resp_desc_3_xuser_14_xuser_f;
   assign int_rd_resp_desc_3_xuser_15_xuser = rd_resp_desc_3_xuser_15_xuser_f;
   assign int_wr_req_desc_3_data_host_addr_0_addr = wr_req_desc_3_data_host_addr_0_addr_f;
   assign int_wr_req_desc_3_data_host_addr_1_addr = wr_req_desc_3_data_host_addr_1_addr_f;
   assign int_wr_req_desc_3_data_host_addr_2_addr = wr_req_desc_3_data_host_addr_2_addr_f;
   assign int_wr_req_desc_3_data_host_addr_3_addr = wr_req_desc_3_data_host_addr_3_addr_f;
   assign int_wr_req_desc_3_wstrb_host_addr_0_addr = wr_req_desc_3_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_3_wstrb_host_addr_1_addr = wr_req_desc_3_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_3_wstrb_host_addr_2_addr = wr_req_desc_3_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_3_wstrb_host_addr_3_addr = wr_req_desc_3_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_3_resp_resp = wr_resp_desc_3_resp_resp_f;
   assign int_wr_resp_desc_3_xid_0_xid = wr_resp_desc_3_xid_0_xid_f;
   assign int_wr_resp_desc_3_xid_1_xid = wr_resp_desc_3_xid_1_xid_f;
   assign int_wr_resp_desc_3_xid_2_xid = wr_resp_desc_3_xid_2_xid_f;
   assign int_wr_resp_desc_3_xid_3_xid = wr_resp_desc_3_xid_3_xid_f;
   assign int_wr_resp_desc_3_xuser_0_xuser = wr_resp_desc_3_xuser_0_xuser_f;
   assign int_wr_resp_desc_3_xuser_1_xuser = wr_resp_desc_3_xuser_1_xuser_f;
   assign int_wr_resp_desc_3_xuser_2_xuser = wr_resp_desc_3_xuser_2_xuser_f;
   assign int_wr_resp_desc_3_xuser_3_xuser = wr_resp_desc_3_xuser_3_xuser_f;
   assign int_wr_resp_desc_3_xuser_4_xuser = wr_resp_desc_3_xuser_4_xuser_f;
   assign int_wr_resp_desc_3_xuser_5_xuser = wr_resp_desc_3_xuser_5_xuser_f;
   assign int_wr_resp_desc_3_xuser_6_xuser = wr_resp_desc_3_xuser_6_xuser_f;
   assign int_wr_resp_desc_3_xuser_7_xuser = wr_resp_desc_3_xuser_7_xuser_f;
   assign int_wr_resp_desc_3_xuser_8_xuser = wr_resp_desc_3_xuser_8_xuser_f;
   assign int_wr_resp_desc_3_xuser_9_xuser = wr_resp_desc_3_xuser_9_xuser_f;
   assign int_wr_resp_desc_3_xuser_10_xuser = wr_resp_desc_3_xuser_10_xuser_f;
   assign int_wr_resp_desc_3_xuser_11_xuser = wr_resp_desc_3_xuser_11_xuser_f;
   assign int_wr_resp_desc_3_xuser_12_xuser = wr_resp_desc_3_xuser_12_xuser_f;
   assign int_wr_resp_desc_3_xuser_13_xuser = wr_resp_desc_3_xuser_13_xuser_f;
   assign int_wr_resp_desc_3_xuser_14_xuser = wr_resp_desc_3_xuser_14_xuser_f;
   assign int_wr_resp_desc_3_xuser_15_xuser = wr_resp_desc_3_xuser_15_xuser_f;
   assign int_sn_req_desc_3_attr_acsnoop = sn_req_desc_3_attr_acsnoop_f;
   assign int_sn_req_desc_3_attr_acprot = sn_req_desc_3_attr_acprot_f;
   assign int_sn_req_desc_3_acaddr_0_addr = sn_req_desc_3_acaddr_0_addr_f;
   assign int_sn_req_desc_3_acaddr_1_addr = sn_req_desc_3_acaddr_1_addr_f;
   assign int_sn_req_desc_3_acaddr_2_addr = sn_req_desc_3_acaddr_2_addr_f;
   assign int_sn_req_desc_3_acaddr_3_addr = sn_req_desc_3_acaddr_3_addr_f;
   assign int_rd_resp_desc_4_data_offset_addr = rd_resp_desc_4_data_offset_addr_f;
   assign int_rd_resp_desc_4_data_size_size = rd_resp_desc_4_data_size_size_f;
   assign int_rd_resp_desc_4_data_host_addr_0_addr = rd_resp_desc_4_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_4_data_host_addr_1_addr = rd_resp_desc_4_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_4_data_host_addr_2_addr = rd_resp_desc_4_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_4_data_host_addr_3_addr = rd_resp_desc_4_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_4_resp_resp = rd_resp_desc_4_resp_resp_f;
   assign int_rd_resp_desc_4_xid_0_xid = rd_resp_desc_4_xid_0_xid_f;
   assign int_rd_resp_desc_4_xid_1_xid = rd_resp_desc_4_xid_1_xid_f;
   assign int_rd_resp_desc_4_xid_2_xid = rd_resp_desc_4_xid_2_xid_f;
   assign int_rd_resp_desc_4_xid_3_xid = rd_resp_desc_4_xid_3_xid_f;
   assign int_rd_resp_desc_4_xuser_0_xuser = rd_resp_desc_4_xuser_0_xuser_f;
   assign int_rd_resp_desc_4_xuser_1_xuser = rd_resp_desc_4_xuser_1_xuser_f;
   assign int_rd_resp_desc_4_xuser_2_xuser = rd_resp_desc_4_xuser_2_xuser_f;
   assign int_rd_resp_desc_4_xuser_3_xuser = rd_resp_desc_4_xuser_3_xuser_f;
   assign int_rd_resp_desc_4_xuser_4_xuser = rd_resp_desc_4_xuser_4_xuser_f;
   assign int_rd_resp_desc_4_xuser_5_xuser = rd_resp_desc_4_xuser_5_xuser_f;
   assign int_rd_resp_desc_4_xuser_6_xuser = rd_resp_desc_4_xuser_6_xuser_f;
   assign int_rd_resp_desc_4_xuser_7_xuser = rd_resp_desc_4_xuser_7_xuser_f;
   assign int_rd_resp_desc_4_xuser_8_xuser = rd_resp_desc_4_xuser_8_xuser_f;
   assign int_rd_resp_desc_4_xuser_9_xuser = rd_resp_desc_4_xuser_9_xuser_f;
   assign int_rd_resp_desc_4_xuser_10_xuser = rd_resp_desc_4_xuser_10_xuser_f;
   assign int_rd_resp_desc_4_xuser_11_xuser = rd_resp_desc_4_xuser_11_xuser_f;
   assign int_rd_resp_desc_4_xuser_12_xuser = rd_resp_desc_4_xuser_12_xuser_f;
   assign int_rd_resp_desc_4_xuser_13_xuser = rd_resp_desc_4_xuser_13_xuser_f;
   assign int_rd_resp_desc_4_xuser_14_xuser = rd_resp_desc_4_xuser_14_xuser_f;
   assign int_rd_resp_desc_4_xuser_15_xuser = rd_resp_desc_4_xuser_15_xuser_f;
   assign int_wr_req_desc_4_data_host_addr_0_addr = wr_req_desc_4_data_host_addr_0_addr_f;
   assign int_wr_req_desc_4_data_host_addr_1_addr = wr_req_desc_4_data_host_addr_1_addr_f;
   assign int_wr_req_desc_4_data_host_addr_2_addr = wr_req_desc_4_data_host_addr_2_addr_f;
   assign int_wr_req_desc_4_data_host_addr_3_addr = wr_req_desc_4_data_host_addr_3_addr_f;
   assign int_wr_req_desc_4_wstrb_host_addr_0_addr = wr_req_desc_4_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_4_wstrb_host_addr_1_addr = wr_req_desc_4_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_4_wstrb_host_addr_2_addr = wr_req_desc_4_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_4_wstrb_host_addr_3_addr = wr_req_desc_4_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_4_resp_resp = wr_resp_desc_4_resp_resp_f;
   assign int_wr_resp_desc_4_xid_0_xid = wr_resp_desc_4_xid_0_xid_f;
   assign int_wr_resp_desc_4_xid_1_xid = wr_resp_desc_4_xid_1_xid_f;
   assign int_wr_resp_desc_4_xid_2_xid = wr_resp_desc_4_xid_2_xid_f;
   assign int_wr_resp_desc_4_xid_3_xid = wr_resp_desc_4_xid_3_xid_f;
   assign int_wr_resp_desc_4_xuser_0_xuser = wr_resp_desc_4_xuser_0_xuser_f;
   assign int_wr_resp_desc_4_xuser_1_xuser = wr_resp_desc_4_xuser_1_xuser_f;
   assign int_wr_resp_desc_4_xuser_2_xuser = wr_resp_desc_4_xuser_2_xuser_f;
   assign int_wr_resp_desc_4_xuser_3_xuser = wr_resp_desc_4_xuser_3_xuser_f;
   assign int_wr_resp_desc_4_xuser_4_xuser = wr_resp_desc_4_xuser_4_xuser_f;
   assign int_wr_resp_desc_4_xuser_5_xuser = wr_resp_desc_4_xuser_5_xuser_f;
   assign int_wr_resp_desc_4_xuser_6_xuser = wr_resp_desc_4_xuser_6_xuser_f;
   assign int_wr_resp_desc_4_xuser_7_xuser = wr_resp_desc_4_xuser_7_xuser_f;
   assign int_wr_resp_desc_4_xuser_8_xuser = wr_resp_desc_4_xuser_8_xuser_f;
   assign int_wr_resp_desc_4_xuser_9_xuser = wr_resp_desc_4_xuser_9_xuser_f;
   assign int_wr_resp_desc_4_xuser_10_xuser = wr_resp_desc_4_xuser_10_xuser_f;
   assign int_wr_resp_desc_4_xuser_11_xuser = wr_resp_desc_4_xuser_11_xuser_f;
   assign int_wr_resp_desc_4_xuser_12_xuser = wr_resp_desc_4_xuser_12_xuser_f;
   assign int_wr_resp_desc_4_xuser_13_xuser = wr_resp_desc_4_xuser_13_xuser_f;
   assign int_wr_resp_desc_4_xuser_14_xuser = wr_resp_desc_4_xuser_14_xuser_f;
   assign int_wr_resp_desc_4_xuser_15_xuser = wr_resp_desc_4_xuser_15_xuser_f;
   assign int_sn_req_desc_4_attr_acsnoop = sn_req_desc_4_attr_acsnoop_f;
   assign int_sn_req_desc_4_attr_acprot = sn_req_desc_4_attr_acprot_f;
   assign int_sn_req_desc_4_acaddr_0_addr = sn_req_desc_4_acaddr_0_addr_f;
   assign int_sn_req_desc_4_acaddr_1_addr = sn_req_desc_4_acaddr_1_addr_f;
   assign int_sn_req_desc_4_acaddr_2_addr = sn_req_desc_4_acaddr_2_addr_f;
   assign int_sn_req_desc_4_acaddr_3_addr = sn_req_desc_4_acaddr_3_addr_f;
   assign int_rd_resp_desc_5_data_offset_addr = rd_resp_desc_5_data_offset_addr_f;
   assign int_rd_resp_desc_5_data_size_size = rd_resp_desc_5_data_size_size_f;
   assign int_rd_resp_desc_5_data_host_addr_0_addr = rd_resp_desc_5_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_5_data_host_addr_1_addr = rd_resp_desc_5_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_5_data_host_addr_2_addr = rd_resp_desc_5_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_5_data_host_addr_3_addr = rd_resp_desc_5_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_5_resp_resp = rd_resp_desc_5_resp_resp_f;
   assign int_rd_resp_desc_5_xid_0_xid = rd_resp_desc_5_xid_0_xid_f;
   assign int_rd_resp_desc_5_xid_1_xid = rd_resp_desc_5_xid_1_xid_f;
   assign int_rd_resp_desc_5_xid_2_xid = rd_resp_desc_5_xid_2_xid_f;
   assign int_rd_resp_desc_5_xid_3_xid = rd_resp_desc_5_xid_3_xid_f;
   assign int_rd_resp_desc_5_xuser_0_xuser = rd_resp_desc_5_xuser_0_xuser_f;
   assign int_rd_resp_desc_5_xuser_1_xuser = rd_resp_desc_5_xuser_1_xuser_f;
   assign int_rd_resp_desc_5_xuser_2_xuser = rd_resp_desc_5_xuser_2_xuser_f;
   assign int_rd_resp_desc_5_xuser_3_xuser = rd_resp_desc_5_xuser_3_xuser_f;
   assign int_rd_resp_desc_5_xuser_4_xuser = rd_resp_desc_5_xuser_4_xuser_f;
   assign int_rd_resp_desc_5_xuser_5_xuser = rd_resp_desc_5_xuser_5_xuser_f;
   assign int_rd_resp_desc_5_xuser_6_xuser = rd_resp_desc_5_xuser_6_xuser_f;
   assign int_rd_resp_desc_5_xuser_7_xuser = rd_resp_desc_5_xuser_7_xuser_f;
   assign int_rd_resp_desc_5_xuser_8_xuser = rd_resp_desc_5_xuser_8_xuser_f;
   assign int_rd_resp_desc_5_xuser_9_xuser = rd_resp_desc_5_xuser_9_xuser_f;
   assign int_rd_resp_desc_5_xuser_10_xuser = rd_resp_desc_5_xuser_10_xuser_f;
   assign int_rd_resp_desc_5_xuser_11_xuser = rd_resp_desc_5_xuser_11_xuser_f;
   assign int_rd_resp_desc_5_xuser_12_xuser = rd_resp_desc_5_xuser_12_xuser_f;
   assign int_rd_resp_desc_5_xuser_13_xuser = rd_resp_desc_5_xuser_13_xuser_f;
   assign int_rd_resp_desc_5_xuser_14_xuser = rd_resp_desc_5_xuser_14_xuser_f;
   assign int_rd_resp_desc_5_xuser_15_xuser = rd_resp_desc_5_xuser_15_xuser_f;
   assign int_wr_req_desc_5_data_host_addr_0_addr = wr_req_desc_5_data_host_addr_0_addr_f;
   assign int_wr_req_desc_5_data_host_addr_1_addr = wr_req_desc_5_data_host_addr_1_addr_f;
   assign int_wr_req_desc_5_data_host_addr_2_addr = wr_req_desc_5_data_host_addr_2_addr_f;
   assign int_wr_req_desc_5_data_host_addr_3_addr = wr_req_desc_5_data_host_addr_3_addr_f;
   assign int_wr_req_desc_5_wstrb_host_addr_0_addr = wr_req_desc_5_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_5_wstrb_host_addr_1_addr = wr_req_desc_5_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_5_wstrb_host_addr_2_addr = wr_req_desc_5_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_5_wstrb_host_addr_3_addr = wr_req_desc_5_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_5_resp_resp = wr_resp_desc_5_resp_resp_f;
   assign int_wr_resp_desc_5_xid_0_xid = wr_resp_desc_5_xid_0_xid_f;
   assign int_wr_resp_desc_5_xid_1_xid = wr_resp_desc_5_xid_1_xid_f;
   assign int_wr_resp_desc_5_xid_2_xid = wr_resp_desc_5_xid_2_xid_f;
   assign int_wr_resp_desc_5_xid_3_xid = wr_resp_desc_5_xid_3_xid_f;
   assign int_wr_resp_desc_5_xuser_0_xuser = wr_resp_desc_5_xuser_0_xuser_f;
   assign int_wr_resp_desc_5_xuser_1_xuser = wr_resp_desc_5_xuser_1_xuser_f;
   assign int_wr_resp_desc_5_xuser_2_xuser = wr_resp_desc_5_xuser_2_xuser_f;
   assign int_wr_resp_desc_5_xuser_3_xuser = wr_resp_desc_5_xuser_3_xuser_f;
   assign int_wr_resp_desc_5_xuser_4_xuser = wr_resp_desc_5_xuser_4_xuser_f;
   assign int_wr_resp_desc_5_xuser_5_xuser = wr_resp_desc_5_xuser_5_xuser_f;
   assign int_wr_resp_desc_5_xuser_6_xuser = wr_resp_desc_5_xuser_6_xuser_f;
   assign int_wr_resp_desc_5_xuser_7_xuser = wr_resp_desc_5_xuser_7_xuser_f;
   assign int_wr_resp_desc_5_xuser_8_xuser = wr_resp_desc_5_xuser_8_xuser_f;
   assign int_wr_resp_desc_5_xuser_9_xuser = wr_resp_desc_5_xuser_9_xuser_f;
   assign int_wr_resp_desc_5_xuser_10_xuser = wr_resp_desc_5_xuser_10_xuser_f;
   assign int_wr_resp_desc_5_xuser_11_xuser = wr_resp_desc_5_xuser_11_xuser_f;
   assign int_wr_resp_desc_5_xuser_12_xuser = wr_resp_desc_5_xuser_12_xuser_f;
   assign int_wr_resp_desc_5_xuser_13_xuser = wr_resp_desc_5_xuser_13_xuser_f;
   assign int_wr_resp_desc_5_xuser_14_xuser = wr_resp_desc_5_xuser_14_xuser_f;
   assign int_wr_resp_desc_5_xuser_15_xuser = wr_resp_desc_5_xuser_15_xuser_f;
   assign int_sn_req_desc_5_attr_acsnoop = sn_req_desc_5_attr_acsnoop_f;
   assign int_sn_req_desc_5_attr_acprot = sn_req_desc_5_attr_acprot_f;
   assign int_sn_req_desc_5_acaddr_0_addr = sn_req_desc_5_acaddr_0_addr_f;
   assign int_sn_req_desc_5_acaddr_1_addr = sn_req_desc_5_acaddr_1_addr_f;
   assign int_sn_req_desc_5_acaddr_2_addr = sn_req_desc_5_acaddr_2_addr_f;
   assign int_sn_req_desc_5_acaddr_3_addr = sn_req_desc_5_acaddr_3_addr_f;
   assign int_rd_resp_desc_6_data_offset_addr = rd_resp_desc_6_data_offset_addr_f;
   assign int_rd_resp_desc_6_data_size_size = rd_resp_desc_6_data_size_size_f;
   assign int_rd_resp_desc_6_data_host_addr_0_addr = rd_resp_desc_6_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_6_data_host_addr_1_addr = rd_resp_desc_6_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_6_data_host_addr_2_addr = rd_resp_desc_6_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_6_data_host_addr_3_addr = rd_resp_desc_6_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_6_resp_resp = rd_resp_desc_6_resp_resp_f;
   assign int_rd_resp_desc_6_xid_0_xid = rd_resp_desc_6_xid_0_xid_f;
   assign int_rd_resp_desc_6_xid_1_xid = rd_resp_desc_6_xid_1_xid_f;
   assign int_rd_resp_desc_6_xid_2_xid = rd_resp_desc_6_xid_2_xid_f;
   assign int_rd_resp_desc_6_xid_3_xid = rd_resp_desc_6_xid_3_xid_f;
   assign int_rd_resp_desc_6_xuser_0_xuser = rd_resp_desc_6_xuser_0_xuser_f;
   assign int_rd_resp_desc_6_xuser_1_xuser = rd_resp_desc_6_xuser_1_xuser_f;
   assign int_rd_resp_desc_6_xuser_2_xuser = rd_resp_desc_6_xuser_2_xuser_f;
   assign int_rd_resp_desc_6_xuser_3_xuser = rd_resp_desc_6_xuser_3_xuser_f;
   assign int_rd_resp_desc_6_xuser_4_xuser = rd_resp_desc_6_xuser_4_xuser_f;
   assign int_rd_resp_desc_6_xuser_5_xuser = rd_resp_desc_6_xuser_5_xuser_f;
   assign int_rd_resp_desc_6_xuser_6_xuser = rd_resp_desc_6_xuser_6_xuser_f;
   assign int_rd_resp_desc_6_xuser_7_xuser = rd_resp_desc_6_xuser_7_xuser_f;
   assign int_rd_resp_desc_6_xuser_8_xuser = rd_resp_desc_6_xuser_8_xuser_f;
   assign int_rd_resp_desc_6_xuser_9_xuser = rd_resp_desc_6_xuser_9_xuser_f;
   assign int_rd_resp_desc_6_xuser_10_xuser = rd_resp_desc_6_xuser_10_xuser_f;
   assign int_rd_resp_desc_6_xuser_11_xuser = rd_resp_desc_6_xuser_11_xuser_f;
   assign int_rd_resp_desc_6_xuser_12_xuser = rd_resp_desc_6_xuser_12_xuser_f;
   assign int_rd_resp_desc_6_xuser_13_xuser = rd_resp_desc_6_xuser_13_xuser_f;
   assign int_rd_resp_desc_6_xuser_14_xuser = rd_resp_desc_6_xuser_14_xuser_f;
   assign int_rd_resp_desc_6_xuser_15_xuser = rd_resp_desc_6_xuser_15_xuser_f;
   assign int_wr_req_desc_6_data_host_addr_0_addr = wr_req_desc_6_data_host_addr_0_addr_f;
   assign int_wr_req_desc_6_data_host_addr_1_addr = wr_req_desc_6_data_host_addr_1_addr_f;
   assign int_wr_req_desc_6_data_host_addr_2_addr = wr_req_desc_6_data_host_addr_2_addr_f;
   assign int_wr_req_desc_6_data_host_addr_3_addr = wr_req_desc_6_data_host_addr_3_addr_f;
   assign int_wr_req_desc_6_wstrb_host_addr_0_addr = wr_req_desc_6_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_6_wstrb_host_addr_1_addr = wr_req_desc_6_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_6_wstrb_host_addr_2_addr = wr_req_desc_6_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_6_wstrb_host_addr_3_addr = wr_req_desc_6_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_6_resp_resp = wr_resp_desc_6_resp_resp_f;
   assign int_wr_resp_desc_6_xid_0_xid = wr_resp_desc_6_xid_0_xid_f;
   assign int_wr_resp_desc_6_xid_1_xid = wr_resp_desc_6_xid_1_xid_f;
   assign int_wr_resp_desc_6_xid_2_xid = wr_resp_desc_6_xid_2_xid_f;
   assign int_wr_resp_desc_6_xid_3_xid = wr_resp_desc_6_xid_3_xid_f;
   assign int_wr_resp_desc_6_xuser_0_xuser = wr_resp_desc_6_xuser_0_xuser_f;
   assign int_wr_resp_desc_6_xuser_1_xuser = wr_resp_desc_6_xuser_1_xuser_f;
   assign int_wr_resp_desc_6_xuser_2_xuser = wr_resp_desc_6_xuser_2_xuser_f;
   assign int_wr_resp_desc_6_xuser_3_xuser = wr_resp_desc_6_xuser_3_xuser_f;
   assign int_wr_resp_desc_6_xuser_4_xuser = wr_resp_desc_6_xuser_4_xuser_f;
   assign int_wr_resp_desc_6_xuser_5_xuser = wr_resp_desc_6_xuser_5_xuser_f;
   assign int_wr_resp_desc_6_xuser_6_xuser = wr_resp_desc_6_xuser_6_xuser_f;
   assign int_wr_resp_desc_6_xuser_7_xuser = wr_resp_desc_6_xuser_7_xuser_f;
   assign int_wr_resp_desc_6_xuser_8_xuser = wr_resp_desc_6_xuser_8_xuser_f;
   assign int_wr_resp_desc_6_xuser_9_xuser = wr_resp_desc_6_xuser_9_xuser_f;
   assign int_wr_resp_desc_6_xuser_10_xuser = wr_resp_desc_6_xuser_10_xuser_f;
   assign int_wr_resp_desc_6_xuser_11_xuser = wr_resp_desc_6_xuser_11_xuser_f;
   assign int_wr_resp_desc_6_xuser_12_xuser = wr_resp_desc_6_xuser_12_xuser_f;
   assign int_wr_resp_desc_6_xuser_13_xuser = wr_resp_desc_6_xuser_13_xuser_f;
   assign int_wr_resp_desc_6_xuser_14_xuser = wr_resp_desc_6_xuser_14_xuser_f;
   assign int_wr_resp_desc_6_xuser_15_xuser = wr_resp_desc_6_xuser_15_xuser_f;
   assign int_sn_req_desc_6_attr_acsnoop = sn_req_desc_6_attr_acsnoop_f;
   assign int_sn_req_desc_6_attr_acprot = sn_req_desc_6_attr_acprot_f;
   assign int_sn_req_desc_6_acaddr_0_addr = sn_req_desc_6_acaddr_0_addr_f;
   assign int_sn_req_desc_6_acaddr_1_addr = sn_req_desc_6_acaddr_1_addr_f;
   assign int_sn_req_desc_6_acaddr_2_addr = sn_req_desc_6_acaddr_2_addr_f;
   assign int_sn_req_desc_6_acaddr_3_addr = sn_req_desc_6_acaddr_3_addr_f;
   assign int_rd_resp_desc_7_data_offset_addr = rd_resp_desc_7_data_offset_addr_f;
   assign int_rd_resp_desc_7_data_size_size = rd_resp_desc_7_data_size_size_f;
   assign int_rd_resp_desc_7_data_host_addr_0_addr = rd_resp_desc_7_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_7_data_host_addr_1_addr = rd_resp_desc_7_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_7_data_host_addr_2_addr = rd_resp_desc_7_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_7_data_host_addr_3_addr = rd_resp_desc_7_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_7_resp_resp = rd_resp_desc_7_resp_resp_f;
   assign int_rd_resp_desc_7_xid_0_xid = rd_resp_desc_7_xid_0_xid_f;
   assign int_rd_resp_desc_7_xid_1_xid = rd_resp_desc_7_xid_1_xid_f;
   assign int_rd_resp_desc_7_xid_2_xid = rd_resp_desc_7_xid_2_xid_f;
   assign int_rd_resp_desc_7_xid_3_xid = rd_resp_desc_7_xid_3_xid_f;
   assign int_rd_resp_desc_7_xuser_0_xuser = rd_resp_desc_7_xuser_0_xuser_f;
   assign int_rd_resp_desc_7_xuser_1_xuser = rd_resp_desc_7_xuser_1_xuser_f;
   assign int_rd_resp_desc_7_xuser_2_xuser = rd_resp_desc_7_xuser_2_xuser_f;
   assign int_rd_resp_desc_7_xuser_3_xuser = rd_resp_desc_7_xuser_3_xuser_f;
   assign int_rd_resp_desc_7_xuser_4_xuser = rd_resp_desc_7_xuser_4_xuser_f;
   assign int_rd_resp_desc_7_xuser_5_xuser = rd_resp_desc_7_xuser_5_xuser_f;
   assign int_rd_resp_desc_7_xuser_6_xuser = rd_resp_desc_7_xuser_6_xuser_f;
   assign int_rd_resp_desc_7_xuser_7_xuser = rd_resp_desc_7_xuser_7_xuser_f;
   assign int_rd_resp_desc_7_xuser_8_xuser = rd_resp_desc_7_xuser_8_xuser_f;
   assign int_rd_resp_desc_7_xuser_9_xuser = rd_resp_desc_7_xuser_9_xuser_f;
   assign int_rd_resp_desc_7_xuser_10_xuser = rd_resp_desc_7_xuser_10_xuser_f;
   assign int_rd_resp_desc_7_xuser_11_xuser = rd_resp_desc_7_xuser_11_xuser_f;
   assign int_rd_resp_desc_7_xuser_12_xuser = rd_resp_desc_7_xuser_12_xuser_f;
   assign int_rd_resp_desc_7_xuser_13_xuser = rd_resp_desc_7_xuser_13_xuser_f;
   assign int_rd_resp_desc_7_xuser_14_xuser = rd_resp_desc_7_xuser_14_xuser_f;
   assign int_rd_resp_desc_7_xuser_15_xuser = rd_resp_desc_7_xuser_15_xuser_f;
   assign int_wr_req_desc_7_data_host_addr_0_addr = wr_req_desc_7_data_host_addr_0_addr_f;
   assign int_wr_req_desc_7_data_host_addr_1_addr = wr_req_desc_7_data_host_addr_1_addr_f;
   assign int_wr_req_desc_7_data_host_addr_2_addr = wr_req_desc_7_data_host_addr_2_addr_f;
   assign int_wr_req_desc_7_data_host_addr_3_addr = wr_req_desc_7_data_host_addr_3_addr_f;
   assign int_wr_req_desc_7_wstrb_host_addr_0_addr = wr_req_desc_7_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_7_wstrb_host_addr_1_addr = wr_req_desc_7_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_7_wstrb_host_addr_2_addr = wr_req_desc_7_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_7_wstrb_host_addr_3_addr = wr_req_desc_7_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_7_resp_resp = wr_resp_desc_7_resp_resp_f;
   assign int_wr_resp_desc_7_xid_0_xid = wr_resp_desc_7_xid_0_xid_f;
   assign int_wr_resp_desc_7_xid_1_xid = wr_resp_desc_7_xid_1_xid_f;
   assign int_wr_resp_desc_7_xid_2_xid = wr_resp_desc_7_xid_2_xid_f;
   assign int_wr_resp_desc_7_xid_3_xid = wr_resp_desc_7_xid_3_xid_f;
   assign int_wr_resp_desc_7_xuser_0_xuser = wr_resp_desc_7_xuser_0_xuser_f;
   assign int_wr_resp_desc_7_xuser_1_xuser = wr_resp_desc_7_xuser_1_xuser_f;
   assign int_wr_resp_desc_7_xuser_2_xuser = wr_resp_desc_7_xuser_2_xuser_f;
   assign int_wr_resp_desc_7_xuser_3_xuser = wr_resp_desc_7_xuser_3_xuser_f;
   assign int_wr_resp_desc_7_xuser_4_xuser = wr_resp_desc_7_xuser_4_xuser_f;
   assign int_wr_resp_desc_7_xuser_5_xuser = wr_resp_desc_7_xuser_5_xuser_f;
   assign int_wr_resp_desc_7_xuser_6_xuser = wr_resp_desc_7_xuser_6_xuser_f;
   assign int_wr_resp_desc_7_xuser_7_xuser = wr_resp_desc_7_xuser_7_xuser_f;
   assign int_wr_resp_desc_7_xuser_8_xuser = wr_resp_desc_7_xuser_8_xuser_f;
   assign int_wr_resp_desc_7_xuser_9_xuser = wr_resp_desc_7_xuser_9_xuser_f;
   assign int_wr_resp_desc_7_xuser_10_xuser = wr_resp_desc_7_xuser_10_xuser_f;
   assign int_wr_resp_desc_7_xuser_11_xuser = wr_resp_desc_7_xuser_11_xuser_f;
   assign int_wr_resp_desc_7_xuser_12_xuser = wr_resp_desc_7_xuser_12_xuser_f;
   assign int_wr_resp_desc_7_xuser_13_xuser = wr_resp_desc_7_xuser_13_xuser_f;
   assign int_wr_resp_desc_7_xuser_14_xuser = wr_resp_desc_7_xuser_14_xuser_f;
   assign int_wr_resp_desc_7_xuser_15_xuser = wr_resp_desc_7_xuser_15_xuser_f;
   assign int_sn_req_desc_7_attr_acsnoop = sn_req_desc_7_attr_acsnoop_f;
   assign int_sn_req_desc_7_attr_acprot = sn_req_desc_7_attr_acprot_f;
   assign int_sn_req_desc_7_acaddr_0_addr = sn_req_desc_7_acaddr_0_addr_f;
   assign int_sn_req_desc_7_acaddr_1_addr = sn_req_desc_7_acaddr_1_addr_f;
   assign int_sn_req_desc_7_acaddr_2_addr = sn_req_desc_7_acaddr_2_addr_f;
   assign int_sn_req_desc_7_acaddr_3_addr = sn_req_desc_7_acaddr_3_addr_f;
   assign int_rd_resp_desc_8_data_offset_addr = rd_resp_desc_8_data_offset_addr_f;
   assign int_rd_resp_desc_8_data_size_size = rd_resp_desc_8_data_size_size_f;
   assign int_rd_resp_desc_8_data_host_addr_0_addr = rd_resp_desc_8_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_8_data_host_addr_1_addr = rd_resp_desc_8_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_8_data_host_addr_2_addr = rd_resp_desc_8_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_8_data_host_addr_3_addr = rd_resp_desc_8_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_8_resp_resp = rd_resp_desc_8_resp_resp_f;
   assign int_rd_resp_desc_8_xid_0_xid = rd_resp_desc_8_xid_0_xid_f;
   assign int_rd_resp_desc_8_xid_1_xid = rd_resp_desc_8_xid_1_xid_f;
   assign int_rd_resp_desc_8_xid_2_xid = rd_resp_desc_8_xid_2_xid_f;
   assign int_rd_resp_desc_8_xid_3_xid = rd_resp_desc_8_xid_3_xid_f;
   assign int_rd_resp_desc_8_xuser_0_xuser = rd_resp_desc_8_xuser_0_xuser_f;
   assign int_rd_resp_desc_8_xuser_1_xuser = rd_resp_desc_8_xuser_1_xuser_f;
   assign int_rd_resp_desc_8_xuser_2_xuser = rd_resp_desc_8_xuser_2_xuser_f;
   assign int_rd_resp_desc_8_xuser_3_xuser = rd_resp_desc_8_xuser_3_xuser_f;
   assign int_rd_resp_desc_8_xuser_4_xuser = rd_resp_desc_8_xuser_4_xuser_f;
   assign int_rd_resp_desc_8_xuser_5_xuser = rd_resp_desc_8_xuser_5_xuser_f;
   assign int_rd_resp_desc_8_xuser_6_xuser = rd_resp_desc_8_xuser_6_xuser_f;
   assign int_rd_resp_desc_8_xuser_7_xuser = rd_resp_desc_8_xuser_7_xuser_f;
   assign int_rd_resp_desc_8_xuser_8_xuser = rd_resp_desc_8_xuser_8_xuser_f;
   assign int_rd_resp_desc_8_xuser_9_xuser = rd_resp_desc_8_xuser_9_xuser_f;
   assign int_rd_resp_desc_8_xuser_10_xuser = rd_resp_desc_8_xuser_10_xuser_f;
   assign int_rd_resp_desc_8_xuser_11_xuser = rd_resp_desc_8_xuser_11_xuser_f;
   assign int_rd_resp_desc_8_xuser_12_xuser = rd_resp_desc_8_xuser_12_xuser_f;
   assign int_rd_resp_desc_8_xuser_13_xuser = rd_resp_desc_8_xuser_13_xuser_f;
   assign int_rd_resp_desc_8_xuser_14_xuser = rd_resp_desc_8_xuser_14_xuser_f;
   assign int_rd_resp_desc_8_xuser_15_xuser = rd_resp_desc_8_xuser_15_xuser_f;
   assign int_wr_req_desc_8_data_host_addr_0_addr = wr_req_desc_8_data_host_addr_0_addr_f;
   assign int_wr_req_desc_8_data_host_addr_1_addr = wr_req_desc_8_data_host_addr_1_addr_f;
   assign int_wr_req_desc_8_data_host_addr_2_addr = wr_req_desc_8_data_host_addr_2_addr_f;
   assign int_wr_req_desc_8_data_host_addr_3_addr = wr_req_desc_8_data_host_addr_3_addr_f;
   assign int_wr_req_desc_8_wstrb_host_addr_0_addr = wr_req_desc_8_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_8_wstrb_host_addr_1_addr = wr_req_desc_8_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_8_wstrb_host_addr_2_addr = wr_req_desc_8_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_8_wstrb_host_addr_3_addr = wr_req_desc_8_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_8_resp_resp = wr_resp_desc_8_resp_resp_f;
   assign int_wr_resp_desc_8_xid_0_xid = wr_resp_desc_8_xid_0_xid_f;
   assign int_wr_resp_desc_8_xid_1_xid = wr_resp_desc_8_xid_1_xid_f;
   assign int_wr_resp_desc_8_xid_2_xid = wr_resp_desc_8_xid_2_xid_f;
   assign int_wr_resp_desc_8_xid_3_xid = wr_resp_desc_8_xid_3_xid_f;
   assign int_wr_resp_desc_8_xuser_0_xuser = wr_resp_desc_8_xuser_0_xuser_f;
   assign int_wr_resp_desc_8_xuser_1_xuser = wr_resp_desc_8_xuser_1_xuser_f;
   assign int_wr_resp_desc_8_xuser_2_xuser = wr_resp_desc_8_xuser_2_xuser_f;
   assign int_wr_resp_desc_8_xuser_3_xuser = wr_resp_desc_8_xuser_3_xuser_f;
   assign int_wr_resp_desc_8_xuser_4_xuser = wr_resp_desc_8_xuser_4_xuser_f;
   assign int_wr_resp_desc_8_xuser_5_xuser = wr_resp_desc_8_xuser_5_xuser_f;
   assign int_wr_resp_desc_8_xuser_6_xuser = wr_resp_desc_8_xuser_6_xuser_f;
   assign int_wr_resp_desc_8_xuser_7_xuser = wr_resp_desc_8_xuser_7_xuser_f;
   assign int_wr_resp_desc_8_xuser_8_xuser = wr_resp_desc_8_xuser_8_xuser_f;
   assign int_wr_resp_desc_8_xuser_9_xuser = wr_resp_desc_8_xuser_9_xuser_f;
   assign int_wr_resp_desc_8_xuser_10_xuser = wr_resp_desc_8_xuser_10_xuser_f;
   assign int_wr_resp_desc_8_xuser_11_xuser = wr_resp_desc_8_xuser_11_xuser_f;
   assign int_wr_resp_desc_8_xuser_12_xuser = wr_resp_desc_8_xuser_12_xuser_f;
   assign int_wr_resp_desc_8_xuser_13_xuser = wr_resp_desc_8_xuser_13_xuser_f;
   assign int_wr_resp_desc_8_xuser_14_xuser = wr_resp_desc_8_xuser_14_xuser_f;
   assign int_wr_resp_desc_8_xuser_15_xuser = wr_resp_desc_8_xuser_15_xuser_f;
   assign int_sn_req_desc_8_attr_acsnoop = sn_req_desc_8_attr_acsnoop_f;
   assign int_sn_req_desc_8_attr_acprot = sn_req_desc_8_attr_acprot_f;
   assign int_sn_req_desc_8_acaddr_0_addr = sn_req_desc_8_acaddr_0_addr_f;
   assign int_sn_req_desc_8_acaddr_1_addr = sn_req_desc_8_acaddr_1_addr_f;
   assign int_sn_req_desc_8_acaddr_2_addr = sn_req_desc_8_acaddr_2_addr_f;
   assign int_sn_req_desc_8_acaddr_3_addr = sn_req_desc_8_acaddr_3_addr_f;
   assign int_rd_resp_desc_9_data_offset_addr = rd_resp_desc_9_data_offset_addr_f;
   assign int_rd_resp_desc_9_data_size_size = rd_resp_desc_9_data_size_size_f;
   assign int_rd_resp_desc_9_data_host_addr_0_addr = rd_resp_desc_9_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_9_data_host_addr_1_addr = rd_resp_desc_9_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_9_data_host_addr_2_addr = rd_resp_desc_9_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_9_data_host_addr_3_addr = rd_resp_desc_9_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_9_resp_resp = rd_resp_desc_9_resp_resp_f;
   assign int_rd_resp_desc_9_xid_0_xid = rd_resp_desc_9_xid_0_xid_f;
   assign int_rd_resp_desc_9_xid_1_xid = rd_resp_desc_9_xid_1_xid_f;
   assign int_rd_resp_desc_9_xid_2_xid = rd_resp_desc_9_xid_2_xid_f;
   assign int_rd_resp_desc_9_xid_3_xid = rd_resp_desc_9_xid_3_xid_f;
   assign int_rd_resp_desc_9_xuser_0_xuser = rd_resp_desc_9_xuser_0_xuser_f;
   assign int_rd_resp_desc_9_xuser_1_xuser = rd_resp_desc_9_xuser_1_xuser_f;
   assign int_rd_resp_desc_9_xuser_2_xuser = rd_resp_desc_9_xuser_2_xuser_f;
   assign int_rd_resp_desc_9_xuser_3_xuser = rd_resp_desc_9_xuser_3_xuser_f;
   assign int_rd_resp_desc_9_xuser_4_xuser = rd_resp_desc_9_xuser_4_xuser_f;
   assign int_rd_resp_desc_9_xuser_5_xuser = rd_resp_desc_9_xuser_5_xuser_f;
   assign int_rd_resp_desc_9_xuser_6_xuser = rd_resp_desc_9_xuser_6_xuser_f;
   assign int_rd_resp_desc_9_xuser_7_xuser = rd_resp_desc_9_xuser_7_xuser_f;
   assign int_rd_resp_desc_9_xuser_8_xuser = rd_resp_desc_9_xuser_8_xuser_f;
   assign int_rd_resp_desc_9_xuser_9_xuser = rd_resp_desc_9_xuser_9_xuser_f;
   assign int_rd_resp_desc_9_xuser_10_xuser = rd_resp_desc_9_xuser_10_xuser_f;
   assign int_rd_resp_desc_9_xuser_11_xuser = rd_resp_desc_9_xuser_11_xuser_f;
   assign int_rd_resp_desc_9_xuser_12_xuser = rd_resp_desc_9_xuser_12_xuser_f;
   assign int_rd_resp_desc_9_xuser_13_xuser = rd_resp_desc_9_xuser_13_xuser_f;
   assign int_rd_resp_desc_9_xuser_14_xuser = rd_resp_desc_9_xuser_14_xuser_f;
   assign int_rd_resp_desc_9_xuser_15_xuser = rd_resp_desc_9_xuser_15_xuser_f;
   assign int_wr_req_desc_9_data_host_addr_0_addr = wr_req_desc_9_data_host_addr_0_addr_f;
   assign int_wr_req_desc_9_data_host_addr_1_addr = wr_req_desc_9_data_host_addr_1_addr_f;
   assign int_wr_req_desc_9_data_host_addr_2_addr = wr_req_desc_9_data_host_addr_2_addr_f;
   assign int_wr_req_desc_9_data_host_addr_3_addr = wr_req_desc_9_data_host_addr_3_addr_f;
   assign int_wr_req_desc_9_wstrb_host_addr_0_addr = wr_req_desc_9_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_9_wstrb_host_addr_1_addr = wr_req_desc_9_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_9_wstrb_host_addr_2_addr = wr_req_desc_9_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_9_wstrb_host_addr_3_addr = wr_req_desc_9_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_9_resp_resp = wr_resp_desc_9_resp_resp_f;
   assign int_wr_resp_desc_9_xid_0_xid = wr_resp_desc_9_xid_0_xid_f;
   assign int_wr_resp_desc_9_xid_1_xid = wr_resp_desc_9_xid_1_xid_f;
   assign int_wr_resp_desc_9_xid_2_xid = wr_resp_desc_9_xid_2_xid_f;
   assign int_wr_resp_desc_9_xid_3_xid = wr_resp_desc_9_xid_3_xid_f;
   assign int_wr_resp_desc_9_xuser_0_xuser = wr_resp_desc_9_xuser_0_xuser_f;
   assign int_wr_resp_desc_9_xuser_1_xuser = wr_resp_desc_9_xuser_1_xuser_f;
   assign int_wr_resp_desc_9_xuser_2_xuser = wr_resp_desc_9_xuser_2_xuser_f;
   assign int_wr_resp_desc_9_xuser_3_xuser = wr_resp_desc_9_xuser_3_xuser_f;
   assign int_wr_resp_desc_9_xuser_4_xuser = wr_resp_desc_9_xuser_4_xuser_f;
   assign int_wr_resp_desc_9_xuser_5_xuser = wr_resp_desc_9_xuser_5_xuser_f;
   assign int_wr_resp_desc_9_xuser_6_xuser = wr_resp_desc_9_xuser_6_xuser_f;
   assign int_wr_resp_desc_9_xuser_7_xuser = wr_resp_desc_9_xuser_7_xuser_f;
   assign int_wr_resp_desc_9_xuser_8_xuser = wr_resp_desc_9_xuser_8_xuser_f;
   assign int_wr_resp_desc_9_xuser_9_xuser = wr_resp_desc_9_xuser_9_xuser_f;
   assign int_wr_resp_desc_9_xuser_10_xuser = wr_resp_desc_9_xuser_10_xuser_f;
   assign int_wr_resp_desc_9_xuser_11_xuser = wr_resp_desc_9_xuser_11_xuser_f;
   assign int_wr_resp_desc_9_xuser_12_xuser = wr_resp_desc_9_xuser_12_xuser_f;
   assign int_wr_resp_desc_9_xuser_13_xuser = wr_resp_desc_9_xuser_13_xuser_f;
   assign int_wr_resp_desc_9_xuser_14_xuser = wr_resp_desc_9_xuser_14_xuser_f;
   assign int_wr_resp_desc_9_xuser_15_xuser = wr_resp_desc_9_xuser_15_xuser_f;
   assign int_sn_req_desc_9_attr_acsnoop = sn_req_desc_9_attr_acsnoop_f;
   assign int_sn_req_desc_9_attr_acprot = sn_req_desc_9_attr_acprot_f;
   assign int_sn_req_desc_9_acaddr_0_addr = sn_req_desc_9_acaddr_0_addr_f;
   assign int_sn_req_desc_9_acaddr_1_addr = sn_req_desc_9_acaddr_1_addr_f;
   assign int_sn_req_desc_9_acaddr_2_addr = sn_req_desc_9_acaddr_2_addr_f;
   assign int_sn_req_desc_9_acaddr_3_addr = sn_req_desc_9_acaddr_3_addr_f;
   assign int_rd_resp_desc_a_data_offset_addr = rd_resp_desc_a_data_offset_addr_f;
   assign int_rd_resp_desc_a_data_size_size = rd_resp_desc_a_data_size_size_f;
   assign int_rd_resp_desc_a_data_host_addr_0_addr = rd_resp_desc_a_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_a_data_host_addr_1_addr = rd_resp_desc_a_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_a_data_host_addr_2_addr = rd_resp_desc_a_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_a_data_host_addr_3_addr = rd_resp_desc_a_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_a_resp_resp = rd_resp_desc_a_resp_resp_f;
   assign int_rd_resp_desc_a_xid_0_xid = rd_resp_desc_a_xid_0_xid_f;
   assign int_rd_resp_desc_a_xid_1_xid = rd_resp_desc_a_xid_1_xid_f;
   assign int_rd_resp_desc_a_xid_2_xid = rd_resp_desc_a_xid_2_xid_f;
   assign int_rd_resp_desc_a_xid_3_xid = rd_resp_desc_a_xid_3_xid_f;
   assign int_rd_resp_desc_a_xuser_0_xuser = rd_resp_desc_a_xuser_0_xuser_f;
   assign int_rd_resp_desc_a_xuser_1_xuser = rd_resp_desc_a_xuser_1_xuser_f;
   assign int_rd_resp_desc_a_xuser_2_xuser = rd_resp_desc_a_xuser_2_xuser_f;
   assign int_rd_resp_desc_a_xuser_3_xuser = rd_resp_desc_a_xuser_3_xuser_f;
   assign int_rd_resp_desc_a_xuser_4_xuser = rd_resp_desc_a_xuser_4_xuser_f;
   assign int_rd_resp_desc_a_xuser_5_xuser = rd_resp_desc_a_xuser_5_xuser_f;
   assign int_rd_resp_desc_a_xuser_6_xuser = rd_resp_desc_a_xuser_6_xuser_f;
   assign int_rd_resp_desc_a_xuser_7_xuser = rd_resp_desc_a_xuser_7_xuser_f;
   assign int_rd_resp_desc_a_xuser_8_xuser = rd_resp_desc_a_xuser_8_xuser_f;
   assign int_rd_resp_desc_a_xuser_9_xuser = rd_resp_desc_a_xuser_9_xuser_f;
   assign int_rd_resp_desc_a_xuser_10_xuser = rd_resp_desc_a_xuser_10_xuser_f;
   assign int_rd_resp_desc_a_xuser_11_xuser = rd_resp_desc_a_xuser_11_xuser_f;
   assign int_rd_resp_desc_a_xuser_12_xuser = rd_resp_desc_a_xuser_12_xuser_f;
   assign int_rd_resp_desc_a_xuser_13_xuser = rd_resp_desc_a_xuser_13_xuser_f;
   assign int_rd_resp_desc_a_xuser_14_xuser = rd_resp_desc_a_xuser_14_xuser_f;
   assign int_rd_resp_desc_a_xuser_15_xuser = rd_resp_desc_a_xuser_15_xuser_f;
   assign int_wr_req_desc_a_data_host_addr_0_addr = wr_req_desc_a_data_host_addr_0_addr_f;
   assign int_wr_req_desc_a_data_host_addr_1_addr = wr_req_desc_a_data_host_addr_1_addr_f;
   assign int_wr_req_desc_a_data_host_addr_2_addr = wr_req_desc_a_data_host_addr_2_addr_f;
   assign int_wr_req_desc_a_data_host_addr_3_addr = wr_req_desc_a_data_host_addr_3_addr_f;
   assign int_wr_req_desc_a_wstrb_host_addr_0_addr = wr_req_desc_a_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_a_wstrb_host_addr_1_addr = wr_req_desc_a_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_a_wstrb_host_addr_2_addr = wr_req_desc_a_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_a_wstrb_host_addr_3_addr = wr_req_desc_a_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_a_resp_resp = wr_resp_desc_a_resp_resp_f;
   assign int_wr_resp_desc_a_xid_0_xid = wr_resp_desc_a_xid_0_xid_f;
   assign int_wr_resp_desc_a_xid_1_xid = wr_resp_desc_a_xid_1_xid_f;
   assign int_wr_resp_desc_a_xid_2_xid = wr_resp_desc_a_xid_2_xid_f;
   assign int_wr_resp_desc_a_xid_3_xid = wr_resp_desc_a_xid_3_xid_f;
   assign int_wr_resp_desc_a_xuser_0_xuser = wr_resp_desc_a_xuser_0_xuser_f;
   assign int_wr_resp_desc_a_xuser_1_xuser = wr_resp_desc_a_xuser_1_xuser_f;
   assign int_wr_resp_desc_a_xuser_2_xuser = wr_resp_desc_a_xuser_2_xuser_f;
   assign int_wr_resp_desc_a_xuser_3_xuser = wr_resp_desc_a_xuser_3_xuser_f;
   assign int_wr_resp_desc_a_xuser_4_xuser = wr_resp_desc_a_xuser_4_xuser_f;
   assign int_wr_resp_desc_a_xuser_5_xuser = wr_resp_desc_a_xuser_5_xuser_f;
   assign int_wr_resp_desc_a_xuser_6_xuser = wr_resp_desc_a_xuser_6_xuser_f;
   assign int_wr_resp_desc_a_xuser_7_xuser = wr_resp_desc_a_xuser_7_xuser_f;
   assign int_wr_resp_desc_a_xuser_8_xuser = wr_resp_desc_a_xuser_8_xuser_f;
   assign int_wr_resp_desc_a_xuser_9_xuser = wr_resp_desc_a_xuser_9_xuser_f;
   assign int_wr_resp_desc_a_xuser_10_xuser = wr_resp_desc_a_xuser_10_xuser_f;
   assign int_wr_resp_desc_a_xuser_11_xuser = wr_resp_desc_a_xuser_11_xuser_f;
   assign int_wr_resp_desc_a_xuser_12_xuser = wr_resp_desc_a_xuser_12_xuser_f;
   assign int_wr_resp_desc_a_xuser_13_xuser = wr_resp_desc_a_xuser_13_xuser_f;
   assign int_wr_resp_desc_a_xuser_14_xuser = wr_resp_desc_a_xuser_14_xuser_f;
   assign int_wr_resp_desc_a_xuser_15_xuser = wr_resp_desc_a_xuser_15_xuser_f;
   assign int_sn_req_desc_a_attr_acsnoop = sn_req_desc_a_attr_acsnoop_f;
   assign int_sn_req_desc_a_attr_acprot = sn_req_desc_a_attr_acprot_f;
   assign int_sn_req_desc_a_acaddr_0_addr = sn_req_desc_a_acaddr_0_addr_f;
   assign int_sn_req_desc_a_acaddr_1_addr = sn_req_desc_a_acaddr_1_addr_f;
   assign int_sn_req_desc_a_acaddr_2_addr = sn_req_desc_a_acaddr_2_addr_f;
   assign int_sn_req_desc_a_acaddr_3_addr = sn_req_desc_a_acaddr_3_addr_f;
   assign int_rd_resp_desc_b_data_offset_addr = rd_resp_desc_b_data_offset_addr_f;
   assign int_rd_resp_desc_b_data_size_size = rd_resp_desc_b_data_size_size_f;
   assign int_rd_resp_desc_b_data_host_addr_0_addr = rd_resp_desc_b_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_b_data_host_addr_1_addr = rd_resp_desc_b_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_b_data_host_addr_2_addr = rd_resp_desc_b_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_b_data_host_addr_3_addr = rd_resp_desc_b_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_b_resp_resp = rd_resp_desc_b_resp_resp_f;
   assign int_rd_resp_desc_b_xid_0_xid = rd_resp_desc_b_xid_0_xid_f;
   assign int_rd_resp_desc_b_xid_1_xid = rd_resp_desc_b_xid_1_xid_f;
   assign int_rd_resp_desc_b_xid_2_xid = rd_resp_desc_b_xid_2_xid_f;
   assign int_rd_resp_desc_b_xid_3_xid = rd_resp_desc_b_xid_3_xid_f;
   assign int_rd_resp_desc_b_xuser_0_xuser = rd_resp_desc_b_xuser_0_xuser_f;
   assign int_rd_resp_desc_b_xuser_1_xuser = rd_resp_desc_b_xuser_1_xuser_f;
   assign int_rd_resp_desc_b_xuser_2_xuser = rd_resp_desc_b_xuser_2_xuser_f;
   assign int_rd_resp_desc_b_xuser_3_xuser = rd_resp_desc_b_xuser_3_xuser_f;
   assign int_rd_resp_desc_b_xuser_4_xuser = rd_resp_desc_b_xuser_4_xuser_f;
   assign int_rd_resp_desc_b_xuser_5_xuser = rd_resp_desc_b_xuser_5_xuser_f;
   assign int_rd_resp_desc_b_xuser_6_xuser = rd_resp_desc_b_xuser_6_xuser_f;
   assign int_rd_resp_desc_b_xuser_7_xuser = rd_resp_desc_b_xuser_7_xuser_f;
   assign int_rd_resp_desc_b_xuser_8_xuser = rd_resp_desc_b_xuser_8_xuser_f;
   assign int_rd_resp_desc_b_xuser_9_xuser = rd_resp_desc_b_xuser_9_xuser_f;
   assign int_rd_resp_desc_b_xuser_10_xuser = rd_resp_desc_b_xuser_10_xuser_f;
   assign int_rd_resp_desc_b_xuser_11_xuser = rd_resp_desc_b_xuser_11_xuser_f;
   assign int_rd_resp_desc_b_xuser_12_xuser = rd_resp_desc_b_xuser_12_xuser_f;
   assign int_rd_resp_desc_b_xuser_13_xuser = rd_resp_desc_b_xuser_13_xuser_f;
   assign int_rd_resp_desc_b_xuser_14_xuser = rd_resp_desc_b_xuser_14_xuser_f;
   assign int_rd_resp_desc_b_xuser_15_xuser = rd_resp_desc_b_xuser_15_xuser_f;
   assign int_wr_req_desc_b_data_host_addr_0_addr = wr_req_desc_b_data_host_addr_0_addr_f;
   assign int_wr_req_desc_b_data_host_addr_1_addr = wr_req_desc_b_data_host_addr_1_addr_f;
   assign int_wr_req_desc_b_data_host_addr_2_addr = wr_req_desc_b_data_host_addr_2_addr_f;
   assign int_wr_req_desc_b_data_host_addr_3_addr = wr_req_desc_b_data_host_addr_3_addr_f;
   assign int_wr_req_desc_b_wstrb_host_addr_0_addr = wr_req_desc_b_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_b_wstrb_host_addr_1_addr = wr_req_desc_b_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_b_wstrb_host_addr_2_addr = wr_req_desc_b_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_b_wstrb_host_addr_3_addr = wr_req_desc_b_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_b_resp_resp = wr_resp_desc_b_resp_resp_f;
   assign int_wr_resp_desc_b_xid_0_xid = wr_resp_desc_b_xid_0_xid_f;
   assign int_wr_resp_desc_b_xid_1_xid = wr_resp_desc_b_xid_1_xid_f;
   assign int_wr_resp_desc_b_xid_2_xid = wr_resp_desc_b_xid_2_xid_f;
   assign int_wr_resp_desc_b_xid_3_xid = wr_resp_desc_b_xid_3_xid_f;
   assign int_wr_resp_desc_b_xuser_0_xuser = wr_resp_desc_b_xuser_0_xuser_f;
   assign int_wr_resp_desc_b_xuser_1_xuser = wr_resp_desc_b_xuser_1_xuser_f;
   assign int_wr_resp_desc_b_xuser_2_xuser = wr_resp_desc_b_xuser_2_xuser_f;
   assign int_wr_resp_desc_b_xuser_3_xuser = wr_resp_desc_b_xuser_3_xuser_f;
   assign int_wr_resp_desc_b_xuser_4_xuser = wr_resp_desc_b_xuser_4_xuser_f;
   assign int_wr_resp_desc_b_xuser_5_xuser = wr_resp_desc_b_xuser_5_xuser_f;
   assign int_wr_resp_desc_b_xuser_6_xuser = wr_resp_desc_b_xuser_6_xuser_f;
   assign int_wr_resp_desc_b_xuser_7_xuser = wr_resp_desc_b_xuser_7_xuser_f;
   assign int_wr_resp_desc_b_xuser_8_xuser = wr_resp_desc_b_xuser_8_xuser_f;
   assign int_wr_resp_desc_b_xuser_9_xuser = wr_resp_desc_b_xuser_9_xuser_f;
   assign int_wr_resp_desc_b_xuser_10_xuser = wr_resp_desc_b_xuser_10_xuser_f;
   assign int_wr_resp_desc_b_xuser_11_xuser = wr_resp_desc_b_xuser_11_xuser_f;
   assign int_wr_resp_desc_b_xuser_12_xuser = wr_resp_desc_b_xuser_12_xuser_f;
   assign int_wr_resp_desc_b_xuser_13_xuser = wr_resp_desc_b_xuser_13_xuser_f;
   assign int_wr_resp_desc_b_xuser_14_xuser = wr_resp_desc_b_xuser_14_xuser_f;
   assign int_wr_resp_desc_b_xuser_15_xuser = wr_resp_desc_b_xuser_15_xuser_f;
   assign int_sn_req_desc_b_attr_acsnoop = sn_req_desc_b_attr_acsnoop_f;
   assign int_sn_req_desc_b_attr_acprot = sn_req_desc_b_attr_acprot_f;
   assign int_sn_req_desc_b_acaddr_0_addr = sn_req_desc_b_acaddr_0_addr_f;
   assign int_sn_req_desc_b_acaddr_1_addr = sn_req_desc_b_acaddr_1_addr_f;
   assign int_sn_req_desc_b_acaddr_2_addr = sn_req_desc_b_acaddr_2_addr_f;
   assign int_sn_req_desc_b_acaddr_3_addr = sn_req_desc_b_acaddr_3_addr_f;
   assign int_rd_resp_desc_c_data_offset_addr = rd_resp_desc_c_data_offset_addr_f;
   assign int_rd_resp_desc_c_data_size_size = rd_resp_desc_c_data_size_size_f;
   assign int_rd_resp_desc_c_data_host_addr_0_addr = rd_resp_desc_c_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_c_data_host_addr_1_addr = rd_resp_desc_c_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_c_data_host_addr_2_addr = rd_resp_desc_c_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_c_data_host_addr_3_addr = rd_resp_desc_c_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_c_resp_resp = rd_resp_desc_c_resp_resp_f;
   assign int_rd_resp_desc_c_xid_0_xid = rd_resp_desc_c_xid_0_xid_f;
   assign int_rd_resp_desc_c_xid_1_xid = rd_resp_desc_c_xid_1_xid_f;
   assign int_rd_resp_desc_c_xid_2_xid = rd_resp_desc_c_xid_2_xid_f;
   assign int_rd_resp_desc_c_xid_3_xid = rd_resp_desc_c_xid_3_xid_f;
   assign int_rd_resp_desc_c_xuser_0_xuser = rd_resp_desc_c_xuser_0_xuser_f;
   assign int_rd_resp_desc_c_xuser_1_xuser = rd_resp_desc_c_xuser_1_xuser_f;
   assign int_rd_resp_desc_c_xuser_2_xuser = rd_resp_desc_c_xuser_2_xuser_f;
   assign int_rd_resp_desc_c_xuser_3_xuser = rd_resp_desc_c_xuser_3_xuser_f;
   assign int_rd_resp_desc_c_xuser_4_xuser = rd_resp_desc_c_xuser_4_xuser_f;
   assign int_rd_resp_desc_c_xuser_5_xuser = rd_resp_desc_c_xuser_5_xuser_f;
   assign int_rd_resp_desc_c_xuser_6_xuser = rd_resp_desc_c_xuser_6_xuser_f;
   assign int_rd_resp_desc_c_xuser_7_xuser = rd_resp_desc_c_xuser_7_xuser_f;
   assign int_rd_resp_desc_c_xuser_8_xuser = rd_resp_desc_c_xuser_8_xuser_f;
   assign int_rd_resp_desc_c_xuser_9_xuser = rd_resp_desc_c_xuser_9_xuser_f;
   assign int_rd_resp_desc_c_xuser_10_xuser = rd_resp_desc_c_xuser_10_xuser_f;
   assign int_rd_resp_desc_c_xuser_11_xuser = rd_resp_desc_c_xuser_11_xuser_f;
   assign int_rd_resp_desc_c_xuser_12_xuser = rd_resp_desc_c_xuser_12_xuser_f;
   assign int_rd_resp_desc_c_xuser_13_xuser = rd_resp_desc_c_xuser_13_xuser_f;
   assign int_rd_resp_desc_c_xuser_14_xuser = rd_resp_desc_c_xuser_14_xuser_f;
   assign int_rd_resp_desc_c_xuser_15_xuser = rd_resp_desc_c_xuser_15_xuser_f;
   assign int_wr_req_desc_c_data_host_addr_0_addr = wr_req_desc_c_data_host_addr_0_addr_f;
   assign int_wr_req_desc_c_data_host_addr_1_addr = wr_req_desc_c_data_host_addr_1_addr_f;
   assign int_wr_req_desc_c_data_host_addr_2_addr = wr_req_desc_c_data_host_addr_2_addr_f;
   assign int_wr_req_desc_c_data_host_addr_3_addr = wr_req_desc_c_data_host_addr_3_addr_f;
   assign int_wr_req_desc_c_wstrb_host_addr_0_addr = wr_req_desc_c_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_c_wstrb_host_addr_1_addr = wr_req_desc_c_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_c_wstrb_host_addr_2_addr = wr_req_desc_c_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_c_wstrb_host_addr_3_addr = wr_req_desc_c_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_c_resp_resp = wr_resp_desc_c_resp_resp_f;
   assign int_wr_resp_desc_c_xid_0_xid = wr_resp_desc_c_xid_0_xid_f;
   assign int_wr_resp_desc_c_xid_1_xid = wr_resp_desc_c_xid_1_xid_f;
   assign int_wr_resp_desc_c_xid_2_xid = wr_resp_desc_c_xid_2_xid_f;
   assign int_wr_resp_desc_c_xid_3_xid = wr_resp_desc_c_xid_3_xid_f;
   assign int_wr_resp_desc_c_xuser_0_xuser = wr_resp_desc_c_xuser_0_xuser_f;
   assign int_wr_resp_desc_c_xuser_1_xuser = wr_resp_desc_c_xuser_1_xuser_f;
   assign int_wr_resp_desc_c_xuser_2_xuser = wr_resp_desc_c_xuser_2_xuser_f;
   assign int_wr_resp_desc_c_xuser_3_xuser = wr_resp_desc_c_xuser_3_xuser_f;
   assign int_wr_resp_desc_c_xuser_4_xuser = wr_resp_desc_c_xuser_4_xuser_f;
   assign int_wr_resp_desc_c_xuser_5_xuser = wr_resp_desc_c_xuser_5_xuser_f;
   assign int_wr_resp_desc_c_xuser_6_xuser = wr_resp_desc_c_xuser_6_xuser_f;
   assign int_wr_resp_desc_c_xuser_7_xuser = wr_resp_desc_c_xuser_7_xuser_f;
   assign int_wr_resp_desc_c_xuser_8_xuser = wr_resp_desc_c_xuser_8_xuser_f;
   assign int_wr_resp_desc_c_xuser_9_xuser = wr_resp_desc_c_xuser_9_xuser_f;
   assign int_wr_resp_desc_c_xuser_10_xuser = wr_resp_desc_c_xuser_10_xuser_f;
   assign int_wr_resp_desc_c_xuser_11_xuser = wr_resp_desc_c_xuser_11_xuser_f;
   assign int_wr_resp_desc_c_xuser_12_xuser = wr_resp_desc_c_xuser_12_xuser_f;
   assign int_wr_resp_desc_c_xuser_13_xuser = wr_resp_desc_c_xuser_13_xuser_f;
   assign int_wr_resp_desc_c_xuser_14_xuser = wr_resp_desc_c_xuser_14_xuser_f;
   assign int_wr_resp_desc_c_xuser_15_xuser = wr_resp_desc_c_xuser_15_xuser_f;
   assign int_sn_req_desc_c_attr_acsnoop = sn_req_desc_c_attr_acsnoop_f;
   assign int_sn_req_desc_c_attr_acprot = sn_req_desc_c_attr_acprot_f;
   assign int_sn_req_desc_c_acaddr_0_addr = sn_req_desc_c_acaddr_0_addr_f;
   assign int_sn_req_desc_c_acaddr_1_addr = sn_req_desc_c_acaddr_1_addr_f;
   assign int_sn_req_desc_c_acaddr_2_addr = sn_req_desc_c_acaddr_2_addr_f;
   assign int_sn_req_desc_c_acaddr_3_addr = sn_req_desc_c_acaddr_3_addr_f;
   assign int_rd_resp_desc_d_data_offset_addr = rd_resp_desc_d_data_offset_addr_f;
   assign int_rd_resp_desc_d_data_size_size = rd_resp_desc_d_data_size_size_f;
   assign int_rd_resp_desc_d_data_host_addr_0_addr = rd_resp_desc_d_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_d_data_host_addr_1_addr = rd_resp_desc_d_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_d_data_host_addr_2_addr = rd_resp_desc_d_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_d_data_host_addr_3_addr = rd_resp_desc_d_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_d_resp_resp = rd_resp_desc_d_resp_resp_f;
   assign int_rd_resp_desc_d_xid_0_xid = rd_resp_desc_d_xid_0_xid_f;
   assign int_rd_resp_desc_d_xid_1_xid = rd_resp_desc_d_xid_1_xid_f;
   assign int_rd_resp_desc_d_xid_2_xid = rd_resp_desc_d_xid_2_xid_f;
   assign int_rd_resp_desc_d_xid_3_xid = rd_resp_desc_d_xid_3_xid_f;
   assign int_rd_resp_desc_d_xuser_0_xuser = rd_resp_desc_d_xuser_0_xuser_f;
   assign int_rd_resp_desc_d_xuser_1_xuser = rd_resp_desc_d_xuser_1_xuser_f;
   assign int_rd_resp_desc_d_xuser_2_xuser = rd_resp_desc_d_xuser_2_xuser_f;
   assign int_rd_resp_desc_d_xuser_3_xuser = rd_resp_desc_d_xuser_3_xuser_f;
   assign int_rd_resp_desc_d_xuser_4_xuser = rd_resp_desc_d_xuser_4_xuser_f;
   assign int_rd_resp_desc_d_xuser_5_xuser = rd_resp_desc_d_xuser_5_xuser_f;
   assign int_rd_resp_desc_d_xuser_6_xuser = rd_resp_desc_d_xuser_6_xuser_f;
   assign int_rd_resp_desc_d_xuser_7_xuser = rd_resp_desc_d_xuser_7_xuser_f;
   assign int_rd_resp_desc_d_xuser_8_xuser = rd_resp_desc_d_xuser_8_xuser_f;
   assign int_rd_resp_desc_d_xuser_9_xuser = rd_resp_desc_d_xuser_9_xuser_f;
   assign int_rd_resp_desc_d_xuser_10_xuser = rd_resp_desc_d_xuser_10_xuser_f;
   assign int_rd_resp_desc_d_xuser_11_xuser = rd_resp_desc_d_xuser_11_xuser_f;
   assign int_rd_resp_desc_d_xuser_12_xuser = rd_resp_desc_d_xuser_12_xuser_f;
   assign int_rd_resp_desc_d_xuser_13_xuser = rd_resp_desc_d_xuser_13_xuser_f;
   assign int_rd_resp_desc_d_xuser_14_xuser = rd_resp_desc_d_xuser_14_xuser_f;
   assign int_rd_resp_desc_d_xuser_15_xuser = rd_resp_desc_d_xuser_15_xuser_f;
   assign int_wr_req_desc_d_data_host_addr_0_addr = wr_req_desc_d_data_host_addr_0_addr_f;
   assign int_wr_req_desc_d_data_host_addr_1_addr = wr_req_desc_d_data_host_addr_1_addr_f;
   assign int_wr_req_desc_d_data_host_addr_2_addr = wr_req_desc_d_data_host_addr_2_addr_f;
   assign int_wr_req_desc_d_data_host_addr_3_addr = wr_req_desc_d_data_host_addr_3_addr_f;
   assign int_wr_req_desc_d_wstrb_host_addr_0_addr = wr_req_desc_d_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_d_wstrb_host_addr_1_addr = wr_req_desc_d_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_d_wstrb_host_addr_2_addr = wr_req_desc_d_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_d_wstrb_host_addr_3_addr = wr_req_desc_d_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_d_resp_resp = wr_resp_desc_d_resp_resp_f;
   assign int_wr_resp_desc_d_xid_0_xid = wr_resp_desc_d_xid_0_xid_f;
   assign int_wr_resp_desc_d_xid_1_xid = wr_resp_desc_d_xid_1_xid_f;
   assign int_wr_resp_desc_d_xid_2_xid = wr_resp_desc_d_xid_2_xid_f;
   assign int_wr_resp_desc_d_xid_3_xid = wr_resp_desc_d_xid_3_xid_f;
   assign int_wr_resp_desc_d_xuser_0_xuser = wr_resp_desc_d_xuser_0_xuser_f;
   assign int_wr_resp_desc_d_xuser_1_xuser = wr_resp_desc_d_xuser_1_xuser_f;
   assign int_wr_resp_desc_d_xuser_2_xuser = wr_resp_desc_d_xuser_2_xuser_f;
   assign int_wr_resp_desc_d_xuser_3_xuser = wr_resp_desc_d_xuser_3_xuser_f;
   assign int_wr_resp_desc_d_xuser_4_xuser = wr_resp_desc_d_xuser_4_xuser_f;
   assign int_wr_resp_desc_d_xuser_5_xuser = wr_resp_desc_d_xuser_5_xuser_f;
   assign int_wr_resp_desc_d_xuser_6_xuser = wr_resp_desc_d_xuser_6_xuser_f;
   assign int_wr_resp_desc_d_xuser_7_xuser = wr_resp_desc_d_xuser_7_xuser_f;
   assign int_wr_resp_desc_d_xuser_8_xuser = wr_resp_desc_d_xuser_8_xuser_f;
   assign int_wr_resp_desc_d_xuser_9_xuser = wr_resp_desc_d_xuser_9_xuser_f;
   assign int_wr_resp_desc_d_xuser_10_xuser = wr_resp_desc_d_xuser_10_xuser_f;
   assign int_wr_resp_desc_d_xuser_11_xuser = wr_resp_desc_d_xuser_11_xuser_f;
   assign int_wr_resp_desc_d_xuser_12_xuser = wr_resp_desc_d_xuser_12_xuser_f;
   assign int_wr_resp_desc_d_xuser_13_xuser = wr_resp_desc_d_xuser_13_xuser_f;
   assign int_wr_resp_desc_d_xuser_14_xuser = wr_resp_desc_d_xuser_14_xuser_f;
   assign int_wr_resp_desc_d_xuser_15_xuser = wr_resp_desc_d_xuser_15_xuser_f;
   assign int_sn_req_desc_d_attr_acsnoop = sn_req_desc_d_attr_acsnoop_f;
   assign int_sn_req_desc_d_attr_acprot = sn_req_desc_d_attr_acprot_f;
   assign int_sn_req_desc_d_acaddr_0_addr = sn_req_desc_d_acaddr_0_addr_f;
   assign int_sn_req_desc_d_acaddr_1_addr = sn_req_desc_d_acaddr_1_addr_f;
   assign int_sn_req_desc_d_acaddr_2_addr = sn_req_desc_d_acaddr_2_addr_f;
   assign int_sn_req_desc_d_acaddr_3_addr = sn_req_desc_d_acaddr_3_addr_f;
   assign int_rd_resp_desc_e_data_offset_addr = rd_resp_desc_e_data_offset_addr_f;
   assign int_rd_resp_desc_e_data_size_size = rd_resp_desc_e_data_size_size_f;
   assign int_rd_resp_desc_e_data_host_addr_0_addr = rd_resp_desc_e_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_e_data_host_addr_1_addr = rd_resp_desc_e_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_e_data_host_addr_2_addr = rd_resp_desc_e_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_e_data_host_addr_3_addr = rd_resp_desc_e_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_e_resp_resp = rd_resp_desc_e_resp_resp_f;
   assign int_rd_resp_desc_e_xid_0_xid = rd_resp_desc_e_xid_0_xid_f;
   assign int_rd_resp_desc_e_xid_1_xid = rd_resp_desc_e_xid_1_xid_f;
   assign int_rd_resp_desc_e_xid_2_xid = rd_resp_desc_e_xid_2_xid_f;
   assign int_rd_resp_desc_e_xid_3_xid = rd_resp_desc_e_xid_3_xid_f;
   assign int_rd_resp_desc_e_xuser_0_xuser = rd_resp_desc_e_xuser_0_xuser_f;
   assign int_rd_resp_desc_e_xuser_1_xuser = rd_resp_desc_e_xuser_1_xuser_f;
   assign int_rd_resp_desc_e_xuser_2_xuser = rd_resp_desc_e_xuser_2_xuser_f;
   assign int_rd_resp_desc_e_xuser_3_xuser = rd_resp_desc_e_xuser_3_xuser_f;
   assign int_rd_resp_desc_e_xuser_4_xuser = rd_resp_desc_e_xuser_4_xuser_f;
   assign int_rd_resp_desc_e_xuser_5_xuser = rd_resp_desc_e_xuser_5_xuser_f;
   assign int_rd_resp_desc_e_xuser_6_xuser = rd_resp_desc_e_xuser_6_xuser_f;
   assign int_rd_resp_desc_e_xuser_7_xuser = rd_resp_desc_e_xuser_7_xuser_f;
   assign int_rd_resp_desc_e_xuser_8_xuser = rd_resp_desc_e_xuser_8_xuser_f;
   assign int_rd_resp_desc_e_xuser_9_xuser = rd_resp_desc_e_xuser_9_xuser_f;
   assign int_rd_resp_desc_e_xuser_10_xuser = rd_resp_desc_e_xuser_10_xuser_f;
   assign int_rd_resp_desc_e_xuser_11_xuser = rd_resp_desc_e_xuser_11_xuser_f;
   assign int_rd_resp_desc_e_xuser_12_xuser = rd_resp_desc_e_xuser_12_xuser_f;
   assign int_rd_resp_desc_e_xuser_13_xuser = rd_resp_desc_e_xuser_13_xuser_f;
   assign int_rd_resp_desc_e_xuser_14_xuser = rd_resp_desc_e_xuser_14_xuser_f;
   assign int_rd_resp_desc_e_xuser_15_xuser = rd_resp_desc_e_xuser_15_xuser_f;
   assign int_wr_req_desc_e_data_host_addr_0_addr = wr_req_desc_e_data_host_addr_0_addr_f;
   assign int_wr_req_desc_e_data_host_addr_1_addr = wr_req_desc_e_data_host_addr_1_addr_f;
   assign int_wr_req_desc_e_data_host_addr_2_addr = wr_req_desc_e_data_host_addr_2_addr_f;
   assign int_wr_req_desc_e_data_host_addr_3_addr = wr_req_desc_e_data_host_addr_3_addr_f;
   assign int_wr_req_desc_e_wstrb_host_addr_0_addr = wr_req_desc_e_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_e_wstrb_host_addr_1_addr = wr_req_desc_e_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_e_wstrb_host_addr_2_addr = wr_req_desc_e_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_e_wstrb_host_addr_3_addr = wr_req_desc_e_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_e_resp_resp = wr_resp_desc_e_resp_resp_f;
   assign int_wr_resp_desc_e_xid_0_xid = wr_resp_desc_e_xid_0_xid_f;
   assign int_wr_resp_desc_e_xid_1_xid = wr_resp_desc_e_xid_1_xid_f;
   assign int_wr_resp_desc_e_xid_2_xid = wr_resp_desc_e_xid_2_xid_f;
   assign int_wr_resp_desc_e_xid_3_xid = wr_resp_desc_e_xid_3_xid_f;
   assign int_wr_resp_desc_e_xuser_0_xuser = wr_resp_desc_e_xuser_0_xuser_f;
   assign int_wr_resp_desc_e_xuser_1_xuser = wr_resp_desc_e_xuser_1_xuser_f;
   assign int_wr_resp_desc_e_xuser_2_xuser = wr_resp_desc_e_xuser_2_xuser_f;
   assign int_wr_resp_desc_e_xuser_3_xuser = wr_resp_desc_e_xuser_3_xuser_f;
   assign int_wr_resp_desc_e_xuser_4_xuser = wr_resp_desc_e_xuser_4_xuser_f;
   assign int_wr_resp_desc_e_xuser_5_xuser = wr_resp_desc_e_xuser_5_xuser_f;
   assign int_wr_resp_desc_e_xuser_6_xuser = wr_resp_desc_e_xuser_6_xuser_f;
   assign int_wr_resp_desc_e_xuser_7_xuser = wr_resp_desc_e_xuser_7_xuser_f;
   assign int_wr_resp_desc_e_xuser_8_xuser = wr_resp_desc_e_xuser_8_xuser_f;
   assign int_wr_resp_desc_e_xuser_9_xuser = wr_resp_desc_e_xuser_9_xuser_f;
   assign int_wr_resp_desc_e_xuser_10_xuser = wr_resp_desc_e_xuser_10_xuser_f;
   assign int_wr_resp_desc_e_xuser_11_xuser = wr_resp_desc_e_xuser_11_xuser_f;
   assign int_wr_resp_desc_e_xuser_12_xuser = wr_resp_desc_e_xuser_12_xuser_f;
   assign int_wr_resp_desc_e_xuser_13_xuser = wr_resp_desc_e_xuser_13_xuser_f;
   assign int_wr_resp_desc_e_xuser_14_xuser = wr_resp_desc_e_xuser_14_xuser_f;
   assign int_wr_resp_desc_e_xuser_15_xuser = wr_resp_desc_e_xuser_15_xuser_f;
   assign int_sn_req_desc_e_attr_acsnoop = sn_req_desc_e_attr_acsnoop_f;
   assign int_sn_req_desc_e_attr_acprot = sn_req_desc_e_attr_acprot_f;
   assign int_sn_req_desc_e_acaddr_0_addr = sn_req_desc_e_acaddr_0_addr_f;
   assign int_sn_req_desc_e_acaddr_1_addr = sn_req_desc_e_acaddr_1_addr_f;
   assign int_sn_req_desc_e_acaddr_2_addr = sn_req_desc_e_acaddr_2_addr_f;
   assign int_sn_req_desc_e_acaddr_3_addr = sn_req_desc_e_acaddr_3_addr_f;
   assign int_rd_resp_desc_f_data_offset_addr = rd_resp_desc_f_data_offset_addr_f;
   assign int_rd_resp_desc_f_data_size_size = rd_resp_desc_f_data_size_size_f;
   assign int_rd_resp_desc_f_data_host_addr_0_addr = rd_resp_desc_f_data_host_addr_0_addr_f;
   assign int_rd_resp_desc_f_data_host_addr_1_addr = rd_resp_desc_f_data_host_addr_1_addr_f;
   assign int_rd_resp_desc_f_data_host_addr_2_addr = rd_resp_desc_f_data_host_addr_2_addr_f;
   assign int_rd_resp_desc_f_data_host_addr_3_addr = rd_resp_desc_f_data_host_addr_3_addr_f;
   assign int_rd_resp_desc_f_resp_resp = rd_resp_desc_f_resp_resp_f;
   assign int_rd_resp_desc_f_xid_0_xid = rd_resp_desc_f_xid_0_xid_f;
   assign int_rd_resp_desc_f_xid_1_xid = rd_resp_desc_f_xid_1_xid_f;
   assign int_rd_resp_desc_f_xid_2_xid = rd_resp_desc_f_xid_2_xid_f;
   assign int_rd_resp_desc_f_xid_3_xid = rd_resp_desc_f_xid_3_xid_f;
   assign int_rd_resp_desc_f_xuser_0_xuser = rd_resp_desc_f_xuser_0_xuser_f;
   assign int_rd_resp_desc_f_xuser_1_xuser = rd_resp_desc_f_xuser_1_xuser_f;
   assign int_rd_resp_desc_f_xuser_2_xuser = rd_resp_desc_f_xuser_2_xuser_f;
   assign int_rd_resp_desc_f_xuser_3_xuser = rd_resp_desc_f_xuser_3_xuser_f;
   assign int_rd_resp_desc_f_xuser_4_xuser = rd_resp_desc_f_xuser_4_xuser_f;
   assign int_rd_resp_desc_f_xuser_5_xuser = rd_resp_desc_f_xuser_5_xuser_f;
   assign int_rd_resp_desc_f_xuser_6_xuser = rd_resp_desc_f_xuser_6_xuser_f;
   assign int_rd_resp_desc_f_xuser_7_xuser = rd_resp_desc_f_xuser_7_xuser_f;
   assign int_rd_resp_desc_f_xuser_8_xuser = rd_resp_desc_f_xuser_8_xuser_f;
   assign int_rd_resp_desc_f_xuser_9_xuser = rd_resp_desc_f_xuser_9_xuser_f;
   assign int_rd_resp_desc_f_xuser_10_xuser = rd_resp_desc_f_xuser_10_xuser_f;
   assign int_rd_resp_desc_f_xuser_11_xuser = rd_resp_desc_f_xuser_11_xuser_f;
   assign int_rd_resp_desc_f_xuser_12_xuser = rd_resp_desc_f_xuser_12_xuser_f;
   assign int_rd_resp_desc_f_xuser_13_xuser = rd_resp_desc_f_xuser_13_xuser_f;
   assign int_rd_resp_desc_f_xuser_14_xuser = rd_resp_desc_f_xuser_14_xuser_f;
   assign int_rd_resp_desc_f_xuser_15_xuser = rd_resp_desc_f_xuser_15_xuser_f;
   assign int_wr_req_desc_f_data_host_addr_0_addr = wr_req_desc_f_data_host_addr_0_addr_f;
   assign int_wr_req_desc_f_data_host_addr_1_addr = wr_req_desc_f_data_host_addr_1_addr_f;
   assign int_wr_req_desc_f_data_host_addr_2_addr = wr_req_desc_f_data_host_addr_2_addr_f;
   assign int_wr_req_desc_f_data_host_addr_3_addr = wr_req_desc_f_data_host_addr_3_addr_f;
   assign int_wr_req_desc_f_wstrb_host_addr_0_addr = wr_req_desc_f_wstrb_host_addr_0_addr_f;
   assign int_wr_req_desc_f_wstrb_host_addr_1_addr = wr_req_desc_f_wstrb_host_addr_1_addr_f;
   assign int_wr_req_desc_f_wstrb_host_addr_2_addr = wr_req_desc_f_wstrb_host_addr_2_addr_f;
   assign int_wr_req_desc_f_wstrb_host_addr_3_addr = wr_req_desc_f_wstrb_host_addr_3_addr_f;
   assign int_wr_resp_desc_f_resp_resp = wr_resp_desc_f_resp_resp_f;
   assign int_wr_resp_desc_f_xid_0_xid = wr_resp_desc_f_xid_0_xid_f;
   assign int_wr_resp_desc_f_xid_1_xid = wr_resp_desc_f_xid_1_xid_f;
   assign int_wr_resp_desc_f_xid_2_xid = wr_resp_desc_f_xid_2_xid_f;
   assign int_wr_resp_desc_f_xid_3_xid = wr_resp_desc_f_xid_3_xid_f;
   assign int_wr_resp_desc_f_xuser_0_xuser = wr_resp_desc_f_xuser_0_xuser_f;
   assign int_wr_resp_desc_f_xuser_1_xuser = wr_resp_desc_f_xuser_1_xuser_f;
   assign int_wr_resp_desc_f_xuser_2_xuser = wr_resp_desc_f_xuser_2_xuser_f;
   assign int_wr_resp_desc_f_xuser_3_xuser = wr_resp_desc_f_xuser_3_xuser_f;
   assign int_wr_resp_desc_f_xuser_4_xuser = wr_resp_desc_f_xuser_4_xuser_f;
   assign int_wr_resp_desc_f_xuser_5_xuser = wr_resp_desc_f_xuser_5_xuser_f;
   assign int_wr_resp_desc_f_xuser_6_xuser = wr_resp_desc_f_xuser_6_xuser_f;
   assign int_wr_resp_desc_f_xuser_7_xuser = wr_resp_desc_f_xuser_7_xuser_f;
   assign int_wr_resp_desc_f_xuser_8_xuser = wr_resp_desc_f_xuser_8_xuser_f;
   assign int_wr_resp_desc_f_xuser_9_xuser = wr_resp_desc_f_xuser_9_xuser_f;
   assign int_wr_resp_desc_f_xuser_10_xuser = wr_resp_desc_f_xuser_10_xuser_f;
   assign int_wr_resp_desc_f_xuser_11_xuser = wr_resp_desc_f_xuser_11_xuser_f;
   assign int_wr_resp_desc_f_xuser_12_xuser = wr_resp_desc_f_xuser_12_xuser_f;
   assign int_wr_resp_desc_f_xuser_13_xuser = wr_resp_desc_f_xuser_13_xuser_f;
   assign int_wr_resp_desc_f_xuser_14_xuser = wr_resp_desc_f_xuser_14_xuser_f;
   assign int_wr_resp_desc_f_xuser_15_xuser = wr_resp_desc_f_xuser_15_xuser_f;
   assign int_sn_req_desc_f_attr_acsnoop = sn_req_desc_f_attr_acsnoop_f;
   assign int_sn_req_desc_f_attr_acprot = sn_req_desc_f_attr_acprot_f;
   assign int_sn_req_desc_f_acaddr_0_addr = sn_req_desc_f_acaddr_0_addr_f;
   assign int_sn_req_desc_f_acaddr_1_addr = sn_req_desc_f_acaddr_1_addr_f;
   assign int_sn_req_desc_f_acaddr_2_addr = sn_req_desc_f_acaddr_2_addr_f;
   assign int_sn_req_desc_f_acaddr_3_addr = sn_req_desc_f_acaddr_3_addr_f;


   //Signals to be given as input to RB

   assign uc2rb_intr_error_status_reg[0] = int_intr_error_status_err_0;
   assign uc2rb_rd_req_fifo_pop_desc_reg[31] = int_rd_req_fifo_pop_desc_valid;
   assign uc2rb_rd_req_fifo_pop_desc_reg[3:0] = int_rd_req_fifo_pop_desc_desc_index;
   assign uc2rb_rd_req_fifo_fill_level_reg[4:0] = int_rd_req_fifo_fill_level_fill;
   assign uc2rb_rd_resp_fifo_free_level_reg[4:0] = int_rd_resp_fifo_free_level_free;
   assign uc2rb_rd_resp_intr_comp_status_reg[15:0] = int_rd_resp_intr_comp_status_comp;
   assign uc2rb_wr_req_fifo_pop_desc_reg[31] = int_wr_req_fifo_pop_desc_valid;
   assign uc2rb_wr_req_fifo_pop_desc_reg[3:0] = int_wr_req_fifo_pop_desc_desc_index;
   assign uc2rb_wr_req_fifo_fill_level_reg[4:0] = int_wr_req_fifo_fill_level_fill;
   assign uc2rb_wr_resp_fifo_free_level_reg[4:0] = int_wr_resp_fifo_free_level_free;
   assign uc2rb_wr_resp_intr_comp_status_reg[15:0] = int_wr_resp_intr_comp_status_comp;
   assign uc2rb_sn_req_fifo_free_level_reg[4:0] = int_sn_req_fifo_free_level_free;
   assign uc2rb_sn_req_intr_comp_status_reg[15:0] = int_sn_req_intr_comp_status_comp;
   assign uc2rb_sn_resp_fifo_pop_desc_reg[31] = int_sn_resp_fifo_pop_desc_valid;
   assign uc2rb_sn_resp_fifo_pop_desc_reg[3:0] = int_sn_resp_fifo_pop_desc_desc_index;
   assign uc2rb_sn_resp_fifo_fill_level_reg[4:0] = int_sn_resp_fifo_fill_level_fill;
   assign uc2rb_sn_data_fifo_pop_desc_reg[31] = int_sn_data_fifo_pop_desc_valid;
   assign uc2rb_sn_data_fifo_pop_desc_reg[3:0] = int_sn_data_fifo_pop_desc_desc_index;
   assign uc2rb_sn_data_fifo_fill_level_reg[4:0] = int_sn_data_fifo_fill_level_fill;
   assign uc2rb_rd_req_desc_0_size_reg[31:0] = int_rd_req_desc_0_size_txn_size;
   assign uc2rb_rd_req_desc_0_axsize_reg[2:0] = int_rd_req_desc_0_axsize_axsize;
   assign uc2rb_rd_req_desc_0_attr_reg[27:24] = int_rd_req_desc_0_attr_axsnoop;
   assign uc2rb_rd_req_desc_0_attr_reg[23:22] = int_rd_req_desc_0_attr_axdomain;
   assign uc2rb_rd_req_desc_0_attr_reg[21:20] = int_rd_req_desc_0_attr_axbar;
   assign uc2rb_rd_req_desc_0_attr_reg[18:15] = int_rd_req_desc_0_attr_axregion;
   assign uc2rb_rd_req_desc_0_attr_reg[14:11] = int_rd_req_desc_0_attr_axqos;
   assign uc2rb_rd_req_desc_0_attr_reg[10:8] = int_rd_req_desc_0_attr_axprot;
   assign uc2rb_rd_req_desc_0_attr_reg[7:4] = int_rd_req_desc_0_attr_axcache;
   assign uc2rb_rd_req_desc_0_attr_reg[2] = int_rd_req_desc_0_attr_axlock;
   assign uc2rb_rd_req_desc_0_attr_reg[1:0] = int_rd_req_desc_0_attr_axburst;
   assign uc2rb_rd_req_desc_0_axaddr_0_reg[31:0] = int_rd_req_desc_0_axaddr_0_addr;
   assign uc2rb_rd_req_desc_0_axaddr_1_reg[31:0] = int_rd_req_desc_0_axaddr_1_addr;
   assign uc2rb_rd_req_desc_0_axaddr_2_reg[31:0] = int_rd_req_desc_0_axaddr_2_addr;
   assign uc2rb_rd_req_desc_0_axaddr_3_reg[31:0] = int_rd_req_desc_0_axaddr_3_addr;
   assign uc2rb_rd_req_desc_0_axid_0_reg[31:0] = int_rd_req_desc_0_axid_0_axid;
   assign uc2rb_rd_req_desc_0_axid_1_reg[31:0] = int_rd_req_desc_0_axid_1_axid;
   assign uc2rb_rd_req_desc_0_axid_2_reg[31:0] = int_rd_req_desc_0_axid_2_axid;
   assign uc2rb_rd_req_desc_0_axid_3_reg[31:0] = int_rd_req_desc_0_axid_3_axid;
   assign uc2rb_rd_req_desc_0_axuser_0_reg[31:0] = int_rd_req_desc_0_axuser_0_axuser;
   assign uc2rb_rd_req_desc_0_axuser_1_reg[31:0] = int_rd_req_desc_0_axuser_1_axuser;
   assign uc2rb_rd_req_desc_0_axuser_2_reg[31:0] = int_rd_req_desc_0_axuser_2_axuser;
   assign uc2rb_rd_req_desc_0_axuser_3_reg[31:0] = int_rd_req_desc_0_axuser_3_axuser;
   assign uc2rb_rd_req_desc_0_axuser_4_reg[31:0] = int_rd_req_desc_0_axuser_4_axuser;
   assign uc2rb_rd_req_desc_0_axuser_5_reg[31:0] = int_rd_req_desc_0_axuser_5_axuser;
   assign uc2rb_rd_req_desc_0_axuser_6_reg[31:0] = int_rd_req_desc_0_axuser_6_axuser;
   assign uc2rb_rd_req_desc_0_axuser_7_reg[31:0] = int_rd_req_desc_0_axuser_7_axuser;
   assign uc2rb_rd_req_desc_0_axuser_8_reg[31:0] = int_rd_req_desc_0_axuser_8_axuser;
   assign uc2rb_rd_req_desc_0_axuser_9_reg[31:0] = int_rd_req_desc_0_axuser_9_axuser;
   assign uc2rb_rd_req_desc_0_axuser_10_reg[31:0] = int_rd_req_desc_0_axuser_10_axuser;
   assign uc2rb_rd_req_desc_0_axuser_11_reg[31:0] = int_rd_req_desc_0_axuser_11_axuser;
   assign uc2rb_rd_req_desc_0_axuser_12_reg[31:0] = int_rd_req_desc_0_axuser_12_axuser;
   assign uc2rb_rd_req_desc_0_axuser_13_reg[31:0] = int_rd_req_desc_0_axuser_13_axuser;
   assign uc2rb_rd_req_desc_0_axuser_14_reg[31:0] = int_rd_req_desc_0_axuser_14_axuser;
   assign uc2rb_rd_req_desc_0_axuser_15_reg[31:0] = int_rd_req_desc_0_axuser_15_axuser;
   assign uc2rb_wr_req_desc_0_txn_type_reg[1] = int_wr_req_desc_0_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_0_size_reg[31:0] = int_wr_req_desc_0_size_txn_size;
   assign uc2rb_wr_req_desc_0_data_offset_reg[13:0] = int_wr_req_desc_0_data_offset_addr;
   assign uc2rb_wr_req_desc_0_axsize_reg[2:0] = int_wr_req_desc_0_axsize_axsize;
   assign uc2rb_wr_req_desc_0_attr_reg[27:24] = int_wr_req_desc_0_attr_axsnoop;
   assign uc2rb_wr_req_desc_0_attr_reg[23:22] = int_wr_req_desc_0_attr_axdomain;
   assign uc2rb_wr_req_desc_0_attr_reg[21:20] = int_wr_req_desc_0_attr_axbar;
   assign uc2rb_wr_req_desc_0_attr_reg[19] = int_wr_req_desc_0_attr_awunique;
   assign uc2rb_wr_req_desc_0_attr_reg[18:15] = int_wr_req_desc_0_attr_axregion;
   assign uc2rb_wr_req_desc_0_attr_reg[14:11] = int_wr_req_desc_0_attr_axqos;
   assign uc2rb_wr_req_desc_0_attr_reg[10:8] = int_wr_req_desc_0_attr_axprot;
   assign uc2rb_wr_req_desc_0_attr_reg[7:4] = int_wr_req_desc_0_attr_axcache;
   assign uc2rb_wr_req_desc_0_attr_reg[2] = int_wr_req_desc_0_attr_axlock;
   assign uc2rb_wr_req_desc_0_attr_reg[1:0] = int_wr_req_desc_0_attr_axburst;
   assign uc2rb_wr_req_desc_0_axaddr_0_reg[31:0] = int_wr_req_desc_0_axaddr_0_addr;
   assign uc2rb_wr_req_desc_0_axaddr_1_reg[31:0] = int_wr_req_desc_0_axaddr_1_addr;
   assign uc2rb_wr_req_desc_0_axaddr_2_reg[31:0] = int_wr_req_desc_0_axaddr_2_addr;
   assign uc2rb_wr_req_desc_0_axaddr_3_reg[31:0] = int_wr_req_desc_0_axaddr_3_addr;
   assign uc2rb_wr_req_desc_0_axid_0_reg[31:0] = int_wr_req_desc_0_axid_0_axid;
   assign uc2rb_wr_req_desc_0_axid_1_reg[31:0] = int_wr_req_desc_0_axid_1_axid;
   assign uc2rb_wr_req_desc_0_axid_2_reg[31:0] = int_wr_req_desc_0_axid_2_axid;
   assign uc2rb_wr_req_desc_0_axid_3_reg[31:0] = int_wr_req_desc_0_axid_3_axid;
   assign uc2rb_wr_req_desc_0_axuser_0_reg[31:0] = int_wr_req_desc_0_axuser_0_axuser;
   assign uc2rb_wr_req_desc_0_axuser_1_reg[31:0] = int_wr_req_desc_0_axuser_1_axuser;
   assign uc2rb_wr_req_desc_0_axuser_2_reg[31:0] = int_wr_req_desc_0_axuser_2_axuser;
   assign uc2rb_wr_req_desc_0_axuser_3_reg[31:0] = int_wr_req_desc_0_axuser_3_axuser;
   assign uc2rb_wr_req_desc_0_axuser_4_reg[31:0] = int_wr_req_desc_0_axuser_4_axuser;
   assign uc2rb_wr_req_desc_0_axuser_5_reg[31:0] = int_wr_req_desc_0_axuser_5_axuser;
   assign uc2rb_wr_req_desc_0_axuser_6_reg[31:0] = int_wr_req_desc_0_axuser_6_axuser;
   assign uc2rb_wr_req_desc_0_axuser_7_reg[31:0] = int_wr_req_desc_0_axuser_7_axuser;
   assign uc2rb_wr_req_desc_0_axuser_8_reg[31:0] = int_wr_req_desc_0_axuser_8_axuser;
   assign uc2rb_wr_req_desc_0_axuser_9_reg[31:0] = int_wr_req_desc_0_axuser_9_axuser;
   assign uc2rb_wr_req_desc_0_axuser_10_reg[31:0] = int_wr_req_desc_0_axuser_10_axuser;
   assign uc2rb_wr_req_desc_0_axuser_11_reg[31:0] = int_wr_req_desc_0_axuser_11_axuser;
   assign uc2rb_wr_req_desc_0_axuser_12_reg[31:0] = int_wr_req_desc_0_axuser_12_axuser;
   assign uc2rb_wr_req_desc_0_axuser_13_reg[31:0] = int_wr_req_desc_0_axuser_13_axuser;
   assign uc2rb_wr_req_desc_0_axuser_14_reg[31:0] = int_wr_req_desc_0_axuser_14_axuser;
   assign uc2rb_wr_req_desc_0_axuser_15_reg[31:0] = int_wr_req_desc_0_axuser_15_axuser;
   assign uc2rb_wr_req_desc_0_wuser_0_reg[31:0] = int_wr_req_desc_0_wuser_0_wuser;
   assign uc2rb_wr_req_desc_0_wuser_1_reg[31:0] = int_wr_req_desc_0_wuser_1_wuser;
   assign uc2rb_wr_req_desc_0_wuser_2_reg[31:0] = int_wr_req_desc_0_wuser_2_wuser;
   assign uc2rb_wr_req_desc_0_wuser_3_reg[31:0] = int_wr_req_desc_0_wuser_3_wuser;
   assign uc2rb_wr_req_desc_0_wuser_4_reg[31:0] = int_wr_req_desc_0_wuser_4_wuser;
   assign uc2rb_wr_req_desc_0_wuser_5_reg[31:0] = int_wr_req_desc_0_wuser_5_wuser;
   assign uc2rb_wr_req_desc_0_wuser_6_reg[31:0] = int_wr_req_desc_0_wuser_6_wuser;
   assign uc2rb_wr_req_desc_0_wuser_7_reg[31:0] = int_wr_req_desc_0_wuser_7_wuser;
   assign uc2rb_wr_req_desc_0_wuser_8_reg[31:0] = int_wr_req_desc_0_wuser_8_wuser;
   assign uc2rb_wr_req_desc_0_wuser_9_reg[31:0] = int_wr_req_desc_0_wuser_9_wuser;
   assign uc2rb_wr_req_desc_0_wuser_10_reg[31:0] = int_wr_req_desc_0_wuser_10_wuser;
   assign uc2rb_wr_req_desc_0_wuser_11_reg[31:0] = int_wr_req_desc_0_wuser_11_wuser;
   assign uc2rb_wr_req_desc_0_wuser_12_reg[31:0] = int_wr_req_desc_0_wuser_12_wuser;
   assign uc2rb_wr_req_desc_0_wuser_13_reg[31:0] = int_wr_req_desc_0_wuser_13_wuser;
   assign uc2rb_wr_req_desc_0_wuser_14_reg[31:0] = int_wr_req_desc_0_wuser_14_wuser;
   assign uc2rb_wr_req_desc_0_wuser_15_reg[31:0] = int_wr_req_desc_0_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_0_resp_reg[4:0] = int_sn_resp_desc_0_resp_resp;
   assign uc2rb_rd_req_desc_1_size_reg[31:0] = int_rd_req_desc_1_size_txn_size;
   assign uc2rb_rd_req_desc_1_axsize_reg[2:0] = int_rd_req_desc_1_axsize_axsize;
   assign uc2rb_rd_req_desc_1_attr_reg[27:24] = int_rd_req_desc_1_attr_axsnoop;
   assign uc2rb_rd_req_desc_1_attr_reg[23:22] = int_rd_req_desc_1_attr_axdomain;
   assign uc2rb_rd_req_desc_1_attr_reg[21:20] = int_rd_req_desc_1_attr_axbar;
   assign uc2rb_rd_req_desc_1_attr_reg[18:15] = int_rd_req_desc_1_attr_axregion;
   assign uc2rb_rd_req_desc_1_attr_reg[14:11] = int_rd_req_desc_1_attr_axqos;
   assign uc2rb_rd_req_desc_1_attr_reg[10:8] = int_rd_req_desc_1_attr_axprot;
   assign uc2rb_rd_req_desc_1_attr_reg[7:4] = int_rd_req_desc_1_attr_axcache;
   assign uc2rb_rd_req_desc_1_attr_reg[2] = int_rd_req_desc_1_attr_axlock;
   assign uc2rb_rd_req_desc_1_attr_reg[1:0] = int_rd_req_desc_1_attr_axburst;
   assign uc2rb_rd_req_desc_1_axaddr_0_reg[31:0] = int_rd_req_desc_1_axaddr_0_addr;
   assign uc2rb_rd_req_desc_1_axaddr_1_reg[31:0] = int_rd_req_desc_1_axaddr_1_addr;
   assign uc2rb_rd_req_desc_1_axaddr_2_reg[31:0] = int_rd_req_desc_1_axaddr_2_addr;
   assign uc2rb_rd_req_desc_1_axaddr_3_reg[31:0] = int_rd_req_desc_1_axaddr_3_addr;
   assign uc2rb_rd_req_desc_1_axid_0_reg[31:0] = int_rd_req_desc_1_axid_0_axid;
   assign uc2rb_rd_req_desc_1_axid_1_reg[31:0] = int_rd_req_desc_1_axid_1_axid;
   assign uc2rb_rd_req_desc_1_axid_2_reg[31:0] = int_rd_req_desc_1_axid_2_axid;
   assign uc2rb_rd_req_desc_1_axid_3_reg[31:0] = int_rd_req_desc_1_axid_3_axid;
   assign uc2rb_rd_req_desc_1_axuser_0_reg[31:0] = int_rd_req_desc_1_axuser_0_axuser;
   assign uc2rb_rd_req_desc_1_axuser_1_reg[31:0] = int_rd_req_desc_1_axuser_1_axuser;
   assign uc2rb_rd_req_desc_1_axuser_2_reg[31:0] = int_rd_req_desc_1_axuser_2_axuser;
   assign uc2rb_rd_req_desc_1_axuser_3_reg[31:0] = int_rd_req_desc_1_axuser_3_axuser;
   assign uc2rb_rd_req_desc_1_axuser_4_reg[31:0] = int_rd_req_desc_1_axuser_4_axuser;
   assign uc2rb_rd_req_desc_1_axuser_5_reg[31:0] = int_rd_req_desc_1_axuser_5_axuser;
   assign uc2rb_rd_req_desc_1_axuser_6_reg[31:0] = int_rd_req_desc_1_axuser_6_axuser;
   assign uc2rb_rd_req_desc_1_axuser_7_reg[31:0] = int_rd_req_desc_1_axuser_7_axuser;
   assign uc2rb_rd_req_desc_1_axuser_8_reg[31:0] = int_rd_req_desc_1_axuser_8_axuser;
   assign uc2rb_rd_req_desc_1_axuser_9_reg[31:0] = int_rd_req_desc_1_axuser_9_axuser;
   assign uc2rb_rd_req_desc_1_axuser_10_reg[31:0] = int_rd_req_desc_1_axuser_10_axuser;
   assign uc2rb_rd_req_desc_1_axuser_11_reg[31:0] = int_rd_req_desc_1_axuser_11_axuser;
   assign uc2rb_rd_req_desc_1_axuser_12_reg[31:0] = int_rd_req_desc_1_axuser_12_axuser;
   assign uc2rb_rd_req_desc_1_axuser_13_reg[31:0] = int_rd_req_desc_1_axuser_13_axuser;
   assign uc2rb_rd_req_desc_1_axuser_14_reg[31:0] = int_rd_req_desc_1_axuser_14_axuser;
   assign uc2rb_rd_req_desc_1_axuser_15_reg[31:0] = int_rd_req_desc_1_axuser_15_axuser;
   assign uc2rb_wr_req_desc_1_txn_type_reg[1] = int_wr_req_desc_1_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_1_size_reg[31:0] = int_wr_req_desc_1_size_txn_size;
   assign uc2rb_wr_req_desc_1_data_offset_reg[13:0] = int_wr_req_desc_1_data_offset_addr;
   assign uc2rb_wr_req_desc_1_axsize_reg[2:0] = int_wr_req_desc_1_axsize_axsize;
   assign uc2rb_wr_req_desc_1_attr_reg[27:24] = int_wr_req_desc_1_attr_axsnoop;
   assign uc2rb_wr_req_desc_1_attr_reg[23:22] = int_wr_req_desc_1_attr_axdomain;
   assign uc2rb_wr_req_desc_1_attr_reg[21:20] = int_wr_req_desc_1_attr_axbar;
   assign uc2rb_wr_req_desc_1_attr_reg[19] = int_wr_req_desc_1_attr_awunique;
   assign uc2rb_wr_req_desc_1_attr_reg[18:15] = int_wr_req_desc_1_attr_axregion;
   assign uc2rb_wr_req_desc_1_attr_reg[14:11] = int_wr_req_desc_1_attr_axqos;
   assign uc2rb_wr_req_desc_1_attr_reg[10:8] = int_wr_req_desc_1_attr_axprot;
   assign uc2rb_wr_req_desc_1_attr_reg[7:4] = int_wr_req_desc_1_attr_axcache;
   assign uc2rb_wr_req_desc_1_attr_reg[2] = int_wr_req_desc_1_attr_axlock;
   assign uc2rb_wr_req_desc_1_attr_reg[1:0] = int_wr_req_desc_1_attr_axburst;
   assign uc2rb_wr_req_desc_1_axaddr_0_reg[31:0] = int_wr_req_desc_1_axaddr_0_addr;
   assign uc2rb_wr_req_desc_1_axaddr_1_reg[31:0] = int_wr_req_desc_1_axaddr_1_addr;
   assign uc2rb_wr_req_desc_1_axaddr_2_reg[31:0] = int_wr_req_desc_1_axaddr_2_addr;
   assign uc2rb_wr_req_desc_1_axaddr_3_reg[31:0] = int_wr_req_desc_1_axaddr_3_addr;
   assign uc2rb_wr_req_desc_1_axid_0_reg[31:0] = int_wr_req_desc_1_axid_0_axid;
   assign uc2rb_wr_req_desc_1_axid_1_reg[31:0] = int_wr_req_desc_1_axid_1_axid;
   assign uc2rb_wr_req_desc_1_axid_2_reg[31:0] = int_wr_req_desc_1_axid_2_axid;
   assign uc2rb_wr_req_desc_1_axid_3_reg[31:0] = int_wr_req_desc_1_axid_3_axid;
   assign uc2rb_wr_req_desc_1_axuser_0_reg[31:0] = int_wr_req_desc_1_axuser_0_axuser;
   assign uc2rb_wr_req_desc_1_axuser_1_reg[31:0] = int_wr_req_desc_1_axuser_1_axuser;
   assign uc2rb_wr_req_desc_1_axuser_2_reg[31:0] = int_wr_req_desc_1_axuser_2_axuser;
   assign uc2rb_wr_req_desc_1_axuser_3_reg[31:0] = int_wr_req_desc_1_axuser_3_axuser;
   assign uc2rb_wr_req_desc_1_axuser_4_reg[31:0] = int_wr_req_desc_1_axuser_4_axuser;
   assign uc2rb_wr_req_desc_1_axuser_5_reg[31:0] = int_wr_req_desc_1_axuser_5_axuser;
   assign uc2rb_wr_req_desc_1_axuser_6_reg[31:0] = int_wr_req_desc_1_axuser_6_axuser;
   assign uc2rb_wr_req_desc_1_axuser_7_reg[31:0] = int_wr_req_desc_1_axuser_7_axuser;
   assign uc2rb_wr_req_desc_1_axuser_8_reg[31:0] = int_wr_req_desc_1_axuser_8_axuser;
   assign uc2rb_wr_req_desc_1_axuser_9_reg[31:0] = int_wr_req_desc_1_axuser_9_axuser;
   assign uc2rb_wr_req_desc_1_axuser_10_reg[31:0] = int_wr_req_desc_1_axuser_10_axuser;
   assign uc2rb_wr_req_desc_1_axuser_11_reg[31:0] = int_wr_req_desc_1_axuser_11_axuser;
   assign uc2rb_wr_req_desc_1_axuser_12_reg[31:0] = int_wr_req_desc_1_axuser_12_axuser;
   assign uc2rb_wr_req_desc_1_axuser_13_reg[31:0] = int_wr_req_desc_1_axuser_13_axuser;
   assign uc2rb_wr_req_desc_1_axuser_14_reg[31:0] = int_wr_req_desc_1_axuser_14_axuser;
   assign uc2rb_wr_req_desc_1_axuser_15_reg[31:0] = int_wr_req_desc_1_axuser_15_axuser;
   assign uc2rb_wr_req_desc_1_wuser_0_reg[31:0] = int_wr_req_desc_1_wuser_0_wuser;
   assign uc2rb_wr_req_desc_1_wuser_1_reg[31:0] = int_wr_req_desc_1_wuser_1_wuser;
   assign uc2rb_wr_req_desc_1_wuser_2_reg[31:0] = int_wr_req_desc_1_wuser_2_wuser;
   assign uc2rb_wr_req_desc_1_wuser_3_reg[31:0] = int_wr_req_desc_1_wuser_3_wuser;
   assign uc2rb_wr_req_desc_1_wuser_4_reg[31:0] = int_wr_req_desc_1_wuser_4_wuser;
   assign uc2rb_wr_req_desc_1_wuser_5_reg[31:0] = int_wr_req_desc_1_wuser_5_wuser;
   assign uc2rb_wr_req_desc_1_wuser_6_reg[31:0] = int_wr_req_desc_1_wuser_6_wuser;
   assign uc2rb_wr_req_desc_1_wuser_7_reg[31:0] = int_wr_req_desc_1_wuser_7_wuser;
   assign uc2rb_wr_req_desc_1_wuser_8_reg[31:0] = int_wr_req_desc_1_wuser_8_wuser;
   assign uc2rb_wr_req_desc_1_wuser_9_reg[31:0] = int_wr_req_desc_1_wuser_9_wuser;
   assign uc2rb_wr_req_desc_1_wuser_10_reg[31:0] = int_wr_req_desc_1_wuser_10_wuser;
   assign uc2rb_wr_req_desc_1_wuser_11_reg[31:0] = int_wr_req_desc_1_wuser_11_wuser;
   assign uc2rb_wr_req_desc_1_wuser_12_reg[31:0] = int_wr_req_desc_1_wuser_12_wuser;
   assign uc2rb_wr_req_desc_1_wuser_13_reg[31:0] = int_wr_req_desc_1_wuser_13_wuser;
   assign uc2rb_wr_req_desc_1_wuser_14_reg[31:0] = int_wr_req_desc_1_wuser_14_wuser;
   assign uc2rb_wr_req_desc_1_wuser_15_reg[31:0] = int_wr_req_desc_1_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_1_resp_reg[4:0] = int_sn_resp_desc_1_resp_resp;
   assign uc2rb_rd_req_desc_2_size_reg[31:0] = int_rd_req_desc_2_size_txn_size;
   assign uc2rb_rd_req_desc_2_axsize_reg[2:0] = int_rd_req_desc_2_axsize_axsize;
   assign uc2rb_rd_req_desc_2_attr_reg[27:24] = int_rd_req_desc_2_attr_axsnoop;
   assign uc2rb_rd_req_desc_2_attr_reg[23:22] = int_rd_req_desc_2_attr_axdomain;
   assign uc2rb_rd_req_desc_2_attr_reg[21:20] = int_rd_req_desc_2_attr_axbar;
   assign uc2rb_rd_req_desc_2_attr_reg[18:15] = int_rd_req_desc_2_attr_axregion;
   assign uc2rb_rd_req_desc_2_attr_reg[14:11] = int_rd_req_desc_2_attr_axqos;
   assign uc2rb_rd_req_desc_2_attr_reg[10:8] = int_rd_req_desc_2_attr_axprot;
   assign uc2rb_rd_req_desc_2_attr_reg[7:4] = int_rd_req_desc_2_attr_axcache;
   assign uc2rb_rd_req_desc_2_attr_reg[2] = int_rd_req_desc_2_attr_axlock;
   assign uc2rb_rd_req_desc_2_attr_reg[1:0] = int_rd_req_desc_2_attr_axburst;
   assign uc2rb_rd_req_desc_2_axaddr_0_reg[31:0] = int_rd_req_desc_2_axaddr_0_addr;
   assign uc2rb_rd_req_desc_2_axaddr_1_reg[31:0] = int_rd_req_desc_2_axaddr_1_addr;
   assign uc2rb_rd_req_desc_2_axaddr_2_reg[31:0] = int_rd_req_desc_2_axaddr_2_addr;
   assign uc2rb_rd_req_desc_2_axaddr_3_reg[31:0] = int_rd_req_desc_2_axaddr_3_addr;
   assign uc2rb_rd_req_desc_2_axid_0_reg[31:0] = int_rd_req_desc_2_axid_0_axid;
   assign uc2rb_rd_req_desc_2_axid_1_reg[31:0] = int_rd_req_desc_2_axid_1_axid;
   assign uc2rb_rd_req_desc_2_axid_2_reg[31:0] = int_rd_req_desc_2_axid_2_axid;
   assign uc2rb_rd_req_desc_2_axid_3_reg[31:0] = int_rd_req_desc_2_axid_3_axid;
   assign uc2rb_rd_req_desc_2_axuser_0_reg[31:0] = int_rd_req_desc_2_axuser_0_axuser;
   assign uc2rb_rd_req_desc_2_axuser_1_reg[31:0] = int_rd_req_desc_2_axuser_1_axuser;
   assign uc2rb_rd_req_desc_2_axuser_2_reg[31:0] = int_rd_req_desc_2_axuser_2_axuser;
   assign uc2rb_rd_req_desc_2_axuser_3_reg[31:0] = int_rd_req_desc_2_axuser_3_axuser;
   assign uc2rb_rd_req_desc_2_axuser_4_reg[31:0] = int_rd_req_desc_2_axuser_4_axuser;
   assign uc2rb_rd_req_desc_2_axuser_5_reg[31:0] = int_rd_req_desc_2_axuser_5_axuser;
   assign uc2rb_rd_req_desc_2_axuser_6_reg[31:0] = int_rd_req_desc_2_axuser_6_axuser;
   assign uc2rb_rd_req_desc_2_axuser_7_reg[31:0] = int_rd_req_desc_2_axuser_7_axuser;
   assign uc2rb_rd_req_desc_2_axuser_8_reg[31:0] = int_rd_req_desc_2_axuser_8_axuser;
   assign uc2rb_rd_req_desc_2_axuser_9_reg[31:0] = int_rd_req_desc_2_axuser_9_axuser;
   assign uc2rb_rd_req_desc_2_axuser_10_reg[31:0] = int_rd_req_desc_2_axuser_10_axuser;
   assign uc2rb_rd_req_desc_2_axuser_11_reg[31:0] = int_rd_req_desc_2_axuser_11_axuser;
   assign uc2rb_rd_req_desc_2_axuser_12_reg[31:0] = int_rd_req_desc_2_axuser_12_axuser;
   assign uc2rb_rd_req_desc_2_axuser_13_reg[31:0] = int_rd_req_desc_2_axuser_13_axuser;
   assign uc2rb_rd_req_desc_2_axuser_14_reg[31:0] = int_rd_req_desc_2_axuser_14_axuser;
   assign uc2rb_rd_req_desc_2_axuser_15_reg[31:0] = int_rd_req_desc_2_axuser_15_axuser;
   assign uc2rb_wr_req_desc_2_txn_type_reg[1] = int_wr_req_desc_2_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_2_size_reg[31:0] = int_wr_req_desc_2_size_txn_size;
   assign uc2rb_wr_req_desc_2_data_offset_reg[13:0] = int_wr_req_desc_2_data_offset_addr;
   assign uc2rb_wr_req_desc_2_axsize_reg[2:0] = int_wr_req_desc_2_axsize_axsize;
   assign uc2rb_wr_req_desc_2_attr_reg[27:24] = int_wr_req_desc_2_attr_axsnoop;
   assign uc2rb_wr_req_desc_2_attr_reg[23:22] = int_wr_req_desc_2_attr_axdomain;
   assign uc2rb_wr_req_desc_2_attr_reg[21:20] = int_wr_req_desc_2_attr_axbar;
   assign uc2rb_wr_req_desc_2_attr_reg[19] = int_wr_req_desc_2_attr_awunique;
   assign uc2rb_wr_req_desc_2_attr_reg[18:15] = int_wr_req_desc_2_attr_axregion;
   assign uc2rb_wr_req_desc_2_attr_reg[14:11] = int_wr_req_desc_2_attr_axqos;
   assign uc2rb_wr_req_desc_2_attr_reg[10:8] = int_wr_req_desc_2_attr_axprot;
   assign uc2rb_wr_req_desc_2_attr_reg[7:4] = int_wr_req_desc_2_attr_axcache;
   assign uc2rb_wr_req_desc_2_attr_reg[2] = int_wr_req_desc_2_attr_axlock;
   assign uc2rb_wr_req_desc_2_attr_reg[1:0] = int_wr_req_desc_2_attr_axburst;
   assign uc2rb_wr_req_desc_2_axaddr_0_reg[31:0] = int_wr_req_desc_2_axaddr_0_addr;
   assign uc2rb_wr_req_desc_2_axaddr_1_reg[31:0] = int_wr_req_desc_2_axaddr_1_addr;
   assign uc2rb_wr_req_desc_2_axaddr_2_reg[31:0] = int_wr_req_desc_2_axaddr_2_addr;
   assign uc2rb_wr_req_desc_2_axaddr_3_reg[31:0] = int_wr_req_desc_2_axaddr_3_addr;
   assign uc2rb_wr_req_desc_2_axid_0_reg[31:0] = int_wr_req_desc_2_axid_0_axid;
   assign uc2rb_wr_req_desc_2_axid_1_reg[31:0] = int_wr_req_desc_2_axid_1_axid;
   assign uc2rb_wr_req_desc_2_axid_2_reg[31:0] = int_wr_req_desc_2_axid_2_axid;
   assign uc2rb_wr_req_desc_2_axid_3_reg[31:0] = int_wr_req_desc_2_axid_3_axid;
   assign uc2rb_wr_req_desc_2_axuser_0_reg[31:0] = int_wr_req_desc_2_axuser_0_axuser;
   assign uc2rb_wr_req_desc_2_axuser_1_reg[31:0] = int_wr_req_desc_2_axuser_1_axuser;
   assign uc2rb_wr_req_desc_2_axuser_2_reg[31:0] = int_wr_req_desc_2_axuser_2_axuser;
   assign uc2rb_wr_req_desc_2_axuser_3_reg[31:0] = int_wr_req_desc_2_axuser_3_axuser;
   assign uc2rb_wr_req_desc_2_axuser_4_reg[31:0] = int_wr_req_desc_2_axuser_4_axuser;
   assign uc2rb_wr_req_desc_2_axuser_5_reg[31:0] = int_wr_req_desc_2_axuser_5_axuser;
   assign uc2rb_wr_req_desc_2_axuser_6_reg[31:0] = int_wr_req_desc_2_axuser_6_axuser;
   assign uc2rb_wr_req_desc_2_axuser_7_reg[31:0] = int_wr_req_desc_2_axuser_7_axuser;
   assign uc2rb_wr_req_desc_2_axuser_8_reg[31:0] = int_wr_req_desc_2_axuser_8_axuser;
   assign uc2rb_wr_req_desc_2_axuser_9_reg[31:0] = int_wr_req_desc_2_axuser_9_axuser;
   assign uc2rb_wr_req_desc_2_axuser_10_reg[31:0] = int_wr_req_desc_2_axuser_10_axuser;
   assign uc2rb_wr_req_desc_2_axuser_11_reg[31:0] = int_wr_req_desc_2_axuser_11_axuser;
   assign uc2rb_wr_req_desc_2_axuser_12_reg[31:0] = int_wr_req_desc_2_axuser_12_axuser;
   assign uc2rb_wr_req_desc_2_axuser_13_reg[31:0] = int_wr_req_desc_2_axuser_13_axuser;
   assign uc2rb_wr_req_desc_2_axuser_14_reg[31:0] = int_wr_req_desc_2_axuser_14_axuser;
   assign uc2rb_wr_req_desc_2_axuser_15_reg[31:0] = int_wr_req_desc_2_axuser_15_axuser;
   assign uc2rb_wr_req_desc_2_wuser_0_reg[31:0] = int_wr_req_desc_2_wuser_0_wuser;
   assign uc2rb_wr_req_desc_2_wuser_1_reg[31:0] = int_wr_req_desc_2_wuser_1_wuser;
   assign uc2rb_wr_req_desc_2_wuser_2_reg[31:0] = int_wr_req_desc_2_wuser_2_wuser;
   assign uc2rb_wr_req_desc_2_wuser_3_reg[31:0] = int_wr_req_desc_2_wuser_3_wuser;
   assign uc2rb_wr_req_desc_2_wuser_4_reg[31:0] = int_wr_req_desc_2_wuser_4_wuser;
   assign uc2rb_wr_req_desc_2_wuser_5_reg[31:0] = int_wr_req_desc_2_wuser_5_wuser;
   assign uc2rb_wr_req_desc_2_wuser_6_reg[31:0] = int_wr_req_desc_2_wuser_6_wuser;
   assign uc2rb_wr_req_desc_2_wuser_7_reg[31:0] = int_wr_req_desc_2_wuser_7_wuser;
   assign uc2rb_wr_req_desc_2_wuser_8_reg[31:0] = int_wr_req_desc_2_wuser_8_wuser;
   assign uc2rb_wr_req_desc_2_wuser_9_reg[31:0] = int_wr_req_desc_2_wuser_9_wuser;
   assign uc2rb_wr_req_desc_2_wuser_10_reg[31:0] = int_wr_req_desc_2_wuser_10_wuser;
   assign uc2rb_wr_req_desc_2_wuser_11_reg[31:0] = int_wr_req_desc_2_wuser_11_wuser;
   assign uc2rb_wr_req_desc_2_wuser_12_reg[31:0] = int_wr_req_desc_2_wuser_12_wuser;
   assign uc2rb_wr_req_desc_2_wuser_13_reg[31:0] = int_wr_req_desc_2_wuser_13_wuser;
   assign uc2rb_wr_req_desc_2_wuser_14_reg[31:0] = int_wr_req_desc_2_wuser_14_wuser;
   assign uc2rb_wr_req_desc_2_wuser_15_reg[31:0] = int_wr_req_desc_2_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_2_resp_reg[4:0] = int_sn_resp_desc_2_resp_resp;
   assign uc2rb_rd_req_desc_3_size_reg[31:0] = int_rd_req_desc_3_size_txn_size;
   assign uc2rb_rd_req_desc_3_axsize_reg[2:0] = int_rd_req_desc_3_axsize_axsize;
   assign uc2rb_rd_req_desc_3_attr_reg[27:24] = int_rd_req_desc_3_attr_axsnoop;
   assign uc2rb_rd_req_desc_3_attr_reg[23:22] = int_rd_req_desc_3_attr_axdomain;
   assign uc2rb_rd_req_desc_3_attr_reg[21:20] = int_rd_req_desc_3_attr_axbar;
   assign uc2rb_rd_req_desc_3_attr_reg[18:15] = int_rd_req_desc_3_attr_axregion;
   assign uc2rb_rd_req_desc_3_attr_reg[14:11] = int_rd_req_desc_3_attr_axqos;
   assign uc2rb_rd_req_desc_3_attr_reg[10:8] = int_rd_req_desc_3_attr_axprot;
   assign uc2rb_rd_req_desc_3_attr_reg[7:4] = int_rd_req_desc_3_attr_axcache;
   assign uc2rb_rd_req_desc_3_attr_reg[2] = int_rd_req_desc_3_attr_axlock;
   assign uc2rb_rd_req_desc_3_attr_reg[1:0] = int_rd_req_desc_3_attr_axburst;
   assign uc2rb_rd_req_desc_3_axaddr_0_reg[31:0] = int_rd_req_desc_3_axaddr_0_addr;
   assign uc2rb_rd_req_desc_3_axaddr_1_reg[31:0] = int_rd_req_desc_3_axaddr_1_addr;
   assign uc2rb_rd_req_desc_3_axaddr_2_reg[31:0] = int_rd_req_desc_3_axaddr_2_addr;
   assign uc2rb_rd_req_desc_3_axaddr_3_reg[31:0] = int_rd_req_desc_3_axaddr_3_addr;
   assign uc2rb_rd_req_desc_3_axid_0_reg[31:0] = int_rd_req_desc_3_axid_0_axid;
   assign uc2rb_rd_req_desc_3_axid_1_reg[31:0] = int_rd_req_desc_3_axid_1_axid;
   assign uc2rb_rd_req_desc_3_axid_2_reg[31:0] = int_rd_req_desc_3_axid_2_axid;
   assign uc2rb_rd_req_desc_3_axid_3_reg[31:0] = int_rd_req_desc_3_axid_3_axid;
   assign uc2rb_rd_req_desc_3_axuser_0_reg[31:0] = int_rd_req_desc_3_axuser_0_axuser;
   assign uc2rb_rd_req_desc_3_axuser_1_reg[31:0] = int_rd_req_desc_3_axuser_1_axuser;
   assign uc2rb_rd_req_desc_3_axuser_2_reg[31:0] = int_rd_req_desc_3_axuser_2_axuser;
   assign uc2rb_rd_req_desc_3_axuser_3_reg[31:0] = int_rd_req_desc_3_axuser_3_axuser;
   assign uc2rb_rd_req_desc_3_axuser_4_reg[31:0] = int_rd_req_desc_3_axuser_4_axuser;
   assign uc2rb_rd_req_desc_3_axuser_5_reg[31:0] = int_rd_req_desc_3_axuser_5_axuser;
   assign uc2rb_rd_req_desc_3_axuser_6_reg[31:0] = int_rd_req_desc_3_axuser_6_axuser;
   assign uc2rb_rd_req_desc_3_axuser_7_reg[31:0] = int_rd_req_desc_3_axuser_7_axuser;
   assign uc2rb_rd_req_desc_3_axuser_8_reg[31:0] = int_rd_req_desc_3_axuser_8_axuser;
   assign uc2rb_rd_req_desc_3_axuser_9_reg[31:0] = int_rd_req_desc_3_axuser_9_axuser;
   assign uc2rb_rd_req_desc_3_axuser_10_reg[31:0] = int_rd_req_desc_3_axuser_10_axuser;
   assign uc2rb_rd_req_desc_3_axuser_11_reg[31:0] = int_rd_req_desc_3_axuser_11_axuser;
   assign uc2rb_rd_req_desc_3_axuser_12_reg[31:0] = int_rd_req_desc_3_axuser_12_axuser;
   assign uc2rb_rd_req_desc_3_axuser_13_reg[31:0] = int_rd_req_desc_3_axuser_13_axuser;
   assign uc2rb_rd_req_desc_3_axuser_14_reg[31:0] = int_rd_req_desc_3_axuser_14_axuser;
   assign uc2rb_rd_req_desc_3_axuser_15_reg[31:0] = int_rd_req_desc_3_axuser_15_axuser;
   assign uc2rb_wr_req_desc_3_txn_type_reg[1] = int_wr_req_desc_3_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_3_size_reg[31:0] = int_wr_req_desc_3_size_txn_size;
   assign uc2rb_wr_req_desc_3_data_offset_reg[13:0] = int_wr_req_desc_3_data_offset_addr;
   assign uc2rb_wr_req_desc_3_axsize_reg[2:0] = int_wr_req_desc_3_axsize_axsize;
   assign uc2rb_wr_req_desc_3_attr_reg[27:24] = int_wr_req_desc_3_attr_axsnoop;
   assign uc2rb_wr_req_desc_3_attr_reg[23:22] = int_wr_req_desc_3_attr_axdomain;
   assign uc2rb_wr_req_desc_3_attr_reg[21:20] = int_wr_req_desc_3_attr_axbar;
   assign uc2rb_wr_req_desc_3_attr_reg[19] = int_wr_req_desc_3_attr_awunique;
   assign uc2rb_wr_req_desc_3_attr_reg[18:15] = int_wr_req_desc_3_attr_axregion;
   assign uc2rb_wr_req_desc_3_attr_reg[14:11] = int_wr_req_desc_3_attr_axqos;
   assign uc2rb_wr_req_desc_3_attr_reg[10:8] = int_wr_req_desc_3_attr_axprot;
   assign uc2rb_wr_req_desc_3_attr_reg[7:4] = int_wr_req_desc_3_attr_axcache;
   assign uc2rb_wr_req_desc_3_attr_reg[2] = int_wr_req_desc_3_attr_axlock;
   assign uc2rb_wr_req_desc_3_attr_reg[1:0] = int_wr_req_desc_3_attr_axburst;
   assign uc2rb_wr_req_desc_3_axaddr_0_reg[31:0] = int_wr_req_desc_3_axaddr_0_addr;
   assign uc2rb_wr_req_desc_3_axaddr_1_reg[31:0] = int_wr_req_desc_3_axaddr_1_addr;
   assign uc2rb_wr_req_desc_3_axaddr_2_reg[31:0] = int_wr_req_desc_3_axaddr_2_addr;
   assign uc2rb_wr_req_desc_3_axaddr_3_reg[31:0] = int_wr_req_desc_3_axaddr_3_addr;
   assign uc2rb_wr_req_desc_3_axid_0_reg[31:0] = int_wr_req_desc_3_axid_0_axid;
   assign uc2rb_wr_req_desc_3_axid_1_reg[31:0] = int_wr_req_desc_3_axid_1_axid;
   assign uc2rb_wr_req_desc_3_axid_2_reg[31:0] = int_wr_req_desc_3_axid_2_axid;
   assign uc2rb_wr_req_desc_3_axid_3_reg[31:0] = int_wr_req_desc_3_axid_3_axid;
   assign uc2rb_wr_req_desc_3_axuser_0_reg[31:0] = int_wr_req_desc_3_axuser_0_axuser;
   assign uc2rb_wr_req_desc_3_axuser_1_reg[31:0] = int_wr_req_desc_3_axuser_1_axuser;
   assign uc2rb_wr_req_desc_3_axuser_2_reg[31:0] = int_wr_req_desc_3_axuser_2_axuser;
   assign uc2rb_wr_req_desc_3_axuser_3_reg[31:0] = int_wr_req_desc_3_axuser_3_axuser;
   assign uc2rb_wr_req_desc_3_axuser_4_reg[31:0] = int_wr_req_desc_3_axuser_4_axuser;
   assign uc2rb_wr_req_desc_3_axuser_5_reg[31:0] = int_wr_req_desc_3_axuser_5_axuser;
   assign uc2rb_wr_req_desc_3_axuser_6_reg[31:0] = int_wr_req_desc_3_axuser_6_axuser;
   assign uc2rb_wr_req_desc_3_axuser_7_reg[31:0] = int_wr_req_desc_3_axuser_7_axuser;
   assign uc2rb_wr_req_desc_3_axuser_8_reg[31:0] = int_wr_req_desc_3_axuser_8_axuser;
   assign uc2rb_wr_req_desc_3_axuser_9_reg[31:0] = int_wr_req_desc_3_axuser_9_axuser;
   assign uc2rb_wr_req_desc_3_axuser_10_reg[31:0] = int_wr_req_desc_3_axuser_10_axuser;
   assign uc2rb_wr_req_desc_3_axuser_11_reg[31:0] = int_wr_req_desc_3_axuser_11_axuser;
   assign uc2rb_wr_req_desc_3_axuser_12_reg[31:0] = int_wr_req_desc_3_axuser_12_axuser;
   assign uc2rb_wr_req_desc_3_axuser_13_reg[31:0] = int_wr_req_desc_3_axuser_13_axuser;
   assign uc2rb_wr_req_desc_3_axuser_14_reg[31:0] = int_wr_req_desc_3_axuser_14_axuser;
   assign uc2rb_wr_req_desc_3_axuser_15_reg[31:0] = int_wr_req_desc_3_axuser_15_axuser;
   assign uc2rb_wr_req_desc_3_wuser_0_reg[31:0] = int_wr_req_desc_3_wuser_0_wuser;
   assign uc2rb_wr_req_desc_3_wuser_1_reg[31:0] = int_wr_req_desc_3_wuser_1_wuser;
   assign uc2rb_wr_req_desc_3_wuser_2_reg[31:0] = int_wr_req_desc_3_wuser_2_wuser;
   assign uc2rb_wr_req_desc_3_wuser_3_reg[31:0] = int_wr_req_desc_3_wuser_3_wuser;
   assign uc2rb_wr_req_desc_3_wuser_4_reg[31:0] = int_wr_req_desc_3_wuser_4_wuser;
   assign uc2rb_wr_req_desc_3_wuser_5_reg[31:0] = int_wr_req_desc_3_wuser_5_wuser;
   assign uc2rb_wr_req_desc_3_wuser_6_reg[31:0] = int_wr_req_desc_3_wuser_6_wuser;
   assign uc2rb_wr_req_desc_3_wuser_7_reg[31:0] = int_wr_req_desc_3_wuser_7_wuser;
   assign uc2rb_wr_req_desc_3_wuser_8_reg[31:0] = int_wr_req_desc_3_wuser_8_wuser;
   assign uc2rb_wr_req_desc_3_wuser_9_reg[31:0] = int_wr_req_desc_3_wuser_9_wuser;
   assign uc2rb_wr_req_desc_3_wuser_10_reg[31:0] = int_wr_req_desc_3_wuser_10_wuser;
   assign uc2rb_wr_req_desc_3_wuser_11_reg[31:0] = int_wr_req_desc_3_wuser_11_wuser;
   assign uc2rb_wr_req_desc_3_wuser_12_reg[31:0] = int_wr_req_desc_3_wuser_12_wuser;
   assign uc2rb_wr_req_desc_3_wuser_13_reg[31:0] = int_wr_req_desc_3_wuser_13_wuser;
   assign uc2rb_wr_req_desc_3_wuser_14_reg[31:0] = int_wr_req_desc_3_wuser_14_wuser;
   assign uc2rb_wr_req_desc_3_wuser_15_reg[31:0] = int_wr_req_desc_3_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_3_resp_reg[4:0] = int_sn_resp_desc_3_resp_resp;
   assign uc2rb_rd_req_desc_4_size_reg[31:0] = int_rd_req_desc_4_size_txn_size;
   assign uc2rb_rd_req_desc_4_axsize_reg[2:0] = int_rd_req_desc_4_axsize_axsize;
   assign uc2rb_rd_req_desc_4_attr_reg[27:24] = int_rd_req_desc_4_attr_axsnoop;
   assign uc2rb_rd_req_desc_4_attr_reg[23:22] = int_rd_req_desc_4_attr_axdomain;
   assign uc2rb_rd_req_desc_4_attr_reg[21:20] = int_rd_req_desc_4_attr_axbar;
   assign uc2rb_rd_req_desc_4_attr_reg[18:15] = int_rd_req_desc_4_attr_axregion;
   assign uc2rb_rd_req_desc_4_attr_reg[14:11] = int_rd_req_desc_4_attr_axqos;
   assign uc2rb_rd_req_desc_4_attr_reg[10:8] = int_rd_req_desc_4_attr_axprot;
   assign uc2rb_rd_req_desc_4_attr_reg[7:4] = int_rd_req_desc_4_attr_axcache;
   assign uc2rb_rd_req_desc_4_attr_reg[2] = int_rd_req_desc_4_attr_axlock;
   assign uc2rb_rd_req_desc_4_attr_reg[1:0] = int_rd_req_desc_4_attr_axburst;
   assign uc2rb_rd_req_desc_4_axaddr_0_reg[31:0] = int_rd_req_desc_4_axaddr_0_addr;
   assign uc2rb_rd_req_desc_4_axaddr_1_reg[31:0] = int_rd_req_desc_4_axaddr_1_addr;
   assign uc2rb_rd_req_desc_4_axaddr_2_reg[31:0] = int_rd_req_desc_4_axaddr_2_addr;
   assign uc2rb_rd_req_desc_4_axaddr_3_reg[31:0] = int_rd_req_desc_4_axaddr_3_addr;
   assign uc2rb_rd_req_desc_4_axid_0_reg[31:0] = int_rd_req_desc_4_axid_0_axid;
   assign uc2rb_rd_req_desc_4_axid_1_reg[31:0] = int_rd_req_desc_4_axid_1_axid;
   assign uc2rb_rd_req_desc_4_axid_2_reg[31:0] = int_rd_req_desc_4_axid_2_axid;
   assign uc2rb_rd_req_desc_4_axid_3_reg[31:0] = int_rd_req_desc_4_axid_3_axid;
   assign uc2rb_rd_req_desc_4_axuser_0_reg[31:0] = int_rd_req_desc_4_axuser_0_axuser;
   assign uc2rb_rd_req_desc_4_axuser_1_reg[31:0] = int_rd_req_desc_4_axuser_1_axuser;
   assign uc2rb_rd_req_desc_4_axuser_2_reg[31:0] = int_rd_req_desc_4_axuser_2_axuser;
   assign uc2rb_rd_req_desc_4_axuser_3_reg[31:0] = int_rd_req_desc_4_axuser_3_axuser;
   assign uc2rb_rd_req_desc_4_axuser_4_reg[31:0] = int_rd_req_desc_4_axuser_4_axuser;
   assign uc2rb_rd_req_desc_4_axuser_5_reg[31:0] = int_rd_req_desc_4_axuser_5_axuser;
   assign uc2rb_rd_req_desc_4_axuser_6_reg[31:0] = int_rd_req_desc_4_axuser_6_axuser;
   assign uc2rb_rd_req_desc_4_axuser_7_reg[31:0] = int_rd_req_desc_4_axuser_7_axuser;
   assign uc2rb_rd_req_desc_4_axuser_8_reg[31:0] = int_rd_req_desc_4_axuser_8_axuser;
   assign uc2rb_rd_req_desc_4_axuser_9_reg[31:0] = int_rd_req_desc_4_axuser_9_axuser;
   assign uc2rb_rd_req_desc_4_axuser_10_reg[31:0] = int_rd_req_desc_4_axuser_10_axuser;
   assign uc2rb_rd_req_desc_4_axuser_11_reg[31:0] = int_rd_req_desc_4_axuser_11_axuser;
   assign uc2rb_rd_req_desc_4_axuser_12_reg[31:0] = int_rd_req_desc_4_axuser_12_axuser;
   assign uc2rb_rd_req_desc_4_axuser_13_reg[31:0] = int_rd_req_desc_4_axuser_13_axuser;
   assign uc2rb_rd_req_desc_4_axuser_14_reg[31:0] = int_rd_req_desc_4_axuser_14_axuser;
   assign uc2rb_rd_req_desc_4_axuser_15_reg[31:0] = int_rd_req_desc_4_axuser_15_axuser;
   assign uc2rb_wr_req_desc_4_txn_type_reg[1] = int_wr_req_desc_4_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_4_size_reg[31:0] = int_wr_req_desc_4_size_txn_size;
   assign uc2rb_wr_req_desc_4_data_offset_reg[13:0] = int_wr_req_desc_4_data_offset_addr;
   assign uc2rb_wr_req_desc_4_axsize_reg[2:0] = int_wr_req_desc_4_axsize_axsize;
   assign uc2rb_wr_req_desc_4_attr_reg[27:24] = int_wr_req_desc_4_attr_axsnoop;
   assign uc2rb_wr_req_desc_4_attr_reg[23:22] = int_wr_req_desc_4_attr_axdomain;
   assign uc2rb_wr_req_desc_4_attr_reg[21:20] = int_wr_req_desc_4_attr_axbar;
   assign uc2rb_wr_req_desc_4_attr_reg[19] = int_wr_req_desc_4_attr_awunique;
   assign uc2rb_wr_req_desc_4_attr_reg[18:15] = int_wr_req_desc_4_attr_axregion;
   assign uc2rb_wr_req_desc_4_attr_reg[14:11] = int_wr_req_desc_4_attr_axqos;
   assign uc2rb_wr_req_desc_4_attr_reg[10:8] = int_wr_req_desc_4_attr_axprot;
   assign uc2rb_wr_req_desc_4_attr_reg[7:4] = int_wr_req_desc_4_attr_axcache;
   assign uc2rb_wr_req_desc_4_attr_reg[2] = int_wr_req_desc_4_attr_axlock;
   assign uc2rb_wr_req_desc_4_attr_reg[1:0] = int_wr_req_desc_4_attr_axburst;
   assign uc2rb_wr_req_desc_4_axaddr_0_reg[31:0] = int_wr_req_desc_4_axaddr_0_addr;
   assign uc2rb_wr_req_desc_4_axaddr_1_reg[31:0] = int_wr_req_desc_4_axaddr_1_addr;
   assign uc2rb_wr_req_desc_4_axaddr_2_reg[31:0] = int_wr_req_desc_4_axaddr_2_addr;
   assign uc2rb_wr_req_desc_4_axaddr_3_reg[31:0] = int_wr_req_desc_4_axaddr_3_addr;
   assign uc2rb_wr_req_desc_4_axid_0_reg[31:0] = int_wr_req_desc_4_axid_0_axid;
   assign uc2rb_wr_req_desc_4_axid_1_reg[31:0] = int_wr_req_desc_4_axid_1_axid;
   assign uc2rb_wr_req_desc_4_axid_2_reg[31:0] = int_wr_req_desc_4_axid_2_axid;
   assign uc2rb_wr_req_desc_4_axid_3_reg[31:0] = int_wr_req_desc_4_axid_3_axid;
   assign uc2rb_wr_req_desc_4_axuser_0_reg[31:0] = int_wr_req_desc_4_axuser_0_axuser;
   assign uc2rb_wr_req_desc_4_axuser_1_reg[31:0] = int_wr_req_desc_4_axuser_1_axuser;
   assign uc2rb_wr_req_desc_4_axuser_2_reg[31:0] = int_wr_req_desc_4_axuser_2_axuser;
   assign uc2rb_wr_req_desc_4_axuser_3_reg[31:0] = int_wr_req_desc_4_axuser_3_axuser;
   assign uc2rb_wr_req_desc_4_axuser_4_reg[31:0] = int_wr_req_desc_4_axuser_4_axuser;
   assign uc2rb_wr_req_desc_4_axuser_5_reg[31:0] = int_wr_req_desc_4_axuser_5_axuser;
   assign uc2rb_wr_req_desc_4_axuser_6_reg[31:0] = int_wr_req_desc_4_axuser_6_axuser;
   assign uc2rb_wr_req_desc_4_axuser_7_reg[31:0] = int_wr_req_desc_4_axuser_7_axuser;
   assign uc2rb_wr_req_desc_4_axuser_8_reg[31:0] = int_wr_req_desc_4_axuser_8_axuser;
   assign uc2rb_wr_req_desc_4_axuser_9_reg[31:0] = int_wr_req_desc_4_axuser_9_axuser;
   assign uc2rb_wr_req_desc_4_axuser_10_reg[31:0] = int_wr_req_desc_4_axuser_10_axuser;
   assign uc2rb_wr_req_desc_4_axuser_11_reg[31:0] = int_wr_req_desc_4_axuser_11_axuser;
   assign uc2rb_wr_req_desc_4_axuser_12_reg[31:0] = int_wr_req_desc_4_axuser_12_axuser;
   assign uc2rb_wr_req_desc_4_axuser_13_reg[31:0] = int_wr_req_desc_4_axuser_13_axuser;
   assign uc2rb_wr_req_desc_4_axuser_14_reg[31:0] = int_wr_req_desc_4_axuser_14_axuser;
   assign uc2rb_wr_req_desc_4_axuser_15_reg[31:0] = int_wr_req_desc_4_axuser_15_axuser;
   assign uc2rb_wr_req_desc_4_wuser_0_reg[31:0] = int_wr_req_desc_4_wuser_0_wuser;
   assign uc2rb_wr_req_desc_4_wuser_1_reg[31:0] = int_wr_req_desc_4_wuser_1_wuser;
   assign uc2rb_wr_req_desc_4_wuser_2_reg[31:0] = int_wr_req_desc_4_wuser_2_wuser;
   assign uc2rb_wr_req_desc_4_wuser_3_reg[31:0] = int_wr_req_desc_4_wuser_3_wuser;
   assign uc2rb_wr_req_desc_4_wuser_4_reg[31:0] = int_wr_req_desc_4_wuser_4_wuser;
   assign uc2rb_wr_req_desc_4_wuser_5_reg[31:0] = int_wr_req_desc_4_wuser_5_wuser;
   assign uc2rb_wr_req_desc_4_wuser_6_reg[31:0] = int_wr_req_desc_4_wuser_6_wuser;
   assign uc2rb_wr_req_desc_4_wuser_7_reg[31:0] = int_wr_req_desc_4_wuser_7_wuser;
   assign uc2rb_wr_req_desc_4_wuser_8_reg[31:0] = int_wr_req_desc_4_wuser_8_wuser;
   assign uc2rb_wr_req_desc_4_wuser_9_reg[31:0] = int_wr_req_desc_4_wuser_9_wuser;
   assign uc2rb_wr_req_desc_4_wuser_10_reg[31:0] = int_wr_req_desc_4_wuser_10_wuser;
   assign uc2rb_wr_req_desc_4_wuser_11_reg[31:0] = int_wr_req_desc_4_wuser_11_wuser;
   assign uc2rb_wr_req_desc_4_wuser_12_reg[31:0] = int_wr_req_desc_4_wuser_12_wuser;
   assign uc2rb_wr_req_desc_4_wuser_13_reg[31:0] = int_wr_req_desc_4_wuser_13_wuser;
   assign uc2rb_wr_req_desc_4_wuser_14_reg[31:0] = int_wr_req_desc_4_wuser_14_wuser;
   assign uc2rb_wr_req_desc_4_wuser_15_reg[31:0] = int_wr_req_desc_4_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_4_resp_reg[4:0] = int_sn_resp_desc_4_resp_resp;
   assign uc2rb_rd_req_desc_5_size_reg[31:0] = int_rd_req_desc_5_size_txn_size;
   assign uc2rb_rd_req_desc_5_axsize_reg[2:0] = int_rd_req_desc_5_axsize_axsize;
   assign uc2rb_rd_req_desc_5_attr_reg[27:24] = int_rd_req_desc_5_attr_axsnoop;
   assign uc2rb_rd_req_desc_5_attr_reg[23:22] = int_rd_req_desc_5_attr_axdomain;
   assign uc2rb_rd_req_desc_5_attr_reg[21:20] = int_rd_req_desc_5_attr_axbar;
   assign uc2rb_rd_req_desc_5_attr_reg[18:15] = int_rd_req_desc_5_attr_axregion;
   assign uc2rb_rd_req_desc_5_attr_reg[14:11] = int_rd_req_desc_5_attr_axqos;
   assign uc2rb_rd_req_desc_5_attr_reg[10:8] = int_rd_req_desc_5_attr_axprot;
   assign uc2rb_rd_req_desc_5_attr_reg[7:4] = int_rd_req_desc_5_attr_axcache;
   assign uc2rb_rd_req_desc_5_attr_reg[2] = int_rd_req_desc_5_attr_axlock;
   assign uc2rb_rd_req_desc_5_attr_reg[1:0] = int_rd_req_desc_5_attr_axburst;
   assign uc2rb_rd_req_desc_5_axaddr_0_reg[31:0] = int_rd_req_desc_5_axaddr_0_addr;
   assign uc2rb_rd_req_desc_5_axaddr_1_reg[31:0] = int_rd_req_desc_5_axaddr_1_addr;
   assign uc2rb_rd_req_desc_5_axaddr_2_reg[31:0] = int_rd_req_desc_5_axaddr_2_addr;
   assign uc2rb_rd_req_desc_5_axaddr_3_reg[31:0] = int_rd_req_desc_5_axaddr_3_addr;
   assign uc2rb_rd_req_desc_5_axid_0_reg[31:0] = int_rd_req_desc_5_axid_0_axid;
   assign uc2rb_rd_req_desc_5_axid_1_reg[31:0] = int_rd_req_desc_5_axid_1_axid;
   assign uc2rb_rd_req_desc_5_axid_2_reg[31:0] = int_rd_req_desc_5_axid_2_axid;
   assign uc2rb_rd_req_desc_5_axid_3_reg[31:0] = int_rd_req_desc_5_axid_3_axid;
   assign uc2rb_rd_req_desc_5_axuser_0_reg[31:0] = int_rd_req_desc_5_axuser_0_axuser;
   assign uc2rb_rd_req_desc_5_axuser_1_reg[31:0] = int_rd_req_desc_5_axuser_1_axuser;
   assign uc2rb_rd_req_desc_5_axuser_2_reg[31:0] = int_rd_req_desc_5_axuser_2_axuser;
   assign uc2rb_rd_req_desc_5_axuser_3_reg[31:0] = int_rd_req_desc_5_axuser_3_axuser;
   assign uc2rb_rd_req_desc_5_axuser_4_reg[31:0] = int_rd_req_desc_5_axuser_4_axuser;
   assign uc2rb_rd_req_desc_5_axuser_5_reg[31:0] = int_rd_req_desc_5_axuser_5_axuser;
   assign uc2rb_rd_req_desc_5_axuser_6_reg[31:0] = int_rd_req_desc_5_axuser_6_axuser;
   assign uc2rb_rd_req_desc_5_axuser_7_reg[31:0] = int_rd_req_desc_5_axuser_7_axuser;
   assign uc2rb_rd_req_desc_5_axuser_8_reg[31:0] = int_rd_req_desc_5_axuser_8_axuser;
   assign uc2rb_rd_req_desc_5_axuser_9_reg[31:0] = int_rd_req_desc_5_axuser_9_axuser;
   assign uc2rb_rd_req_desc_5_axuser_10_reg[31:0] = int_rd_req_desc_5_axuser_10_axuser;
   assign uc2rb_rd_req_desc_5_axuser_11_reg[31:0] = int_rd_req_desc_5_axuser_11_axuser;
   assign uc2rb_rd_req_desc_5_axuser_12_reg[31:0] = int_rd_req_desc_5_axuser_12_axuser;
   assign uc2rb_rd_req_desc_5_axuser_13_reg[31:0] = int_rd_req_desc_5_axuser_13_axuser;
   assign uc2rb_rd_req_desc_5_axuser_14_reg[31:0] = int_rd_req_desc_5_axuser_14_axuser;
   assign uc2rb_rd_req_desc_5_axuser_15_reg[31:0] = int_rd_req_desc_5_axuser_15_axuser;
   assign uc2rb_wr_req_desc_5_txn_type_reg[1] = int_wr_req_desc_5_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_5_size_reg[31:0] = int_wr_req_desc_5_size_txn_size;
   assign uc2rb_wr_req_desc_5_data_offset_reg[13:0] = int_wr_req_desc_5_data_offset_addr;
   assign uc2rb_wr_req_desc_5_axsize_reg[2:0] = int_wr_req_desc_5_axsize_axsize;
   assign uc2rb_wr_req_desc_5_attr_reg[27:24] = int_wr_req_desc_5_attr_axsnoop;
   assign uc2rb_wr_req_desc_5_attr_reg[23:22] = int_wr_req_desc_5_attr_axdomain;
   assign uc2rb_wr_req_desc_5_attr_reg[21:20] = int_wr_req_desc_5_attr_axbar;
   assign uc2rb_wr_req_desc_5_attr_reg[19] = int_wr_req_desc_5_attr_awunique;
   assign uc2rb_wr_req_desc_5_attr_reg[18:15] = int_wr_req_desc_5_attr_axregion;
   assign uc2rb_wr_req_desc_5_attr_reg[14:11] = int_wr_req_desc_5_attr_axqos;
   assign uc2rb_wr_req_desc_5_attr_reg[10:8] = int_wr_req_desc_5_attr_axprot;
   assign uc2rb_wr_req_desc_5_attr_reg[7:4] = int_wr_req_desc_5_attr_axcache;
   assign uc2rb_wr_req_desc_5_attr_reg[2] = int_wr_req_desc_5_attr_axlock;
   assign uc2rb_wr_req_desc_5_attr_reg[1:0] = int_wr_req_desc_5_attr_axburst;
   assign uc2rb_wr_req_desc_5_axaddr_0_reg[31:0] = int_wr_req_desc_5_axaddr_0_addr;
   assign uc2rb_wr_req_desc_5_axaddr_1_reg[31:0] = int_wr_req_desc_5_axaddr_1_addr;
   assign uc2rb_wr_req_desc_5_axaddr_2_reg[31:0] = int_wr_req_desc_5_axaddr_2_addr;
   assign uc2rb_wr_req_desc_5_axaddr_3_reg[31:0] = int_wr_req_desc_5_axaddr_3_addr;
   assign uc2rb_wr_req_desc_5_axid_0_reg[31:0] = int_wr_req_desc_5_axid_0_axid;
   assign uc2rb_wr_req_desc_5_axid_1_reg[31:0] = int_wr_req_desc_5_axid_1_axid;
   assign uc2rb_wr_req_desc_5_axid_2_reg[31:0] = int_wr_req_desc_5_axid_2_axid;
   assign uc2rb_wr_req_desc_5_axid_3_reg[31:0] = int_wr_req_desc_5_axid_3_axid;
   assign uc2rb_wr_req_desc_5_axuser_0_reg[31:0] = int_wr_req_desc_5_axuser_0_axuser;
   assign uc2rb_wr_req_desc_5_axuser_1_reg[31:0] = int_wr_req_desc_5_axuser_1_axuser;
   assign uc2rb_wr_req_desc_5_axuser_2_reg[31:0] = int_wr_req_desc_5_axuser_2_axuser;
   assign uc2rb_wr_req_desc_5_axuser_3_reg[31:0] = int_wr_req_desc_5_axuser_3_axuser;
   assign uc2rb_wr_req_desc_5_axuser_4_reg[31:0] = int_wr_req_desc_5_axuser_4_axuser;
   assign uc2rb_wr_req_desc_5_axuser_5_reg[31:0] = int_wr_req_desc_5_axuser_5_axuser;
   assign uc2rb_wr_req_desc_5_axuser_6_reg[31:0] = int_wr_req_desc_5_axuser_6_axuser;
   assign uc2rb_wr_req_desc_5_axuser_7_reg[31:0] = int_wr_req_desc_5_axuser_7_axuser;
   assign uc2rb_wr_req_desc_5_axuser_8_reg[31:0] = int_wr_req_desc_5_axuser_8_axuser;
   assign uc2rb_wr_req_desc_5_axuser_9_reg[31:0] = int_wr_req_desc_5_axuser_9_axuser;
   assign uc2rb_wr_req_desc_5_axuser_10_reg[31:0] = int_wr_req_desc_5_axuser_10_axuser;
   assign uc2rb_wr_req_desc_5_axuser_11_reg[31:0] = int_wr_req_desc_5_axuser_11_axuser;
   assign uc2rb_wr_req_desc_5_axuser_12_reg[31:0] = int_wr_req_desc_5_axuser_12_axuser;
   assign uc2rb_wr_req_desc_5_axuser_13_reg[31:0] = int_wr_req_desc_5_axuser_13_axuser;
   assign uc2rb_wr_req_desc_5_axuser_14_reg[31:0] = int_wr_req_desc_5_axuser_14_axuser;
   assign uc2rb_wr_req_desc_5_axuser_15_reg[31:0] = int_wr_req_desc_5_axuser_15_axuser;
   assign uc2rb_wr_req_desc_5_wuser_0_reg[31:0] = int_wr_req_desc_5_wuser_0_wuser;
   assign uc2rb_wr_req_desc_5_wuser_1_reg[31:0] = int_wr_req_desc_5_wuser_1_wuser;
   assign uc2rb_wr_req_desc_5_wuser_2_reg[31:0] = int_wr_req_desc_5_wuser_2_wuser;
   assign uc2rb_wr_req_desc_5_wuser_3_reg[31:0] = int_wr_req_desc_5_wuser_3_wuser;
   assign uc2rb_wr_req_desc_5_wuser_4_reg[31:0] = int_wr_req_desc_5_wuser_4_wuser;
   assign uc2rb_wr_req_desc_5_wuser_5_reg[31:0] = int_wr_req_desc_5_wuser_5_wuser;
   assign uc2rb_wr_req_desc_5_wuser_6_reg[31:0] = int_wr_req_desc_5_wuser_6_wuser;
   assign uc2rb_wr_req_desc_5_wuser_7_reg[31:0] = int_wr_req_desc_5_wuser_7_wuser;
   assign uc2rb_wr_req_desc_5_wuser_8_reg[31:0] = int_wr_req_desc_5_wuser_8_wuser;
   assign uc2rb_wr_req_desc_5_wuser_9_reg[31:0] = int_wr_req_desc_5_wuser_9_wuser;
   assign uc2rb_wr_req_desc_5_wuser_10_reg[31:0] = int_wr_req_desc_5_wuser_10_wuser;
   assign uc2rb_wr_req_desc_5_wuser_11_reg[31:0] = int_wr_req_desc_5_wuser_11_wuser;
   assign uc2rb_wr_req_desc_5_wuser_12_reg[31:0] = int_wr_req_desc_5_wuser_12_wuser;
   assign uc2rb_wr_req_desc_5_wuser_13_reg[31:0] = int_wr_req_desc_5_wuser_13_wuser;
   assign uc2rb_wr_req_desc_5_wuser_14_reg[31:0] = int_wr_req_desc_5_wuser_14_wuser;
   assign uc2rb_wr_req_desc_5_wuser_15_reg[31:0] = int_wr_req_desc_5_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_5_resp_reg[4:0] = int_sn_resp_desc_5_resp_resp;
   assign uc2rb_rd_req_desc_6_size_reg[31:0] = int_rd_req_desc_6_size_txn_size;
   assign uc2rb_rd_req_desc_6_axsize_reg[2:0] = int_rd_req_desc_6_axsize_axsize;
   assign uc2rb_rd_req_desc_6_attr_reg[27:24] = int_rd_req_desc_6_attr_axsnoop;
   assign uc2rb_rd_req_desc_6_attr_reg[23:22] = int_rd_req_desc_6_attr_axdomain;
   assign uc2rb_rd_req_desc_6_attr_reg[21:20] = int_rd_req_desc_6_attr_axbar;
   assign uc2rb_rd_req_desc_6_attr_reg[18:15] = int_rd_req_desc_6_attr_axregion;
   assign uc2rb_rd_req_desc_6_attr_reg[14:11] = int_rd_req_desc_6_attr_axqos;
   assign uc2rb_rd_req_desc_6_attr_reg[10:8] = int_rd_req_desc_6_attr_axprot;
   assign uc2rb_rd_req_desc_6_attr_reg[7:4] = int_rd_req_desc_6_attr_axcache;
   assign uc2rb_rd_req_desc_6_attr_reg[2] = int_rd_req_desc_6_attr_axlock;
   assign uc2rb_rd_req_desc_6_attr_reg[1:0] = int_rd_req_desc_6_attr_axburst;
   assign uc2rb_rd_req_desc_6_axaddr_0_reg[31:0] = int_rd_req_desc_6_axaddr_0_addr;
   assign uc2rb_rd_req_desc_6_axaddr_1_reg[31:0] = int_rd_req_desc_6_axaddr_1_addr;
   assign uc2rb_rd_req_desc_6_axaddr_2_reg[31:0] = int_rd_req_desc_6_axaddr_2_addr;
   assign uc2rb_rd_req_desc_6_axaddr_3_reg[31:0] = int_rd_req_desc_6_axaddr_3_addr;
   assign uc2rb_rd_req_desc_6_axid_0_reg[31:0] = int_rd_req_desc_6_axid_0_axid;
   assign uc2rb_rd_req_desc_6_axid_1_reg[31:0] = int_rd_req_desc_6_axid_1_axid;
   assign uc2rb_rd_req_desc_6_axid_2_reg[31:0] = int_rd_req_desc_6_axid_2_axid;
   assign uc2rb_rd_req_desc_6_axid_3_reg[31:0] = int_rd_req_desc_6_axid_3_axid;
   assign uc2rb_rd_req_desc_6_axuser_0_reg[31:0] = int_rd_req_desc_6_axuser_0_axuser;
   assign uc2rb_rd_req_desc_6_axuser_1_reg[31:0] = int_rd_req_desc_6_axuser_1_axuser;
   assign uc2rb_rd_req_desc_6_axuser_2_reg[31:0] = int_rd_req_desc_6_axuser_2_axuser;
   assign uc2rb_rd_req_desc_6_axuser_3_reg[31:0] = int_rd_req_desc_6_axuser_3_axuser;
   assign uc2rb_rd_req_desc_6_axuser_4_reg[31:0] = int_rd_req_desc_6_axuser_4_axuser;
   assign uc2rb_rd_req_desc_6_axuser_5_reg[31:0] = int_rd_req_desc_6_axuser_5_axuser;
   assign uc2rb_rd_req_desc_6_axuser_6_reg[31:0] = int_rd_req_desc_6_axuser_6_axuser;
   assign uc2rb_rd_req_desc_6_axuser_7_reg[31:0] = int_rd_req_desc_6_axuser_7_axuser;
   assign uc2rb_rd_req_desc_6_axuser_8_reg[31:0] = int_rd_req_desc_6_axuser_8_axuser;
   assign uc2rb_rd_req_desc_6_axuser_9_reg[31:0] = int_rd_req_desc_6_axuser_9_axuser;
   assign uc2rb_rd_req_desc_6_axuser_10_reg[31:0] = int_rd_req_desc_6_axuser_10_axuser;
   assign uc2rb_rd_req_desc_6_axuser_11_reg[31:0] = int_rd_req_desc_6_axuser_11_axuser;
   assign uc2rb_rd_req_desc_6_axuser_12_reg[31:0] = int_rd_req_desc_6_axuser_12_axuser;
   assign uc2rb_rd_req_desc_6_axuser_13_reg[31:0] = int_rd_req_desc_6_axuser_13_axuser;
   assign uc2rb_rd_req_desc_6_axuser_14_reg[31:0] = int_rd_req_desc_6_axuser_14_axuser;
   assign uc2rb_rd_req_desc_6_axuser_15_reg[31:0] = int_rd_req_desc_6_axuser_15_axuser;
   assign uc2rb_wr_req_desc_6_txn_type_reg[1] = int_wr_req_desc_6_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_6_size_reg[31:0] = int_wr_req_desc_6_size_txn_size;
   assign uc2rb_wr_req_desc_6_data_offset_reg[13:0] = int_wr_req_desc_6_data_offset_addr;
   assign uc2rb_wr_req_desc_6_axsize_reg[2:0] = int_wr_req_desc_6_axsize_axsize;
   assign uc2rb_wr_req_desc_6_attr_reg[27:24] = int_wr_req_desc_6_attr_axsnoop;
   assign uc2rb_wr_req_desc_6_attr_reg[23:22] = int_wr_req_desc_6_attr_axdomain;
   assign uc2rb_wr_req_desc_6_attr_reg[21:20] = int_wr_req_desc_6_attr_axbar;
   assign uc2rb_wr_req_desc_6_attr_reg[19] = int_wr_req_desc_6_attr_awunique;
   assign uc2rb_wr_req_desc_6_attr_reg[18:15] = int_wr_req_desc_6_attr_axregion;
   assign uc2rb_wr_req_desc_6_attr_reg[14:11] = int_wr_req_desc_6_attr_axqos;
   assign uc2rb_wr_req_desc_6_attr_reg[10:8] = int_wr_req_desc_6_attr_axprot;
   assign uc2rb_wr_req_desc_6_attr_reg[7:4] = int_wr_req_desc_6_attr_axcache;
   assign uc2rb_wr_req_desc_6_attr_reg[2] = int_wr_req_desc_6_attr_axlock;
   assign uc2rb_wr_req_desc_6_attr_reg[1:0] = int_wr_req_desc_6_attr_axburst;
   assign uc2rb_wr_req_desc_6_axaddr_0_reg[31:0] = int_wr_req_desc_6_axaddr_0_addr;
   assign uc2rb_wr_req_desc_6_axaddr_1_reg[31:0] = int_wr_req_desc_6_axaddr_1_addr;
   assign uc2rb_wr_req_desc_6_axaddr_2_reg[31:0] = int_wr_req_desc_6_axaddr_2_addr;
   assign uc2rb_wr_req_desc_6_axaddr_3_reg[31:0] = int_wr_req_desc_6_axaddr_3_addr;
   assign uc2rb_wr_req_desc_6_axid_0_reg[31:0] = int_wr_req_desc_6_axid_0_axid;
   assign uc2rb_wr_req_desc_6_axid_1_reg[31:0] = int_wr_req_desc_6_axid_1_axid;
   assign uc2rb_wr_req_desc_6_axid_2_reg[31:0] = int_wr_req_desc_6_axid_2_axid;
   assign uc2rb_wr_req_desc_6_axid_3_reg[31:0] = int_wr_req_desc_6_axid_3_axid;
   assign uc2rb_wr_req_desc_6_axuser_0_reg[31:0] = int_wr_req_desc_6_axuser_0_axuser;
   assign uc2rb_wr_req_desc_6_axuser_1_reg[31:0] = int_wr_req_desc_6_axuser_1_axuser;
   assign uc2rb_wr_req_desc_6_axuser_2_reg[31:0] = int_wr_req_desc_6_axuser_2_axuser;
   assign uc2rb_wr_req_desc_6_axuser_3_reg[31:0] = int_wr_req_desc_6_axuser_3_axuser;
   assign uc2rb_wr_req_desc_6_axuser_4_reg[31:0] = int_wr_req_desc_6_axuser_4_axuser;
   assign uc2rb_wr_req_desc_6_axuser_5_reg[31:0] = int_wr_req_desc_6_axuser_5_axuser;
   assign uc2rb_wr_req_desc_6_axuser_6_reg[31:0] = int_wr_req_desc_6_axuser_6_axuser;
   assign uc2rb_wr_req_desc_6_axuser_7_reg[31:0] = int_wr_req_desc_6_axuser_7_axuser;
   assign uc2rb_wr_req_desc_6_axuser_8_reg[31:0] = int_wr_req_desc_6_axuser_8_axuser;
   assign uc2rb_wr_req_desc_6_axuser_9_reg[31:0] = int_wr_req_desc_6_axuser_9_axuser;
   assign uc2rb_wr_req_desc_6_axuser_10_reg[31:0] = int_wr_req_desc_6_axuser_10_axuser;
   assign uc2rb_wr_req_desc_6_axuser_11_reg[31:0] = int_wr_req_desc_6_axuser_11_axuser;
   assign uc2rb_wr_req_desc_6_axuser_12_reg[31:0] = int_wr_req_desc_6_axuser_12_axuser;
   assign uc2rb_wr_req_desc_6_axuser_13_reg[31:0] = int_wr_req_desc_6_axuser_13_axuser;
   assign uc2rb_wr_req_desc_6_axuser_14_reg[31:0] = int_wr_req_desc_6_axuser_14_axuser;
   assign uc2rb_wr_req_desc_6_axuser_15_reg[31:0] = int_wr_req_desc_6_axuser_15_axuser;
   assign uc2rb_wr_req_desc_6_wuser_0_reg[31:0] = int_wr_req_desc_6_wuser_0_wuser;
   assign uc2rb_wr_req_desc_6_wuser_1_reg[31:0] = int_wr_req_desc_6_wuser_1_wuser;
   assign uc2rb_wr_req_desc_6_wuser_2_reg[31:0] = int_wr_req_desc_6_wuser_2_wuser;
   assign uc2rb_wr_req_desc_6_wuser_3_reg[31:0] = int_wr_req_desc_6_wuser_3_wuser;
   assign uc2rb_wr_req_desc_6_wuser_4_reg[31:0] = int_wr_req_desc_6_wuser_4_wuser;
   assign uc2rb_wr_req_desc_6_wuser_5_reg[31:0] = int_wr_req_desc_6_wuser_5_wuser;
   assign uc2rb_wr_req_desc_6_wuser_6_reg[31:0] = int_wr_req_desc_6_wuser_6_wuser;
   assign uc2rb_wr_req_desc_6_wuser_7_reg[31:0] = int_wr_req_desc_6_wuser_7_wuser;
   assign uc2rb_wr_req_desc_6_wuser_8_reg[31:0] = int_wr_req_desc_6_wuser_8_wuser;
   assign uc2rb_wr_req_desc_6_wuser_9_reg[31:0] = int_wr_req_desc_6_wuser_9_wuser;
   assign uc2rb_wr_req_desc_6_wuser_10_reg[31:0] = int_wr_req_desc_6_wuser_10_wuser;
   assign uc2rb_wr_req_desc_6_wuser_11_reg[31:0] = int_wr_req_desc_6_wuser_11_wuser;
   assign uc2rb_wr_req_desc_6_wuser_12_reg[31:0] = int_wr_req_desc_6_wuser_12_wuser;
   assign uc2rb_wr_req_desc_6_wuser_13_reg[31:0] = int_wr_req_desc_6_wuser_13_wuser;
   assign uc2rb_wr_req_desc_6_wuser_14_reg[31:0] = int_wr_req_desc_6_wuser_14_wuser;
   assign uc2rb_wr_req_desc_6_wuser_15_reg[31:0] = int_wr_req_desc_6_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_6_resp_reg[4:0] = int_sn_resp_desc_6_resp_resp;
   assign uc2rb_rd_req_desc_7_size_reg[31:0] = int_rd_req_desc_7_size_txn_size;
   assign uc2rb_rd_req_desc_7_axsize_reg[2:0] = int_rd_req_desc_7_axsize_axsize;
   assign uc2rb_rd_req_desc_7_attr_reg[27:24] = int_rd_req_desc_7_attr_axsnoop;
   assign uc2rb_rd_req_desc_7_attr_reg[23:22] = int_rd_req_desc_7_attr_axdomain;
   assign uc2rb_rd_req_desc_7_attr_reg[21:20] = int_rd_req_desc_7_attr_axbar;
   assign uc2rb_rd_req_desc_7_attr_reg[18:15] = int_rd_req_desc_7_attr_axregion;
   assign uc2rb_rd_req_desc_7_attr_reg[14:11] = int_rd_req_desc_7_attr_axqos;
   assign uc2rb_rd_req_desc_7_attr_reg[10:8] = int_rd_req_desc_7_attr_axprot;
   assign uc2rb_rd_req_desc_7_attr_reg[7:4] = int_rd_req_desc_7_attr_axcache;
   assign uc2rb_rd_req_desc_7_attr_reg[2] = int_rd_req_desc_7_attr_axlock;
   assign uc2rb_rd_req_desc_7_attr_reg[1:0] = int_rd_req_desc_7_attr_axburst;
   assign uc2rb_rd_req_desc_7_axaddr_0_reg[31:0] = int_rd_req_desc_7_axaddr_0_addr;
   assign uc2rb_rd_req_desc_7_axaddr_1_reg[31:0] = int_rd_req_desc_7_axaddr_1_addr;
   assign uc2rb_rd_req_desc_7_axaddr_2_reg[31:0] = int_rd_req_desc_7_axaddr_2_addr;
   assign uc2rb_rd_req_desc_7_axaddr_3_reg[31:0] = int_rd_req_desc_7_axaddr_3_addr;
   assign uc2rb_rd_req_desc_7_axid_0_reg[31:0] = int_rd_req_desc_7_axid_0_axid;
   assign uc2rb_rd_req_desc_7_axid_1_reg[31:0] = int_rd_req_desc_7_axid_1_axid;
   assign uc2rb_rd_req_desc_7_axid_2_reg[31:0] = int_rd_req_desc_7_axid_2_axid;
   assign uc2rb_rd_req_desc_7_axid_3_reg[31:0] = int_rd_req_desc_7_axid_3_axid;
   assign uc2rb_rd_req_desc_7_axuser_0_reg[31:0] = int_rd_req_desc_7_axuser_0_axuser;
   assign uc2rb_rd_req_desc_7_axuser_1_reg[31:0] = int_rd_req_desc_7_axuser_1_axuser;
   assign uc2rb_rd_req_desc_7_axuser_2_reg[31:0] = int_rd_req_desc_7_axuser_2_axuser;
   assign uc2rb_rd_req_desc_7_axuser_3_reg[31:0] = int_rd_req_desc_7_axuser_3_axuser;
   assign uc2rb_rd_req_desc_7_axuser_4_reg[31:0] = int_rd_req_desc_7_axuser_4_axuser;
   assign uc2rb_rd_req_desc_7_axuser_5_reg[31:0] = int_rd_req_desc_7_axuser_5_axuser;
   assign uc2rb_rd_req_desc_7_axuser_6_reg[31:0] = int_rd_req_desc_7_axuser_6_axuser;
   assign uc2rb_rd_req_desc_7_axuser_7_reg[31:0] = int_rd_req_desc_7_axuser_7_axuser;
   assign uc2rb_rd_req_desc_7_axuser_8_reg[31:0] = int_rd_req_desc_7_axuser_8_axuser;
   assign uc2rb_rd_req_desc_7_axuser_9_reg[31:0] = int_rd_req_desc_7_axuser_9_axuser;
   assign uc2rb_rd_req_desc_7_axuser_10_reg[31:0] = int_rd_req_desc_7_axuser_10_axuser;
   assign uc2rb_rd_req_desc_7_axuser_11_reg[31:0] = int_rd_req_desc_7_axuser_11_axuser;
   assign uc2rb_rd_req_desc_7_axuser_12_reg[31:0] = int_rd_req_desc_7_axuser_12_axuser;
   assign uc2rb_rd_req_desc_7_axuser_13_reg[31:0] = int_rd_req_desc_7_axuser_13_axuser;
   assign uc2rb_rd_req_desc_7_axuser_14_reg[31:0] = int_rd_req_desc_7_axuser_14_axuser;
   assign uc2rb_rd_req_desc_7_axuser_15_reg[31:0] = int_rd_req_desc_7_axuser_15_axuser;
   assign uc2rb_wr_req_desc_7_txn_type_reg[1] = int_wr_req_desc_7_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_7_size_reg[31:0] = int_wr_req_desc_7_size_txn_size;
   assign uc2rb_wr_req_desc_7_data_offset_reg[13:0] = int_wr_req_desc_7_data_offset_addr;
   assign uc2rb_wr_req_desc_7_axsize_reg[2:0] = int_wr_req_desc_7_axsize_axsize;
   assign uc2rb_wr_req_desc_7_attr_reg[27:24] = int_wr_req_desc_7_attr_axsnoop;
   assign uc2rb_wr_req_desc_7_attr_reg[23:22] = int_wr_req_desc_7_attr_axdomain;
   assign uc2rb_wr_req_desc_7_attr_reg[21:20] = int_wr_req_desc_7_attr_axbar;
   assign uc2rb_wr_req_desc_7_attr_reg[19] = int_wr_req_desc_7_attr_awunique;
   assign uc2rb_wr_req_desc_7_attr_reg[18:15] = int_wr_req_desc_7_attr_axregion;
   assign uc2rb_wr_req_desc_7_attr_reg[14:11] = int_wr_req_desc_7_attr_axqos;
   assign uc2rb_wr_req_desc_7_attr_reg[10:8] = int_wr_req_desc_7_attr_axprot;
   assign uc2rb_wr_req_desc_7_attr_reg[7:4] = int_wr_req_desc_7_attr_axcache;
   assign uc2rb_wr_req_desc_7_attr_reg[2] = int_wr_req_desc_7_attr_axlock;
   assign uc2rb_wr_req_desc_7_attr_reg[1:0] = int_wr_req_desc_7_attr_axburst;
   assign uc2rb_wr_req_desc_7_axaddr_0_reg[31:0] = int_wr_req_desc_7_axaddr_0_addr;
   assign uc2rb_wr_req_desc_7_axaddr_1_reg[31:0] = int_wr_req_desc_7_axaddr_1_addr;
   assign uc2rb_wr_req_desc_7_axaddr_2_reg[31:0] = int_wr_req_desc_7_axaddr_2_addr;
   assign uc2rb_wr_req_desc_7_axaddr_3_reg[31:0] = int_wr_req_desc_7_axaddr_3_addr;
   assign uc2rb_wr_req_desc_7_axid_0_reg[31:0] = int_wr_req_desc_7_axid_0_axid;
   assign uc2rb_wr_req_desc_7_axid_1_reg[31:0] = int_wr_req_desc_7_axid_1_axid;
   assign uc2rb_wr_req_desc_7_axid_2_reg[31:0] = int_wr_req_desc_7_axid_2_axid;
   assign uc2rb_wr_req_desc_7_axid_3_reg[31:0] = int_wr_req_desc_7_axid_3_axid;
   assign uc2rb_wr_req_desc_7_axuser_0_reg[31:0] = int_wr_req_desc_7_axuser_0_axuser;
   assign uc2rb_wr_req_desc_7_axuser_1_reg[31:0] = int_wr_req_desc_7_axuser_1_axuser;
   assign uc2rb_wr_req_desc_7_axuser_2_reg[31:0] = int_wr_req_desc_7_axuser_2_axuser;
   assign uc2rb_wr_req_desc_7_axuser_3_reg[31:0] = int_wr_req_desc_7_axuser_3_axuser;
   assign uc2rb_wr_req_desc_7_axuser_4_reg[31:0] = int_wr_req_desc_7_axuser_4_axuser;
   assign uc2rb_wr_req_desc_7_axuser_5_reg[31:0] = int_wr_req_desc_7_axuser_5_axuser;
   assign uc2rb_wr_req_desc_7_axuser_6_reg[31:0] = int_wr_req_desc_7_axuser_6_axuser;
   assign uc2rb_wr_req_desc_7_axuser_7_reg[31:0] = int_wr_req_desc_7_axuser_7_axuser;
   assign uc2rb_wr_req_desc_7_axuser_8_reg[31:0] = int_wr_req_desc_7_axuser_8_axuser;
   assign uc2rb_wr_req_desc_7_axuser_9_reg[31:0] = int_wr_req_desc_7_axuser_9_axuser;
   assign uc2rb_wr_req_desc_7_axuser_10_reg[31:0] = int_wr_req_desc_7_axuser_10_axuser;
   assign uc2rb_wr_req_desc_7_axuser_11_reg[31:0] = int_wr_req_desc_7_axuser_11_axuser;
   assign uc2rb_wr_req_desc_7_axuser_12_reg[31:0] = int_wr_req_desc_7_axuser_12_axuser;
   assign uc2rb_wr_req_desc_7_axuser_13_reg[31:0] = int_wr_req_desc_7_axuser_13_axuser;
   assign uc2rb_wr_req_desc_7_axuser_14_reg[31:0] = int_wr_req_desc_7_axuser_14_axuser;
   assign uc2rb_wr_req_desc_7_axuser_15_reg[31:0] = int_wr_req_desc_7_axuser_15_axuser;
   assign uc2rb_wr_req_desc_7_wuser_0_reg[31:0] = int_wr_req_desc_7_wuser_0_wuser;
   assign uc2rb_wr_req_desc_7_wuser_1_reg[31:0] = int_wr_req_desc_7_wuser_1_wuser;
   assign uc2rb_wr_req_desc_7_wuser_2_reg[31:0] = int_wr_req_desc_7_wuser_2_wuser;
   assign uc2rb_wr_req_desc_7_wuser_3_reg[31:0] = int_wr_req_desc_7_wuser_3_wuser;
   assign uc2rb_wr_req_desc_7_wuser_4_reg[31:0] = int_wr_req_desc_7_wuser_4_wuser;
   assign uc2rb_wr_req_desc_7_wuser_5_reg[31:0] = int_wr_req_desc_7_wuser_5_wuser;
   assign uc2rb_wr_req_desc_7_wuser_6_reg[31:0] = int_wr_req_desc_7_wuser_6_wuser;
   assign uc2rb_wr_req_desc_7_wuser_7_reg[31:0] = int_wr_req_desc_7_wuser_7_wuser;
   assign uc2rb_wr_req_desc_7_wuser_8_reg[31:0] = int_wr_req_desc_7_wuser_8_wuser;
   assign uc2rb_wr_req_desc_7_wuser_9_reg[31:0] = int_wr_req_desc_7_wuser_9_wuser;
   assign uc2rb_wr_req_desc_7_wuser_10_reg[31:0] = int_wr_req_desc_7_wuser_10_wuser;
   assign uc2rb_wr_req_desc_7_wuser_11_reg[31:0] = int_wr_req_desc_7_wuser_11_wuser;
   assign uc2rb_wr_req_desc_7_wuser_12_reg[31:0] = int_wr_req_desc_7_wuser_12_wuser;
   assign uc2rb_wr_req_desc_7_wuser_13_reg[31:0] = int_wr_req_desc_7_wuser_13_wuser;
   assign uc2rb_wr_req_desc_7_wuser_14_reg[31:0] = int_wr_req_desc_7_wuser_14_wuser;
   assign uc2rb_wr_req_desc_7_wuser_15_reg[31:0] = int_wr_req_desc_7_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_7_resp_reg[4:0] = int_sn_resp_desc_7_resp_resp;
   assign uc2rb_rd_req_desc_8_size_reg[31:0] = int_rd_req_desc_8_size_txn_size;
   assign uc2rb_rd_req_desc_8_axsize_reg[2:0] = int_rd_req_desc_8_axsize_axsize;
   assign uc2rb_rd_req_desc_8_attr_reg[27:24] = int_rd_req_desc_8_attr_axsnoop;
   assign uc2rb_rd_req_desc_8_attr_reg[23:22] = int_rd_req_desc_8_attr_axdomain;
   assign uc2rb_rd_req_desc_8_attr_reg[21:20] = int_rd_req_desc_8_attr_axbar;
   assign uc2rb_rd_req_desc_8_attr_reg[18:15] = int_rd_req_desc_8_attr_axregion;
   assign uc2rb_rd_req_desc_8_attr_reg[14:11] = int_rd_req_desc_8_attr_axqos;
   assign uc2rb_rd_req_desc_8_attr_reg[10:8] = int_rd_req_desc_8_attr_axprot;
   assign uc2rb_rd_req_desc_8_attr_reg[7:4] = int_rd_req_desc_8_attr_axcache;
   assign uc2rb_rd_req_desc_8_attr_reg[2] = int_rd_req_desc_8_attr_axlock;
   assign uc2rb_rd_req_desc_8_attr_reg[1:0] = int_rd_req_desc_8_attr_axburst;
   assign uc2rb_rd_req_desc_8_axaddr_0_reg[31:0] = int_rd_req_desc_8_axaddr_0_addr;
   assign uc2rb_rd_req_desc_8_axaddr_1_reg[31:0] = int_rd_req_desc_8_axaddr_1_addr;
   assign uc2rb_rd_req_desc_8_axaddr_2_reg[31:0] = int_rd_req_desc_8_axaddr_2_addr;
   assign uc2rb_rd_req_desc_8_axaddr_3_reg[31:0] = int_rd_req_desc_8_axaddr_3_addr;
   assign uc2rb_rd_req_desc_8_axid_0_reg[31:0] = int_rd_req_desc_8_axid_0_axid;
   assign uc2rb_rd_req_desc_8_axid_1_reg[31:0] = int_rd_req_desc_8_axid_1_axid;
   assign uc2rb_rd_req_desc_8_axid_2_reg[31:0] = int_rd_req_desc_8_axid_2_axid;
   assign uc2rb_rd_req_desc_8_axid_3_reg[31:0] = int_rd_req_desc_8_axid_3_axid;
   assign uc2rb_rd_req_desc_8_axuser_0_reg[31:0] = int_rd_req_desc_8_axuser_0_axuser;
   assign uc2rb_rd_req_desc_8_axuser_1_reg[31:0] = int_rd_req_desc_8_axuser_1_axuser;
   assign uc2rb_rd_req_desc_8_axuser_2_reg[31:0] = int_rd_req_desc_8_axuser_2_axuser;
   assign uc2rb_rd_req_desc_8_axuser_3_reg[31:0] = int_rd_req_desc_8_axuser_3_axuser;
   assign uc2rb_rd_req_desc_8_axuser_4_reg[31:0] = int_rd_req_desc_8_axuser_4_axuser;
   assign uc2rb_rd_req_desc_8_axuser_5_reg[31:0] = int_rd_req_desc_8_axuser_5_axuser;
   assign uc2rb_rd_req_desc_8_axuser_6_reg[31:0] = int_rd_req_desc_8_axuser_6_axuser;
   assign uc2rb_rd_req_desc_8_axuser_7_reg[31:0] = int_rd_req_desc_8_axuser_7_axuser;
   assign uc2rb_rd_req_desc_8_axuser_8_reg[31:0] = int_rd_req_desc_8_axuser_8_axuser;
   assign uc2rb_rd_req_desc_8_axuser_9_reg[31:0] = int_rd_req_desc_8_axuser_9_axuser;
   assign uc2rb_rd_req_desc_8_axuser_10_reg[31:0] = int_rd_req_desc_8_axuser_10_axuser;
   assign uc2rb_rd_req_desc_8_axuser_11_reg[31:0] = int_rd_req_desc_8_axuser_11_axuser;
   assign uc2rb_rd_req_desc_8_axuser_12_reg[31:0] = int_rd_req_desc_8_axuser_12_axuser;
   assign uc2rb_rd_req_desc_8_axuser_13_reg[31:0] = int_rd_req_desc_8_axuser_13_axuser;
   assign uc2rb_rd_req_desc_8_axuser_14_reg[31:0] = int_rd_req_desc_8_axuser_14_axuser;
   assign uc2rb_rd_req_desc_8_axuser_15_reg[31:0] = int_rd_req_desc_8_axuser_15_axuser;
   assign uc2rb_wr_req_desc_8_txn_type_reg[1] = int_wr_req_desc_8_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_8_size_reg[31:0] = int_wr_req_desc_8_size_txn_size;
   assign uc2rb_wr_req_desc_8_data_offset_reg[13:0] = int_wr_req_desc_8_data_offset_addr;
   assign uc2rb_wr_req_desc_8_axsize_reg[2:0] = int_wr_req_desc_8_axsize_axsize;
   assign uc2rb_wr_req_desc_8_attr_reg[27:24] = int_wr_req_desc_8_attr_axsnoop;
   assign uc2rb_wr_req_desc_8_attr_reg[23:22] = int_wr_req_desc_8_attr_axdomain;
   assign uc2rb_wr_req_desc_8_attr_reg[21:20] = int_wr_req_desc_8_attr_axbar;
   assign uc2rb_wr_req_desc_8_attr_reg[19] = int_wr_req_desc_8_attr_awunique;
   assign uc2rb_wr_req_desc_8_attr_reg[18:15] = int_wr_req_desc_8_attr_axregion;
   assign uc2rb_wr_req_desc_8_attr_reg[14:11] = int_wr_req_desc_8_attr_axqos;
   assign uc2rb_wr_req_desc_8_attr_reg[10:8] = int_wr_req_desc_8_attr_axprot;
   assign uc2rb_wr_req_desc_8_attr_reg[7:4] = int_wr_req_desc_8_attr_axcache;
   assign uc2rb_wr_req_desc_8_attr_reg[2] = int_wr_req_desc_8_attr_axlock;
   assign uc2rb_wr_req_desc_8_attr_reg[1:0] = int_wr_req_desc_8_attr_axburst;
   assign uc2rb_wr_req_desc_8_axaddr_0_reg[31:0] = int_wr_req_desc_8_axaddr_0_addr;
   assign uc2rb_wr_req_desc_8_axaddr_1_reg[31:0] = int_wr_req_desc_8_axaddr_1_addr;
   assign uc2rb_wr_req_desc_8_axaddr_2_reg[31:0] = int_wr_req_desc_8_axaddr_2_addr;
   assign uc2rb_wr_req_desc_8_axaddr_3_reg[31:0] = int_wr_req_desc_8_axaddr_3_addr;
   assign uc2rb_wr_req_desc_8_axid_0_reg[31:0] = int_wr_req_desc_8_axid_0_axid;
   assign uc2rb_wr_req_desc_8_axid_1_reg[31:0] = int_wr_req_desc_8_axid_1_axid;
   assign uc2rb_wr_req_desc_8_axid_2_reg[31:0] = int_wr_req_desc_8_axid_2_axid;
   assign uc2rb_wr_req_desc_8_axid_3_reg[31:0] = int_wr_req_desc_8_axid_3_axid;
   assign uc2rb_wr_req_desc_8_axuser_0_reg[31:0] = int_wr_req_desc_8_axuser_0_axuser;
   assign uc2rb_wr_req_desc_8_axuser_1_reg[31:0] = int_wr_req_desc_8_axuser_1_axuser;
   assign uc2rb_wr_req_desc_8_axuser_2_reg[31:0] = int_wr_req_desc_8_axuser_2_axuser;
   assign uc2rb_wr_req_desc_8_axuser_3_reg[31:0] = int_wr_req_desc_8_axuser_3_axuser;
   assign uc2rb_wr_req_desc_8_axuser_4_reg[31:0] = int_wr_req_desc_8_axuser_4_axuser;
   assign uc2rb_wr_req_desc_8_axuser_5_reg[31:0] = int_wr_req_desc_8_axuser_5_axuser;
   assign uc2rb_wr_req_desc_8_axuser_6_reg[31:0] = int_wr_req_desc_8_axuser_6_axuser;
   assign uc2rb_wr_req_desc_8_axuser_7_reg[31:0] = int_wr_req_desc_8_axuser_7_axuser;
   assign uc2rb_wr_req_desc_8_axuser_8_reg[31:0] = int_wr_req_desc_8_axuser_8_axuser;
   assign uc2rb_wr_req_desc_8_axuser_9_reg[31:0] = int_wr_req_desc_8_axuser_9_axuser;
   assign uc2rb_wr_req_desc_8_axuser_10_reg[31:0] = int_wr_req_desc_8_axuser_10_axuser;
   assign uc2rb_wr_req_desc_8_axuser_11_reg[31:0] = int_wr_req_desc_8_axuser_11_axuser;
   assign uc2rb_wr_req_desc_8_axuser_12_reg[31:0] = int_wr_req_desc_8_axuser_12_axuser;
   assign uc2rb_wr_req_desc_8_axuser_13_reg[31:0] = int_wr_req_desc_8_axuser_13_axuser;
   assign uc2rb_wr_req_desc_8_axuser_14_reg[31:0] = int_wr_req_desc_8_axuser_14_axuser;
   assign uc2rb_wr_req_desc_8_axuser_15_reg[31:0] = int_wr_req_desc_8_axuser_15_axuser;
   assign uc2rb_wr_req_desc_8_wuser_0_reg[31:0] = int_wr_req_desc_8_wuser_0_wuser;
   assign uc2rb_wr_req_desc_8_wuser_1_reg[31:0] = int_wr_req_desc_8_wuser_1_wuser;
   assign uc2rb_wr_req_desc_8_wuser_2_reg[31:0] = int_wr_req_desc_8_wuser_2_wuser;
   assign uc2rb_wr_req_desc_8_wuser_3_reg[31:0] = int_wr_req_desc_8_wuser_3_wuser;
   assign uc2rb_wr_req_desc_8_wuser_4_reg[31:0] = int_wr_req_desc_8_wuser_4_wuser;
   assign uc2rb_wr_req_desc_8_wuser_5_reg[31:0] = int_wr_req_desc_8_wuser_5_wuser;
   assign uc2rb_wr_req_desc_8_wuser_6_reg[31:0] = int_wr_req_desc_8_wuser_6_wuser;
   assign uc2rb_wr_req_desc_8_wuser_7_reg[31:0] = int_wr_req_desc_8_wuser_7_wuser;
   assign uc2rb_wr_req_desc_8_wuser_8_reg[31:0] = int_wr_req_desc_8_wuser_8_wuser;
   assign uc2rb_wr_req_desc_8_wuser_9_reg[31:0] = int_wr_req_desc_8_wuser_9_wuser;
   assign uc2rb_wr_req_desc_8_wuser_10_reg[31:0] = int_wr_req_desc_8_wuser_10_wuser;
   assign uc2rb_wr_req_desc_8_wuser_11_reg[31:0] = int_wr_req_desc_8_wuser_11_wuser;
   assign uc2rb_wr_req_desc_8_wuser_12_reg[31:0] = int_wr_req_desc_8_wuser_12_wuser;
   assign uc2rb_wr_req_desc_8_wuser_13_reg[31:0] = int_wr_req_desc_8_wuser_13_wuser;
   assign uc2rb_wr_req_desc_8_wuser_14_reg[31:0] = int_wr_req_desc_8_wuser_14_wuser;
   assign uc2rb_wr_req_desc_8_wuser_15_reg[31:0] = int_wr_req_desc_8_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_8_resp_reg[4:0] = int_sn_resp_desc_8_resp_resp;
   assign uc2rb_rd_req_desc_9_size_reg[31:0] = int_rd_req_desc_9_size_txn_size;
   assign uc2rb_rd_req_desc_9_axsize_reg[2:0] = int_rd_req_desc_9_axsize_axsize;
   assign uc2rb_rd_req_desc_9_attr_reg[27:24] = int_rd_req_desc_9_attr_axsnoop;
   assign uc2rb_rd_req_desc_9_attr_reg[23:22] = int_rd_req_desc_9_attr_axdomain;
   assign uc2rb_rd_req_desc_9_attr_reg[21:20] = int_rd_req_desc_9_attr_axbar;
   assign uc2rb_rd_req_desc_9_attr_reg[18:15] = int_rd_req_desc_9_attr_axregion;
   assign uc2rb_rd_req_desc_9_attr_reg[14:11] = int_rd_req_desc_9_attr_axqos;
   assign uc2rb_rd_req_desc_9_attr_reg[10:8] = int_rd_req_desc_9_attr_axprot;
   assign uc2rb_rd_req_desc_9_attr_reg[7:4] = int_rd_req_desc_9_attr_axcache;
   assign uc2rb_rd_req_desc_9_attr_reg[2] = int_rd_req_desc_9_attr_axlock;
   assign uc2rb_rd_req_desc_9_attr_reg[1:0] = int_rd_req_desc_9_attr_axburst;
   assign uc2rb_rd_req_desc_9_axaddr_0_reg[31:0] = int_rd_req_desc_9_axaddr_0_addr;
   assign uc2rb_rd_req_desc_9_axaddr_1_reg[31:0] = int_rd_req_desc_9_axaddr_1_addr;
   assign uc2rb_rd_req_desc_9_axaddr_2_reg[31:0] = int_rd_req_desc_9_axaddr_2_addr;
   assign uc2rb_rd_req_desc_9_axaddr_3_reg[31:0] = int_rd_req_desc_9_axaddr_3_addr;
   assign uc2rb_rd_req_desc_9_axid_0_reg[31:0] = int_rd_req_desc_9_axid_0_axid;
   assign uc2rb_rd_req_desc_9_axid_1_reg[31:0] = int_rd_req_desc_9_axid_1_axid;
   assign uc2rb_rd_req_desc_9_axid_2_reg[31:0] = int_rd_req_desc_9_axid_2_axid;
   assign uc2rb_rd_req_desc_9_axid_3_reg[31:0] = int_rd_req_desc_9_axid_3_axid;
   assign uc2rb_rd_req_desc_9_axuser_0_reg[31:0] = int_rd_req_desc_9_axuser_0_axuser;
   assign uc2rb_rd_req_desc_9_axuser_1_reg[31:0] = int_rd_req_desc_9_axuser_1_axuser;
   assign uc2rb_rd_req_desc_9_axuser_2_reg[31:0] = int_rd_req_desc_9_axuser_2_axuser;
   assign uc2rb_rd_req_desc_9_axuser_3_reg[31:0] = int_rd_req_desc_9_axuser_3_axuser;
   assign uc2rb_rd_req_desc_9_axuser_4_reg[31:0] = int_rd_req_desc_9_axuser_4_axuser;
   assign uc2rb_rd_req_desc_9_axuser_5_reg[31:0] = int_rd_req_desc_9_axuser_5_axuser;
   assign uc2rb_rd_req_desc_9_axuser_6_reg[31:0] = int_rd_req_desc_9_axuser_6_axuser;
   assign uc2rb_rd_req_desc_9_axuser_7_reg[31:0] = int_rd_req_desc_9_axuser_7_axuser;
   assign uc2rb_rd_req_desc_9_axuser_8_reg[31:0] = int_rd_req_desc_9_axuser_8_axuser;
   assign uc2rb_rd_req_desc_9_axuser_9_reg[31:0] = int_rd_req_desc_9_axuser_9_axuser;
   assign uc2rb_rd_req_desc_9_axuser_10_reg[31:0] = int_rd_req_desc_9_axuser_10_axuser;
   assign uc2rb_rd_req_desc_9_axuser_11_reg[31:0] = int_rd_req_desc_9_axuser_11_axuser;
   assign uc2rb_rd_req_desc_9_axuser_12_reg[31:0] = int_rd_req_desc_9_axuser_12_axuser;
   assign uc2rb_rd_req_desc_9_axuser_13_reg[31:0] = int_rd_req_desc_9_axuser_13_axuser;
   assign uc2rb_rd_req_desc_9_axuser_14_reg[31:0] = int_rd_req_desc_9_axuser_14_axuser;
   assign uc2rb_rd_req_desc_9_axuser_15_reg[31:0] = int_rd_req_desc_9_axuser_15_axuser;
   assign uc2rb_wr_req_desc_9_txn_type_reg[1] = int_wr_req_desc_9_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_9_size_reg[31:0] = int_wr_req_desc_9_size_txn_size;
   assign uc2rb_wr_req_desc_9_data_offset_reg[13:0] = int_wr_req_desc_9_data_offset_addr;
   assign uc2rb_wr_req_desc_9_axsize_reg[2:0] = int_wr_req_desc_9_axsize_axsize;
   assign uc2rb_wr_req_desc_9_attr_reg[27:24] = int_wr_req_desc_9_attr_axsnoop;
   assign uc2rb_wr_req_desc_9_attr_reg[23:22] = int_wr_req_desc_9_attr_axdomain;
   assign uc2rb_wr_req_desc_9_attr_reg[21:20] = int_wr_req_desc_9_attr_axbar;
   assign uc2rb_wr_req_desc_9_attr_reg[19] = int_wr_req_desc_9_attr_awunique;
   assign uc2rb_wr_req_desc_9_attr_reg[18:15] = int_wr_req_desc_9_attr_axregion;
   assign uc2rb_wr_req_desc_9_attr_reg[14:11] = int_wr_req_desc_9_attr_axqos;
   assign uc2rb_wr_req_desc_9_attr_reg[10:8] = int_wr_req_desc_9_attr_axprot;
   assign uc2rb_wr_req_desc_9_attr_reg[7:4] = int_wr_req_desc_9_attr_axcache;
   assign uc2rb_wr_req_desc_9_attr_reg[2] = int_wr_req_desc_9_attr_axlock;
   assign uc2rb_wr_req_desc_9_attr_reg[1:0] = int_wr_req_desc_9_attr_axburst;
   assign uc2rb_wr_req_desc_9_axaddr_0_reg[31:0] = int_wr_req_desc_9_axaddr_0_addr;
   assign uc2rb_wr_req_desc_9_axaddr_1_reg[31:0] = int_wr_req_desc_9_axaddr_1_addr;
   assign uc2rb_wr_req_desc_9_axaddr_2_reg[31:0] = int_wr_req_desc_9_axaddr_2_addr;
   assign uc2rb_wr_req_desc_9_axaddr_3_reg[31:0] = int_wr_req_desc_9_axaddr_3_addr;
   assign uc2rb_wr_req_desc_9_axid_0_reg[31:0] = int_wr_req_desc_9_axid_0_axid;
   assign uc2rb_wr_req_desc_9_axid_1_reg[31:0] = int_wr_req_desc_9_axid_1_axid;
   assign uc2rb_wr_req_desc_9_axid_2_reg[31:0] = int_wr_req_desc_9_axid_2_axid;
   assign uc2rb_wr_req_desc_9_axid_3_reg[31:0] = int_wr_req_desc_9_axid_3_axid;
   assign uc2rb_wr_req_desc_9_axuser_0_reg[31:0] = int_wr_req_desc_9_axuser_0_axuser;
   assign uc2rb_wr_req_desc_9_axuser_1_reg[31:0] = int_wr_req_desc_9_axuser_1_axuser;
   assign uc2rb_wr_req_desc_9_axuser_2_reg[31:0] = int_wr_req_desc_9_axuser_2_axuser;
   assign uc2rb_wr_req_desc_9_axuser_3_reg[31:0] = int_wr_req_desc_9_axuser_3_axuser;
   assign uc2rb_wr_req_desc_9_axuser_4_reg[31:0] = int_wr_req_desc_9_axuser_4_axuser;
   assign uc2rb_wr_req_desc_9_axuser_5_reg[31:0] = int_wr_req_desc_9_axuser_5_axuser;
   assign uc2rb_wr_req_desc_9_axuser_6_reg[31:0] = int_wr_req_desc_9_axuser_6_axuser;
   assign uc2rb_wr_req_desc_9_axuser_7_reg[31:0] = int_wr_req_desc_9_axuser_7_axuser;
   assign uc2rb_wr_req_desc_9_axuser_8_reg[31:0] = int_wr_req_desc_9_axuser_8_axuser;
   assign uc2rb_wr_req_desc_9_axuser_9_reg[31:0] = int_wr_req_desc_9_axuser_9_axuser;
   assign uc2rb_wr_req_desc_9_axuser_10_reg[31:0] = int_wr_req_desc_9_axuser_10_axuser;
   assign uc2rb_wr_req_desc_9_axuser_11_reg[31:0] = int_wr_req_desc_9_axuser_11_axuser;
   assign uc2rb_wr_req_desc_9_axuser_12_reg[31:0] = int_wr_req_desc_9_axuser_12_axuser;
   assign uc2rb_wr_req_desc_9_axuser_13_reg[31:0] = int_wr_req_desc_9_axuser_13_axuser;
   assign uc2rb_wr_req_desc_9_axuser_14_reg[31:0] = int_wr_req_desc_9_axuser_14_axuser;
   assign uc2rb_wr_req_desc_9_axuser_15_reg[31:0] = int_wr_req_desc_9_axuser_15_axuser;
   assign uc2rb_wr_req_desc_9_wuser_0_reg[31:0] = int_wr_req_desc_9_wuser_0_wuser;
   assign uc2rb_wr_req_desc_9_wuser_1_reg[31:0] = int_wr_req_desc_9_wuser_1_wuser;
   assign uc2rb_wr_req_desc_9_wuser_2_reg[31:0] = int_wr_req_desc_9_wuser_2_wuser;
   assign uc2rb_wr_req_desc_9_wuser_3_reg[31:0] = int_wr_req_desc_9_wuser_3_wuser;
   assign uc2rb_wr_req_desc_9_wuser_4_reg[31:0] = int_wr_req_desc_9_wuser_4_wuser;
   assign uc2rb_wr_req_desc_9_wuser_5_reg[31:0] = int_wr_req_desc_9_wuser_5_wuser;
   assign uc2rb_wr_req_desc_9_wuser_6_reg[31:0] = int_wr_req_desc_9_wuser_6_wuser;
   assign uc2rb_wr_req_desc_9_wuser_7_reg[31:0] = int_wr_req_desc_9_wuser_7_wuser;
   assign uc2rb_wr_req_desc_9_wuser_8_reg[31:0] = int_wr_req_desc_9_wuser_8_wuser;
   assign uc2rb_wr_req_desc_9_wuser_9_reg[31:0] = int_wr_req_desc_9_wuser_9_wuser;
   assign uc2rb_wr_req_desc_9_wuser_10_reg[31:0] = int_wr_req_desc_9_wuser_10_wuser;
   assign uc2rb_wr_req_desc_9_wuser_11_reg[31:0] = int_wr_req_desc_9_wuser_11_wuser;
   assign uc2rb_wr_req_desc_9_wuser_12_reg[31:0] = int_wr_req_desc_9_wuser_12_wuser;
   assign uc2rb_wr_req_desc_9_wuser_13_reg[31:0] = int_wr_req_desc_9_wuser_13_wuser;
   assign uc2rb_wr_req_desc_9_wuser_14_reg[31:0] = int_wr_req_desc_9_wuser_14_wuser;
   assign uc2rb_wr_req_desc_9_wuser_15_reg[31:0] = int_wr_req_desc_9_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_9_resp_reg[4:0] = int_sn_resp_desc_9_resp_resp;
   assign uc2rb_rd_req_desc_a_size_reg[31:0] = int_rd_req_desc_a_size_txn_size;
   assign uc2rb_rd_req_desc_a_axsize_reg[2:0] = int_rd_req_desc_a_axsize_axsize;
   assign uc2rb_rd_req_desc_a_attr_reg[27:24] = int_rd_req_desc_a_attr_axsnoop;
   assign uc2rb_rd_req_desc_a_attr_reg[23:22] = int_rd_req_desc_a_attr_axdomain;
   assign uc2rb_rd_req_desc_a_attr_reg[21:20] = int_rd_req_desc_a_attr_axbar;
   assign uc2rb_rd_req_desc_a_attr_reg[18:15] = int_rd_req_desc_a_attr_axregion;
   assign uc2rb_rd_req_desc_a_attr_reg[14:11] = int_rd_req_desc_a_attr_axqos;
   assign uc2rb_rd_req_desc_a_attr_reg[10:8] = int_rd_req_desc_a_attr_axprot;
   assign uc2rb_rd_req_desc_a_attr_reg[7:4] = int_rd_req_desc_a_attr_axcache;
   assign uc2rb_rd_req_desc_a_attr_reg[2] = int_rd_req_desc_a_attr_axlock;
   assign uc2rb_rd_req_desc_a_attr_reg[1:0] = int_rd_req_desc_a_attr_axburst;
   assign uc2rb_rd_req_desc_a_axaddr_0_reg[31:0] = int_rd_req_desc_a_axaddr_0_addr;
   assign uc2rb_rd_req_desc_a_axaddr_1_reg[31:0] = int_rd_req_desc_a_axaddr_1_addr;
   assign uc2rb_rd_req_desc_a_axaddr_2_reg[31:0] = int_rd_req_desc_a_axaddr_2_addr;
   assign uc2rb_rd_req_desc_a_axaddr_3_reg[31:0] = int_rd_req_desc_a_axaddr_3_addr;
   assign uc2rb_rd_req_desc_a_axid_0_reg[31:0] = int_rd_req_desc_a_axid_0_axid;
   assign uc2rb_rd_req_desc_a_axid_1_reg[31:0] = int_rd_req_desc_a_axid_1_axid;
   assign uc2rb_rd_req_desc_a_axid_2_reg[31:0] = int_rd_req_desc_a_axid_2_axid;
   assign uc2rb_rd_req_desc_a_axid_3_reg[31:0] = int_rd_req_desc_a_axid_3_axid;
   assign uc2rb_rd_req_desc_a_axuser_0_reg[31:0] = int_rd_req_desc_a_axuser_0_axuser;
   assign uc2rb_rd_req_desc_a_axuser_1_reg[31:0] = int_rd_req_desc_a_axuser_1_axuser;
   assign uc2rb_rd_req_desc_a_axuser_2_reg[31:0] = int_rd_req_desc_a_axuser_2_axuser;
   assign uc2rb_rd_req_desc_a_axuser_3_reg[31:0] = int_rd_req_desc_a_axuser_3_axuser;
   assign uc2rb_rd_req_desc_a_axuser_4_reg[31:0] = int_rd_req_desc_a_axuser_4_axuser;
   assign uc2rb_rd_req_desc_a_axuser_5_reg[31:0] = int_rd_req_desc_a_axuser_5_axuser;
   assign uc2rb_rd_req_desc_a_axuser_6_reg[31:0] = int_rd_req_desc_a_axuser_6_axuser;
   assign uc2rb_rd_req_desc_a_axuser_7_reg[31:0] = int_rd_req_desc_a_axuser_7_axuser;
   assign uc2rb_rd_req_desc_a_axuser_8_reg[31:0] = int_rd_req_desc_a_axuser_8_axuser;
   assign uc2rb_rd_req_desc_a_axuser_9_reg[31:0] = int_rd_req_desc_a_axuser_9_axuser;
   assign uc2rb_rd_req_desc_a_axuser_10_reg[31:0] = int_rd_req_desc_a_axuser_10_axuser;
   assign uc2rb_rd_req_desc_a_axuser_11_reg[31:0] = int_rd_req_desc_a_axuser_11_axuser;
   assign uc2rb_rd_req_desc_a_axuser_12_reg[31:0] = int_rd_req_desc_a_axuser_12_axuser;
   assign uc2rb_rd_req_desc_a_axuser_13_reg[31:0] = int_rd_req_desc_a_axuser_13_axuser;
   assign uc2rb_rd_req_desc_a_axuser_14_reg[31:0] = int_rd_req_desc_a_axuser_14_axuser;
   assign uc2rb_rd_req_desc_a_axuser_15_reg[31:0] = int_rd_req_desc_a_axuser_15_axuser;
   assign uc2rb_wr_req_desc_a_txn_type_reg[1] = int_wr_req_desc_a_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_a_size_reg[31:0] = int_wr_req_desc_a_size_txn_size;
   assign uc2rb_wr_req_desc_a_data_offset_reg[13:0] = int_wr_req_desc_a_data_offset_addr;
   assign uc2rb_wr_req_desc_a_axsize_reg[2:0] = int_wr_req_desc_a_axsize_axsize;
   assign uc2rb_wr_req_desc_a_attr_reg[27:24] = int_wr_req_desc_a_attr_axsnoop;
   assign uc2rb_wr_req_desc_a_attr_reg[23:22] = int_wr_req_desc_a_attr_axdomain;
   assign uc2rb_wr_req_desc_a_attr_reg[21:20] = int_wr_req_desc_a_attr_axbar;
   assign uc2rb_wr_req_desc_a_attr_reg[19] = int_wr_req_desc_a_attr_awunique;
   assign uc2rb_wr_req_desc_a_attr_reg[18:15] = int_wr_req_desc_a_attr_axregion;
   assign uc2rb_wr_req_desc_a_attr_reg[14:11] = int_wr_req_desc_a_attr_axqos;
   assign uc2rb_wr_req_desc_a_attr_reg[10:8] = int_wr_req_desc_a_attr_axprot;
   assign uc2rb_wr_req_desc_a_attr_reg[7:4] = int_wr_req_desc_a_attr_axcache;
   assign uc2rb_wr_req_desc_a_attr_reg[2] = int_wr_req_desc_a_attr_axlock;
   assign uc2rb_wr_req_desc_a_attr_reg[1:0] = int_wr_req_desc_a_attr_axburst;
   assign uc2rb_wr_req_desc_a_axaddr_0_reg[31:0] = int_wr_req_desc_a_axaddr_0_addr;
   assign uc2rb_wr_req_desc_a_axaddr_1_reg[31:0] = int_wr_req_desc_a_axaddr_1_addr;
   assign uc2rb_wr_req_desc_a_axaddr_2_reg[31:0] = int_wr_req_desc_a_axaddr_2_addr;
   assign uc2rb_wr_req_desc_a_axaddr_3_reg[31:0] = int_wr_req_desc_a_axaddr_3_addr;
   assign uc2rb_wr_req_desc_a_axid_0_reg[31:0] = int_wr_req_desc_a_axid_0_axid;
   assign uc2rb_wr_req_desc_a_axid_1_reg[31:0] = int_wr_req_desc_a_axid_1_axid;
   assign uc2rb_wr_req_desc_a_axid_2_reg[31:0] = int_wr_req_desc_a_axid_2_axid;
   assign uc2rb_wr_req_desc_a_axid_3_reg[31:0] = int_wr_req_desc_a_axid_3_axid;
   assign uc2rb_wr_req_desc_a_axuser_0_reg[31:0] = int_wr_req_desc_a_axuser_0_axuser;
   assign uc2rb_wr_req_desc_a_axuser_1_reg[31:0] = int_wr_req_desc_a_axuser_1_axuser;
   assign uc2rb_wr_req_desc_a_axuser_2_reg[31:0] = int_wr_req_desc_a_axuser_2_axuser;
   assign uc2rb_wr_req_desc_a_axuser_3_reg[31:0] = int_wr_req_desc_a_axuser_3_axuser;
   assign uc2rb_wr_req_desc_a_axuser_4_reg[31:0] = int_wr_req_desc_a_axuser_4_axuser;
   assign uc2rb_wr_req_desc_a_axuser_5_reg[31:0] = int_wr_req_desc_a_axuser_5_axuser;
   assign uc2rb_wr_req_desc_a_axuser_6_reg[31:0] = int_wr_req_desc_a_axuser_6_axuser;
   assign uc2rb_wr_req_desc_a_axuser_7_reg[31:0] = int_wr_req_desc_a_axuser_7_axuser;
   assign uc2rb_wr_req_desc_a_axuser_8_reg[31:0] = int_wr_req_desc_a_axuser_8_axuser;
   assign uc2rb_wr_req_desc_a_axuser_9_reg[31:0] = int_wr_req_desc_a_axuser_9_axuser;
   assign uc2rb_wr_req_desc_a_axuser_10_reg[31:0] = int_wr_req_desc_a_axuser_10_axuser;
   assign uc2rb_wr_req_desc_a_axuser_11_reg[31:0] = int_wr_req_desc_a_axuser_11_axuser;
   assign uc2rb_wr_req_desc_a_axuser_12_reg[31:0] = int_wr_req_desc_a_axuser_12_axuser;
   assign uc2rb_wr_req_desc_a_axuser_13_reg[31:0] = int_wr_req_desc_a_axuser_13_axuser;
   assign uc2rb_wr_req_desc_a_axuser_14_reg[31:0] = int_wr_req_desc_a_axuser_14_axuser;
   assign uc2rb_wr_req_desc_a_axuser_15_reg[31:0] = int_wr_req_desc_a_axuser_15_axuser;
   assign uc2rb_wr_req_desc_a_wuser_0_reg[31:0] = int_wr_req_desc_a_wuser_0_wuser;
   assign uc2rb_wr_req_desc_a_wuser_1_reg[31:0] = int_wr_req_desc_a_wuser_1_wuser;
   assign uc2rb_wr_req_desc_a_wuser_2_reg[31:0] = int_wr_req_desc_a_wuser_2_wuser;
   assign uc2rb_wr_req_desc_a_wuser_3_reg[31:0] = int_wr_req_desc_a_wuser_3_wuser;
   assign uc2rb_wr_req_desc_a_wuser_4_reg[31:0] = int_wr_req_desc_a_wuser_4_wuser;
   assign uc2rb_wr_req_desc_a_wuser_5_reg[31:0] = int_wr_req_desc_a_wuser_5_wuser;
   assign uc2rb_wr_req_desc_a_wuser_6_reg[31:0] = int_wr_req_desc_a_wuser_6_wuser;
   assign uc2rb_wr_req_desc_a_wuser_7_reg[31:0] = int_wr_req_desc_a_wuser_7_wuser;
   assign uc2rb_wr_req_desc_a_wuser_8_reg[31:0] = int_wr_req_desc_a_wuser_8_wuser;
   assign uc2rb_wr_req_desc_a_wuser_9_reg[31:0] = int_wr_req_desc_a_wuser_9_wuser;
   assign uc2rb_wr_req_desc_a_wuser_10_reg[31:0] = int_wr_req_desc_a_wuser_10_wuser;
   assign uc2rb_wr_req_desc_a_wuser_11_reg[31:0] = int_wr_req_desc_a_wuser_11_wuser;
   assign uc2rb_wr_req_desc_a_wuser_12_reg[31:0] = int_wr_req_desc_a_wuser_12_wuser;
   assign uc2rb_wr_req_desc_a_wuser_13_reg[31:0] = int_wr_req_desc_a_wuser_13_wuser;
   assign uc2rb_wr_req_desc_a_wuser_14_reg[31:0] = int_wr_req_desc_a_wuser_14_wuser;
   assign uc2rb_wr_req_desc_a_wuser_15_reg[31:0] = int_wr_req_desc_a_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_a_resp_reg[4:0] = int_sn_resp_desc_a_resp_resp;
   assign uc2rb_rd_req_desc_b_size_reg[31:0] = int_rd_req_desc_b_size_txn_size;
   assign uc2rb_rd_req_desc_b_axsize_reg[2:0] = int_rd_req_desc_b_axsize_axsize;
   assign uc2rb_rd_req_desc_b_attr_reg[27:24] = int_rd_req_desc_b_attr_axsnoop;
   assign uc2rb_rd_req_desc_b_attr_reg[23:22] = int_rd_req_desc_b_attr_axdomain;
   assign uc2rb_rd_req_desc_b_attr_reg[21:20] = int_rd_req_desc_b_attr_axbar;
   assign uc2rb_rd_req_desc_b_attr_reg[18:15] = int_rd_req_desc_b_attr_axregion;
   assign uc2rb_rd_req_desc_b_attr_reg[14:11] = int_rd_req_desc_b_attr_axqos;
   assign uc2rb_rd_req_desc_b_attr_reg[10:8] = int_rd_req_desc_b_attr_axprot;
   assign uc2rb_rd_req_desc_b_attr_reg[7:4] = int_rd_req_desc_b_attr_axcache;
   assign uc2rb_rd_req_desc_b_attr_reg[2] = int_rd_req_desc_b_attr_axlock;
   assign uc2rb_rd_req_desc_b_attr_reg[1:0] = int_rd_req_desc_b_attr_axburst;
   assign uc2rb_rd_req_desc_b_axaddr_0_reg[31:0] = int_rd_req_desc_b_axaddr_0_addr;
   assign uc2rb_rd_req_desc_b_axaddr_1_reg[31:0] = int_rd_req_desc_b_axaddr_1_addr;
   assign uc2rb_rd_req_desc_b_axaddr_2_reg[31:0] = int_rd_req_desc_b_axaddr_2_addr;
   assign uc2rb_rd_req_desc_b_axaddr_3_reg[31:0] = int_rd_req_desc_b_axaddr_3_addr;
   assign uc2rb_rd_req_desc_b_axid_0_reg[31:0] = int_rd_req_desc_b_axid_0_axid;
   assign uc2rb_rd_req_desc_b_axid_1_reg[31:0] = int_rd_req_desc_b_axid_1_axid;
   assign uc2rb_rd_req_desc_b_axid_2_reg[31:0] = int_rd_req_desc_b_axid_2_axid;
   assign uc2rb_rd_req_desc_b_axid_3_reg[31:0] = int_rd_req_desc_b_axid_3_axid;
   assign uc2rb_rd_req_desc_b_axuser_0_reg[31:0] = int_rd_req_desc_b_axuser_0_axuser;
   assign uc2rb_rd_req_desc_b_axuser_1_reg[31:0] = int_rd_req_desc_b_axuser_1_axuser;
   assign uc2rb_rd_req_desc_b_axuser_2_reg[31:0] = int_rd_req_desc_b_axuser_2_axuser;
   assign uc2rb_rd_req_desc_b_axuser_3_reg[31:0] = int_rd_req_desc_b_axuser_3_axuser;
   assign uc2rb_rd_req_desc_b_axuser_4_reg[31:0] = int_rd_req_desc_b_axuser_4_axuser;
   assign uc2rb_rd_req_desc_b_axuser_5_reg[31:0] = int_rd_req_desc_b_axuser_5_axuser;
   assign uc2rb_rd_req_desc_b_axuser_6_reg[31:0] = int_rd_req_desc_b_axuser_6_axuser;
   assign uc2rb_rd_req_desc_b_axuser_7_reg[31:0] = int_rd_req_desc_b_axuser_7_axuser;
   assign uc2rb_rd_req_desc_b_axuser_8_reg[31:0] = int_rd_req_desc_b_axuser_8_axuser;
   assign uc2rb_rd_req_desc_b_axuser_9_reg[31:0] = int_rd_req_desc_b_axuser_9_axuser;
   assign uc2rb_rd_req_desc_b_axuser_10_reg[31:0] = int_rd_req_desc_b_axuser_10_axuser;
   assign uc2rb_rd_req_desc_b_axuser_11_reg[31:0] = int_rd_req_desc_b_axuser_11_axuser;
   assign uc2rb_rd_req_desc_b_axuser_12_reg[31:0] = int_rd_req_desc_b_axuser_12_axuser;
   assign uc2rb_rd_req_desc_b_axuser_13_reg[31:0] = int_rd_req_desc_b_axuser_13_axuser;
   assign uc2rb_rd_req_desc_b_axuser_14_reg[31:0] = int_rd_req_desc_b_axuser_14_axuser;
   assign uc2rb_rd_req_desc_b_axuser_15_reg[31:0] = int_rd_req_desc_b_axuser_15_axuser;
   assign uc2rb_wr_req_desc_b_txn_type_reg[1] = int_wr_req_desc_b_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_b_size_reg[31:0] = int_wr_req_desc_b_size_txn_size;
   assign uc2rb_wr_req_desc_b_data_offset_reg[13:0] = int_wr_req_desc_b_data_offset_addr;
   assign uc2rb_wr_req_desc_b_axsize_reg[2:0] = int_wr_req_desc_b_axsize_axsize;
   assign uc2rb_wr_req_desc_b_attr_reg[27:24] = int_wr_req_desc_b_attr_axsnoop;
   assign uc2rb_wr_req_desc_b_attr_reg[23:22] = int_wr_req_desc_b_attr_axdomain;
   assign uc2rb_wr_req_desc_b_attr_reg[21:20] = int_wr_req_desc_b_attr_axbar;
   assign uc2rb_wr_req_desc_b_attr_reg[19] = int_wr_req_desc_b_attr_awunique;
   assign uc2rb_wr_req_desc_b_attr_reg[18:15] = int_wr_req_desc_b_attr_axregion;
   assign uc2rb_wr_req_desc_b_attr_reg[14:11] = int_wr_req_desc_b_attr_axqos;
   assign uc2rb_wr_req_desc_b_attr_reg[10:8] = int_wr_req_desc_b_attr_axprot;
   assign uc2rb_wr_req_desc_b_attr_reg[7:4] = int_wr_req_desc_b_attr_axcache;
   assign uc2rb_wr_req_desc_b_attr_reg[2] = int_wr_req_desc_b_attr_axlock;
   assign uc2rb_wr_req_desc_b_attr_reg[1:0] = int_wr_req_desc_b_attr_axburst;
   assign uc2rb_wr_req_desc_b_axaddr_0_reg[31:0] = int_wr_req_desc_b_axaddr_0_addr;
   assign uc2rb_wr_req_desc_b_axaddr_1_reg[31:0] = int_wr_req_desc_b_axaddr_1_addr;
   assign uc2rb_wr_req_desc_b_axaddr_2_reg[31:0] = int_wr_req_desc_b_axaddr_2_addr;
   assign uc2rb_wr_req_desc_b_axaddr_3_reg[31:0] = int_wr_req_desc_b_axaddr_3_addr;
   assign uc2rb_wr_req_desc_b_axid_0_reg[31:0] = int_wr_req_desc_b_axid_0_axid;
   assign uc2rb_wr_req_desc_b_axid_1_reg[31:0] = int_wr_req_desc_b_axid_1_axid;
   assign uc2rb_wr_req_desc_b_axid_2_reg[31:0] = int_wr_req_desc_b_axid_2_axid;
   assign uc2rb_wr_req_desc_b_axid_3_reg[31:0] = int_wr_req_desc_b_axid_3_axid;
   assign uc2rb_wr_req_desc_b_axuser_0_reg[31:0] = int_wr_req_desc_b_axuser_0_axuser;
   assign uc2rb_wr_req_desc_b_axuser_1_reg[31:0] = int_wr_req_desc_b_axuser_1_axuser;
   assign uc2rb_wr_req_desc_b_axuser_2_reg[31:0] = int_wr_req_desc_b_axuser_2_axuser;
   assign uc2rb_wr_req_desc_b_axuser_3_reg[31:0] = int_wr_req_desc_b_axuser_3_axuser;
   assign uc2rb_wr_req_desc_b_axuser_4_reg[31:0] = int_wr_req_desc_b_axuser_4_axuser;
   assign uc2rb_wr_req_desc_b_axuser_5_reg[31:0] = int_wr_req_desc_b_axuser_5_axuser;
   assign uc2rb_wr_req_desc_b_axuser_6_reg[31:0] = int_wr_req_desc_b_axuser_6_axuser;
   assign uc2rb_wr_req_desc_b_axuser_7_reg[31:0] = int_wr_req_desc_b_axuser_7_axuser;
   assign uc2rb_wr_req_desc_b_axuser_8_reg[31:0] = int_wr_req_desc_b_axuser_8_axuser;
   assign uc2rb_wr_req_desc_b_axuser_9_reg[31:0] = int_wr_req_desc_b_axuser_9_axuser;
   assign uc2rb_wr_req_desc_b_axuser_10_reg[31:0] = int_wr_req_desc_b_axuser_10_axuser;
   assign uc2rb_wr_req_desc_b_axuser_11_reg[31:0] = int_wr_req_desc_b_axuser_11_axuser;
   assign uc2rb_wr_req_desc_b_axuser_12_reg[31:0] = int_wr_req_desc_b_axuser_12_axuser;
   assign uc2rb_wr_req_desc_b_axuser_13_reg[31:0] = int_wr_req_desc_b_axuser_13_axuser;
   assign uc2rb_wr_req_desc_b_axuser_14_reg[31:0] = int_wr_req_desc_b_axuser_14_axuser;
   assign uc2rb_wr_req_desc_b_axuser_15_reg[31:0] = int_wr_req_desc_b_axuser_15_axuser;
   assign uc2rb_wr_req_desc_b_wuser_0_reg[31:0] = int_wr_req_desc_b_wuser_0_wuser;
   assign uc2rb_wr_req_desc_b_wuser_1_reg[31:0] = int_wr_req_desc_b_wuser_1_wuser;
   assign uc2rb_wr_req_desc_b_wuser_2_reg[31:0] = int_wr_req_desc_b_wuser_2_wuser;
   assign uc2rb_wr_req_desc_b_wuser_3_reg[31:0] = int_wr_req_desc_b_wuser_3_wuser;
   assign uc2rb_wr_req_desc_b_wuser_4_reg[31:0] = int_wr_req_desc_b_wuser_4_wuser;
   assign uc2rb_wr_req_desc_b_wuser_5_reg[31:0] = int_wr_req_desc_b_wuser_5_wuser;
   assign uc2rb_wr_req_desc_b_wuser_6_reg[31:0] = int_wr_req_desc_b_wuser_6_wuser;
   assign uc2rb_wr_req_desc_b_wuser_7_reg[31:0] = int_wr_req_desc_b_wuser_7_wuser;
   assign uc2rb_wr_req_desc_b_wuser_8_reg[31:0] = int_wr_req_desc_b_wuser_8_wuser;
   assign uc2rb_wr_req_desc_b_wuser_9_reg[31:0] = int_wr_req_desc_b_wuser_9_wuser;
   assign uc2rb_wr_req_desc_b_wuser_10_reg[31:0] = int_wr_req_desc_b_wuser_10_wuser;
   assign uc2rb_wr_req_desc_b_wuser_11_reg[31:0] = int_wr_req_desc_b_wuser_11_wuser;
   assign uc2rb_wr_req_desc_b_wuser_12_reg[31:0] = int_wr_req_desc_b_wuser_12_wuser;
   assign uc2rb_wr_req_desc_b_wuser_13_reg[31:0] = int_wr_req_desc_b_wuser_13_wuser;
   assign uc2rb_wr_req_desc_b_wuser_14_reg[31:0] = int_wr_req_desc_b_wuser_14_wuser;
   assign uc2rb_wr_req_desc_b_wuser_15_reg[31:0] = int_wr_req_desc_b_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_b_resp_reg[4:0] = int_sn_resp_desc_b_resp_resp;
   assign uc2rb_rd_req_desc_c_size_reg[31:0] = int_rd_req_desc_c_size_txn_size;
   assign uc2rb_rd_req_desc_c_axsize_reg[2:0] = int_rd_req_desc_c_axsize_axsize;
   assign uc2rb_rd_req_desc_c_attr_reg[27:24] = int_rd_req_desc_c_attr_axsnoop;
   assign uc2rb_rd_req_desc_c_attr_reg[23:22] = int_rd_req_desc_c_attr_axdomain;
   assign uc2rb_rd_req_desc_c_attr_reg[21:20] = int_rd_req_desc_c_attr_axbar;
   assign uc2rb_rd_req_desc_c_attr_reg[18:15] = int_rd_req_desc_c_attr_axregion;
   assign uc2rb_rd_req_desc_c_attr_reg[14:11] = int_rd_req_desc_c_attr_axqos;
   assign uc2rb_rd_req_desc_c_attr_reg[10:8] = int_rd_req_desc_c_attr_axprot;
   assign uc2rb_rd_req_desc_c_attr_reg[7:4] = int_rd_req_desc_c_attr_axcache;
   assign uc2rb_rd_req_desc_c_attr_reg[2] = int_rd_req_desc_c_attr_axlock;
   assign uc2rb_rd_req_desc_c_attr_reg[1:0] = int_rd_req_desc_c_attr_axburst;
   assign uc2rb_rd_req_desc_c_axaddr_0_reg[31:0] = int_rd_req_desc_c_axaddr_0_addr;
   assign uc2rb_rd_req_desc_c_axaddr_1_reg[31:0] = int_rd_req_desc_c_axaddr_1_addr;
   assign uc2rb_rd_req_desc_c_axaddr_2_reg[31:0] = int_rd_req_desc_c_axaddr_2_addr;
   assign uc2rb_rd_req_desc_c_axaddr_3_reg[31:0] = int_rd_req_desc_c_axaddr_3_addr;
   assign uc2rb_rd_req_desc_c_axid_0_reg[31:0] = int_rd_req_desc_c_axid_0_axid;
   assign uc2rb_rd_req_desc_c_axid_1_reg[31:0] = int_rd_req_desc_c_axid_1_axid;
   assign uc2rb_rd_req_desc_c_axid_2_reg[31:0] = int_rd_req_desc_c_axid_2_axid;
   assign uc2rb_rd_req_desc_c_axid_3_reg[31:0] = int_rd_req_desc_c_axid_3_axid;
   assign uc2rb_rd_req_desc_c_axuser_0_reg[31:0] = int_rd_req_desc_c_axuser_0_axuser;
   assign uc2rb_rd_req_desc_c_axuser_1_reg[31:0] = int_rd_req_desc_c_axuser_1_axuser;
   assign uc2rb_rd_req_desc_c_axuser_2_reg[31:0] = int_rd_req_desc_c_axuser_2_axuser;
   assign uc2rb_rd_req_desc_c_axuser_3_reg[31:0] = int_rd_req_desc_c_axuser_3_axuser;
   assign uc2rb_rd_req_desc_c_axuser_4_reg[31:0] = int_rd_req_desc_c_axuser_4_axuser;
   assign uc2rb_rd_req_desc_c_axuser_5_reg[31:0] = int_rd_req_desc_c_axuser_5_axuser;
   assign uc2rb_rd_req_desc_c_axuser_6_reg[31:0] = int_rd_req_desc_c_axuser_6_axuser;
   assign uc2rb_rd_req_desc_c_axuser_7_reg[31:0] = int_rd_req_desc_c_axuser_7_axuser;
   assign uc2rb_rd_req_desc_c_axuser_8_reg[31:0] = int_rd_req_desc_c_axuser_8_axuser;
   assign uc2rb_rd_req_desc_c_axuser_9_reg[31:0] = int_rd_req_desc_c_axuser_9_axuser;
   assign uc2rb_rd_req_desc_c_axuser_10_reg[31:0] = int_rd_req_desc_c_axuser_10_axuser;
   assign uc2rb_rd_req_desc_c_axuser_11_reg[31:0] = int_rd_req_desc_c_axuser_11_axuser;
   assign uc2rb_rd_req_desc_c_axuser_12_reg[31:0] = int_rd_req_desc_c_axuser_12_axuser;
   assign uc2rb_rd_req_desc_c_axuser_13_reg[31:0] = int_rd_req_desc_c_axuser_13_axuser;
   assign uc2rb_rd_req_desc_c_axuser_14_reg[31:0] = int_rd_req_desc_c_axuser_14_axuser;
   assign uc2rb_rd_req_desc_c_axuser_15_reg[31:0] = int_rd_req_desc_c_axuser_15_axuser;
   assign uc2rb_wr_req_desc_c_txn_type_reg[1] = int_wr_req_desc_c_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_c_size_reg[31:0] = int_wr_req_desc_c_size_txn_size;
   assign uc2rb_wr_req_desc_c_data_offset_reg[13:0] = int_wr_req_desc_c_data_offset_addr;
   assign uc2rb_wr_req_desc_c_axsize_reg[2:0] = int_wr_req_desc_c_axsize_axsize;
   assign uc2rb_wr_req_desc_c_attr_reg[27:24] = int_wr_req_desc_c_attr_axsnoop;
   assign uc2rb_wr_req_desc_c_attr_reg[23:22] = int_wr_req_desc_c_attr_axdomain;
   assign uc2rb_wr_req_desc_c_attr_reg[21:20] = int_wr_req_desc_c_attr_axbar;
   assign uc2rb_wr_req_desc_c_attr_reg[19] = int_wr_req_desc_c_attr_awunique;
   assign uc2rb_wr_req_desc_c_attr_reg[18:15] = int_wr_req_desc_c_attr_axregion;
   assign uc2rb_wr_req_desc_c_attr_reg[14:11] = int_wr_req_desc_c_attr_axqos;
   assign uc2rb_wr_req_desc_c_attr_reg[10:8] = int_wr_req_desc_c_attr_axprot;
   assign uc2rb_wr_req_desc_c_attr_reg[7:4] = int_wr_req_desc_c_attr_axcache;
   assign uc2rb_wr_req_desc_c_attr_reg[2] = int_wr_req_desc_c_attr_axlock;
   assign uc2rb_wr_req_desc_c_attr_reg[1:0] = int_wr_req_desc_c_attr_axburst;
   assign uc2rb_wr_req_desc_c_axaddr_0_reg[31:0] = int_wr_req_desc_c_axaddr_0_addr;
   assign uc2rb_wr_req_desc_c_axaddr_1_reg[31:0] = int_wr_req_desc_c_axaddr_1_addr;
   assign uc2rb_wr_req_desc_c_axaddr_2_reg[31:0] = int_wr_req_desc_c_axaddr_2_addr;
   assign uc2rb_wr_req_desc_c_axaddr_3_reg[31:0] = int_wr_req_desc_c_axaddr_3_addr;
   assign uc2rb_wr_req_desc_c_axid_0_reg[31:0] = int_wr_req_desc_c_axid_0_axid;
   assign uc2rb_wr_req_desc_c_axid_1_reg[31:0] = int_wr_req_desc_c_axid_1_axid;
   assign uc2rb_wr_req_desc_c_axid_2_reg[31:0] = int_wr_req_desc_c_axid_2_axid;
   assign uc2rb_wr_req_desc_c_axid_3_reg[31:0] = int_wr_req_desc_c_axid_3_axid;
   assign uc2rb_wr_req_desc_c_axuser_0_reg[31:0] = int_wr_req_desc_c_axuser_0_axuser;
   assign uc2rb_wr_req_desc_c_axuser_1_reg[31:0] = int_wr_req_desc_c_axuser_1_axuser;
   assign uc2rb_wr_req_desc_c_axuser_2_reg[31:0] = int_wr_req_desc_c_axuser_2_axuser;
   assign uc2rb_wr_req_desc_c_axuser_3_reg[31:0] = int_wr_req_desc_c_axuser_3_axuser;
   assign uc2rb_wr_req_desc_c_axuser_4_reg[31:0] = int_wr_req_desc_c_axuser_4_axuser;
   assign uc2rb_wr_req_desc_c_axuser_5_reg[31:0] = int_wr_req_desc_c_axuser_5_axuser;
   assign uc2rb_wr_req_desc_c_axuser_6_reg[31:0] = int_wr_req_desc_c_axuser_6_axuser;
   assign uc2rb_wr_req_desc_c_axuser_7_reg[31:0] = int_wr_req_desc_c_axuser_7_axuser;
   assign uc2rb_wr_req_desc_c_axuser_8_reg[31:0] = int_wr_req_desc_c_axuser_8_axuser;
   assign uc2rb_wr_req_desc_c_axuser_9_reg[31:0] = int_wr_req_desc_c_axuser_9_axuser;
   assign uc2rb_wr_req_desc_c_axuser_10_reg[31:0] = int_wr_req_desc_c_axuser_10_axuser;
   assign uc2rb_wr_req_desc_c_axuser_11_reg[31:0] = int_wr_req_desc_c_axuser_11_axuser;
   assign uc2rb_wr_req_desc_c_axuser_12_reg[31:0] = int_wr_req_desc_c_axuser_12_axuser;
   assign uc2rb_wr_req_desc_c_axuser_13_reg[31:0] = int_wr_req_desc_c_axuser_13_axuser;
   assign uc2rb_wr_req_desc_c_axuser_14_reg[31:0] = int_wr_req_desc_c_axuser_14_axuser;
   assign uc2rb_wr_req_desc_c_axuser_15_reg[31:0] = int_wr_req_desc_c_axuser_15_axuser;
   assign uc2rb_wr_req_desc_c_wuser_0_reg[31:0] = int_wr_req_desc_c_wuser_0_wuser;
   assign uc2rb_wr_req_desc_c_wuser_1_reg[31:0] = int_wr_req_desc_c_wuser_1_wuser;
   assign uc2rb_wr_req_desc_c_wuser_2_reg[31:0] = int_wr_req_desc_c_wuser_2_wuser;
   assign uc2rb_wr_req_desc_c_wuser_3_reg[31:0] = int_wr_req_desc_c_wuser_3_wuser;
   assign uc2rb_wr_req_desc_c_wuser_4_reg[31:0] = int_wr_req_desc_c_wuser_4_wuser;
   assign uc2rb_wr_req_desc_c_wuser_5_reg[31:0] = int_wr_req_desc_c_wuser_5_wuser;
   assign uc2rb_wr_req_desc_c_wuser_6_reg[31:0] = int_wr_req_desc_c_wuser_6_wuser;
   assign uc2rb_wr_req_desc_c_wuser_7_reg[31:0] = int_wr_req_desc_c_wuser_7_wuser;
   assign uc2rb_wr_req_desc_c_wuser_8_reg[31:0] = int_wr_req_desc_c_wuser_8_wuser;
   assign uc2rb_wr_req_desc_c_wuser_9_reg[31:0] = int_wr_req_desc_c_wuser_9_wuser;
   assign uc2rb_wr_req_desc_c_wuser_10_reg[31:0] = int_wr_req_desc_c_wuser_10_wuser;
   assign uc2rb_wr_req_desc_c_wuser_11_reg[31:0] = int_wr_req_desc_c_wuser_11_wuser;
   assign uc2rb_wr_req_desc_c_wuser_12_reg[31:0] = int_wr_req_desc_c_wuser_12_wuser;
   assign uc2rb_wr_req_desc_c_wuser_13_reg[31:0] = int_wr_req_desc_c_wuser_13_wuser;
   assign uc2rb_wr_req_desc_c_wuser_14_reg[31:0] = int_wr_req_desc_c_wuser_14_wuser;
   assign uc2rb_wr_req_desc_c_wuser_15_reg[31:0] = int_wr_req_desc_c_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_c_resp_reg[4:0] = int_sn_resp_desc_c_resp_resp;
   assign uc2rb_rd_req_desc_d_size_reg[31:0] = int_rd_req_desc_d_size_txn_size;
   assign uc2rb_rd_req_desc_d_axsize_reg[2:0] = int_rd_req_desc_d_axsize_axsize;
   assign uc2rb_rd_req_desc_d_attr_reg[27:24] = int_rd_req_desc_d_attr_axsnoop;
   assign uc2rb_rd_req_desc_d_attr_reg[23:22] = int_rd_req_desc_d_attr_axdomain;
   assign uc2rb_rd_req_desc_d_attr_reg[21:20] = int_rd_req_desc_d_attr_axbar;
   assign uc2rb_rd_req_desc_d_attr_reg[18:15] = int_rd_req_desc_d_attr_axregion;
   assign uc2rb_rd_req_desc_d_attr_reg[14:11] = int_rd_req_desc_d_attr_axqos;
   assign uc2rb_rd_req_desc_d_attr_reg[10:8] = int_rd_req_desc_d_attr_axprot;
   assign uc2rb_rd_req_desc_d_attr_reg[7:4] = int_rd_req_desc_d_attr_axcache;
   assign uc2rb_rd_req_desc_d_attr_reg[2] = int_rd_req_desc_d_attr_axlock;
   assign uc2rb_rd_req_desc_d_attr_reg[1:0] = int_rd_req_desc_d_attr_axburst;
   assign uc2rb_rd_req_desc_d_axaddr_0_reg[31:0] = int_rd_req_desc_d_axaddr_0_addr;
   assign uc2rb_rd_req_desc_d_axaddr_1_reg[31:0] = int_rd_req_desc_d_axaddr_1_addr;
   assign uc2rb_rd_req_desc_d_axaddr_2_reg[31:0] = int_rd_req_desc_d_axaddr_2_addr;
   assign uc2rb_rd_req_desc_d_axaddr_3_reg[31:0] = int_rd_req_desc_d_axaddr_3_addr;
   assign uc2rb_rd_req_desc_d_axid_0_reg[31:0] = int_rd_req_desc_d_axid_0_axid;
   assign uc2rb_rd_req_desc_d_axid_1_reg[31:0] = int_rd_req_desc_d_axid_1_axid;
   assign uc2rb_rd_req_desc_d_axid_2_reg[31:0] = int_rd_req_desc_d_axid_2_axid;
   assign uc2rb_rd_req_desc_d_axid_3_reg[31:0] = int_rd_req_desc_d_axid_3_axid;
   assign uc2rb_rd_req_desc_d_axuser_0_reg[31:0] = int_rd_req_desc_d_axuser_0_axuser;
   assign uc2rb_rd_req_desc_d_axuser_1_reg[31:0] = int_rd_req_desc_d_axuser_1_axuser;
   assign uc2rb_rd_req_desc_d_axuser_2_reg[31:0] = int_rd_req_desc_d_axuser_2_axuser;
   assign uc2rb_rd_req_desc_d_axuser_3_reg[31:0] = int_rd_req_desc_d_axuser_3_axuser;
   assign uc2rb_rd_req_desc_d_axuser_4_reg[31:0] = int_rd_req_desc_d_axuser_4_axuser;
   assign uc2rb_rd_req_desc_d_axuser_5_reg[31:0] = int_rd_req_desc_d_axuser_5_axuser;
   assign uc2rb_rd_req_desc_d_axuser_6_reg[31:0] = int_rd_req_desc_d_axuser_6_axuser;
   assign uc2rb_rd_req_desc_d_axuser_7_reg[31:0] = int_rd_req_desc_d_axuser_7_axuser;
   assign uc2rb_rd_req_desc_d_axuser_8_reg[31:0] = int_rd_req_desc_d_axuser_8_axuser;
   assign uc2rb_rd_req_desc_d_axuser_9_reg[31:0] = int_rd_req_desc_d_axuser_9_axuser;
   assign uc2rb_rd_req_desc_d_axuser_10_reg[31:0] = int_rd_req_desc_d_axuser_10_axuser;
   assign uc2rb_rd_req_desc_d_axuser_11_reg[31:0] = int_rd_req_desc_d_axuser_11_axuser;
   assign uc2rb_rd_req_desc_d_axuser_12_reg[31:0] = int_rd_req_desc_d_axuser_12_axuser;
   assign uc2rb_rd_req_desc_d_axuser_13_reg[31:0] = int_rd_req_desc_d_axuser_13_axuser;
   assign uc2rb_rd_req_desc_d_axuser_14_reg[31:0] = int_rd_req_desc_d_axuser_14_axuser;
   assign uc2rb_rd_req_desc_d_axuser_15_reg[31:0] = int_rd_req_desc_d_axuser_15_axuser;
   assign uc2rb_wr_req_desc_d_txn_type_reg[1] = int_wr_req_desc_d_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_d_size_reg[31:0] = int_wr_req_desc_d_size_txn_size;
   assign uc2rb_wr_req_desc_d_data_offset_reg[13:0] = int_wr_req_desc_d_data_offset_addr;
   assign uc2rb_wr_req_desc_d_axsize_reg[2:0] = int_wr_req_desc_d_axsize_axsize;
   assign uc2rb_wr_req_desc_d_attr_reg[27:24] = int_wr_req_desc_d_attr_axsnoop;
   assign uc2rb_wr_req_desc_d_attr_reg[23:22] = int_wr_req_desc_d_attr_axdomain;
   assign uc2rb_wr_req_desc_d_attr_reg[21:20] = int_wr_req_desc_d_attr_axbar;
   assign uc2rb_wr_req_desc_d_attr_reg[19] = int_wr_req_desc_d_attr_awunique;
   assign uc2rb_wr_req_desc_d_attr_reg[18:15] = int_wr_req_desc_d_attr_axregion;
   assign uc2rb_wr_req_desc_d_attr_reg[14:11] = int_wr_req_desc_d_attr_axqos;
   assign uc2rb_wr_req_desc_d_attr_reg[10:8] = int_wr_req_desc_d_attr_axprot;
   assign uc2rb_wr_req_desc_d_attr_reg[7:4] = int_wr_req_desc_d_attr_axcache;
   assign uc2rb_wr_req_desc_d_attr_reg[2] = int_wr_req_desc_d_attr_axlock;
   assign uc2rb_wr_req_desc_d_attr_reg[1:0] = int_wr_req_desc_d_attr_axburst;
   assign uc2rb_wr_req_desc_d_axaddr_0_reg[31:0] = int_wr_req_desc_d_axaddr_0_addr;
   assign uc2rb_wr_req_desc_d_axaddr_1_reg[31:0] = int_wr_req_desc_d_axaddr_1_addr;
   assign uc2rb_wr_req_desc_d_axaddr_2_reg[31:0] = int_wr_req_desc_d_axaddr_2_addr;
   assign uc2rb_wr_req_desc_d_axaddr_3_reg[31:0] = int_wr_req_desc_d_axaddr_3_addr;
   assign uc2rb_wr_req_desc_d_axid_0_reg[31:0] = int_wr_req_desc_d_axid_0_axid;
   assign uc2rb_wr_req_desc_d_axid_1_reg[31:0] = int_wr_req_desc_d_axid_1_axid;
   assign uc2rb_wr_req_desc_d_axid_2_reg[31:0] = int_wr_req_desc_d_axid_2_axid;
   assign uc2rb_wr_req_desc_d_axid_3_reg[31:0] = int_wr_req_desc_d_axid_3_axid;
   assign uc2rb_wr_req_desc_d_axuser_0_reg[31:0] = int_wr_req_desc_d_axuser_0_axuser;
   assign uc2rb_wr_req_desc_d_axuser_1_reg[31:0] = int_wr_req_desc_d_axuser_1_axuser;
   assign uc2rb_wr_req_desc_d_axuser_2_reg[31:0] = int_wr_req_desc_d_axuser_2_axuser;
   assign uc2rb_wr_req_desc_d_axuser_3_reg[31:0] = int_wr_req_desc_d_axuser_3_axuser;
   assign uc2rb_wr_req_desc_d_axuser_4_reg[31:0] = int_wr_req_desc_d_axuser_4_axuser;
   assign uc2rb_wr_req_desc_d_axuser_5_reg[31:0] = int_wr_req_desc_d_axuser_5_axuser;
   assign uc2rb_wr_req_desc_d_axuser_6_reg[31:0] = int_wr_req_desc_d_axuser_6_axuser;
   assign uc2rb_wr_req_desc_d_axuser_7_reg[31:0] = int_wr_req_desc_d_axuser_7_axuser;
   assign uc2rb_wr_req_desc_d_axuser_8_reg[31:0] = int_wr_req_desc_d_axuser_8_axuser;
   assign uc2rb_wr_req_desc_d_axuser_9_reg[31:0] = int_wr_req_desc_d_axuser_9_axuser;
   assign uc2rb_wr_req_desc_d_axuser_10_reg[31:0] = int_wr_req_desc_d_axuser_10_axuser;
   assign uc2rb_wr_req_desc_d_axuser_11_reg[31:0] = int_wr_req_desc_d_axuser_11_axuser;
   assign uc2rb_wr_req_desc_d_axuser_12_reg[31:0] = int_wr_req_desc_d_axuser_12_axuser;
   assign uc2rb_wr_req_desc_d_axuser_13_reg[31:0] = int_wr_req_desc_d_axuser_13_axuser;
   assign uc2rb_wr_req_desc_d_axuser_14_reg[31:0] = int_wr_req_desc_d_axuser_14_axuser;
   assign uc2rb_wr_req_desc_d_axuser_15_reg[31:0] = int_wr_req_desc_d_axuser_15_axuser;
   assign uc2rb_wr_req_desc_d_wuser_0_reg[31:0] = int_wr_req_desc_d_wuser_0_wuser;
   assign uc2rb_wr_req_desc_d_wuser_1_reg[31:0] = int_wr_req_desc_d_wuser_1_wuser;
   assign uc2rb_wr_req_desc_d_wuser_2_reg[31:0] = int_wr_req_desc_d_wuser_2_wuser;
   assign uc2rb_wr_req_desc_d_wuser_3_reg[31:0] = int_wr_req_desc_d_wuser_3_wuser;
   assign uc2rb_wr_req_desc_d_wuser_4_reg[31:0] = int_wr_req_desc_d_wuser_4_wuser;
   assign uc2rb_wr_req_desc_d_wuser_5_reg[31:0] = int_wr_req_desc_d_wuser_5_wuser;
   assign uc2rb_wr_req_desc_d_wuser_6_reg[31:0] = int_wr_req_desc_d_wuser_6_wuser;
   assign uc2rb_wr_req_desc_d_wuser_7_reg[31:0] = int_wr_req_desc_d_wuser_7_wuser;
   assign uc2rb_wr_req_desc_d_wuser_8_reg[31:0] = int_wr_req_desc_d_wuser_8_wuser;
   assign uc2rb_wr_req_desc_d_wuser_9_reg[31:0] = int_wr_req_desc_d_wuser_9_wuser;
   assign uc2rb_wr_req_desc_d_wuser_10_reg[31:0] = int_wr_req_desc_d_wuser_10_wuser;
   assign uc2rb_wr_req_desc_d_wuser_11_reg[31:0] = int_wr_req_desc_d_wuser_11_wuser;
   assign uc2rb_wr_req_desc_d_wuser_12_reg[31:0] = int_wr_req_desc_d_wuser_12_wuser;
   assign uc2rb_wr_req_desc_d_wuser_13_reg[31:0] = int_wr_req_desc_d_wuser_13_wuser;
   assign uc2rb_wr_req_desc_d_wuser_14_reg[31:0] = int_wr_req_desc_d_wuser_14_wuser;
   assign uc2rb_wr_req_desc_d_wuser_15_reg[31:0] = int_wr_req_desc_d_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_d_resp_reg[4:0] = int_sn_resp_desc_d_resp_resp;
   assign uc2rb_rd_req_desc_e_size_reg[31:0] = int_rd_req_desc_e_size_txn_size;
   assign uc2rb_rd_req_desc_e_axsize_reg[2:0] = int_rd_req_desc_e_axsize_axsize;
   assign uc2rb_rd_req_desc_e_attr_reg[27:24] = int_rd_req_desc_e_attr_axsnoop;
   assign uc2rb_rd_req_desc_e_attr_reg[23:22] = int_rd_req_desc_e_attr_axdomain;
   assign uc2rb_rd_req_desc_e_attr_reg[21:20] = int_rd_req_desc_e_attr_axbar;
   assign uc2rb_rd_req_desc_e_attr_reg[18:15] = int_rd_req_desc_e_attr_axregion;
   assign uc2rb_rd_req_desc_e_attr_reg[14:11] = int_rd_req_desc_e_attr_axqos;
   assign uc2rb_rd_req_desc_e_attr_reg[10:8] = int_rd_req_desc_e_attr_axprot;
   assign uc2rb_rd_req_desc_e_attr_reg[7:4] = int_rd_req_desc_e_attr_axcache;
   assign uc2rb_rd_req_desc_e_attr_reg[2] = int_rd_req_desc_e_attr_axlock;
   assign uc2rb_rd_req_desc_e_attr_reg[1:0] = int_rd_req_desc_e_attr_axburst;
   assign uc2rb_rd_req_desc_e_axaddr_0_reg[31:0] = int_rd_req_desc_e_axaddr_0_addr;
   assign uc2rb_rd_req_desc_e_axaddr_1_reg[31:0] = int_rd_req_desc_e_axaddr_1_addr;
   assign uc2rb_rd_req_desc_e_axaddr_2_reg[31:0] = int_rd_req_desc_e_axaddr_2_addr;
   assign uc2rb_rd_req_desc_e_axaddr_3_reg[31:0] = int_rd_req_desc_e_axaddr_3_addr;
   assign uc2rb_rd_req_desc_e_axid_0_reg[31:0] = int_rd_req_desc_e_axid_0_axid;
   assign uc2rb_rd_req_desc_e_axid_1_reg[31:0] = int_rd_req_desc_e_axid_1_axid;
   assign uc2rb_rd_req_desc_e_axid_2_reg[31:0] = int_rd_req_desc_e_axid_2_axid;
   assign uc2rb_rd_req_desc_e_axid_3_reg[31:0] = int_rd_req_desc_e_axid_3_axid;
   assign uc2rb_rd_req_desc_e_axuser_0_reg[31:0] = int_rd_req_desc_e_axuser_0_axuser;
   assign uc2rb_rd_req_desc_e_axuser_1_reg[31:0] = int_rd_req_desc_e_axuser_1_axuser;
   assign uc2rb_rd_req_desc_e_axuser_2_reg[31:0] = int_rd_req_desc_e_axuser_2_axuser;
   assign uc2rb_rd_req_desc_e_axuser_3_reg[31:0] = int_rd_req_desc_e_axuser_3_axuser;
   assign uc2rb_rd_req_desc_e_axuser_4_reg[31:0] = int_rd_req_desc_e_axuser_4_axuser;
   assign uc2rb_rd_req_desc_e_axuser_5_reg[31:0] = int_rd_req_desc_e_axuser_5_axuser;
   assign uc2rb_rd_req_desc_e_axuser_6_reg[31:0] = int_rd_req_desc_e_axuser_6_axuser;
   assign uc2rb_rd_req_desc_e_axuser_7_reg[31:0] = int_rd_req_desc_e_axuser_7_axuser;
   assign uc2rb_rd_req_desc_e_axuser_8_reg[31:0] = int_rd_req_desc_e_axuser_8_axuser;
   assign uc2rb_rd_req_desc_e_axuser_9_reg[31:0] = int_rd_req_desc_e_axuser_9_axuser;
   assign uc2rb_rd_req_desc_e_axuser_10_reg[31:0] = int_rd_req_desc_e_axuser_10_axuser;
   assign uc2rb_rd_req_desc_e_axuser_11_reg[31:0] = int_rd_req_desc_e_axuser_11_axuser;
   assign uc2rb_rd_req_desc_e_axuser_12_reg[31:0] = int_rd_req_desc_e_axuser_12_axuser;
   assign uc2rb_rd_req_desc_e_axuser_13_reg[31:0] = int_rd_req_desc_e_axuser_13_axuser;
   assign uc2rb_rd_req_desc_e_axuser_14_reg[31:0] = int_rd_req_desc_e_axuser_14_axuser;
   assign uc2rb_rd_req_desc_e_axuser_15_reg[31:0] = int_rd_req_desc_e_axuser_15_axuser;
   assign uc2rb_wr_req_desc_e_txn_type_reg[1] = int_wr_req_desc_e_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_e_size_reg[31:0] = int_wr_req_desc_e_size_txn_size;
   assign uc2rb_wr_req_desc_e_data_offset_reg[13:0] = int_wr_req_desc_e_data_offset_addr;
   assign uc2rb_wr_req_desc_e_axsize_reg[2:0] = int_wr_req_desc_e_axsize_axsize;
   assign uc2rb_wr_req_desc_e_attr_reg[27:24] = int_wr_req_desc_e_attr_axsnoop;
   assign uc2rb_wr_req_desc_e_attr_reg[23:22] = int_wr_req_desc_e_attr_axdomain;
   assign uc2rb_wr_req_desc_e_attr_reg[21:20] = int_wr_req_desc_e_attr_axbar;
   assign uc2rb_wr_req_desc_e_attr_reg[19] = int_wr_req_desc_e_attr_awunique;
   assign uc2rb_wr_req_desc_e_attr_reg[18:15] = int_wr_req_desc_e_attr_axregion;
   assign uc2rb_wr_req_desc_e_attr_reg[14:11] = int_wr_req_desc_e_attr_axqos;
   assign uc2rb_wr_req_desc_e_attr_reg[10:8] = int_wr_req_desc_e_attr_axprot;
   assign uc2rb_wr_req_desc_e_attr_reg[7:4] = int_wr_req_desc_e_attr_axcache;
   assign uc2rb_wr_req_desc_e_attr_reg[2] = int_wr_req_desc_e_attr_axlock;
   assign uc2rb_wr_req_desc_e_attr_reg[1:0] = int_wr_req_desc_e_attr_axburst;
   assign uc2rb_wr_req_desc_e_axaddr_0_reg[31:0] = int_wr_req_desc_e_axaddr_0_addr;
   assign uc2rb_wr_req_desc_e_axaddr_1_reg[31:0] = int_wr_req_desc_e_axaddr_1_addr;
   assign uc2rb_wr_req_desc_e_axaddr_2_reg[31:0] = int_wr_req_desc_e_axaddr_2_addr;
   assign uc2rb_wr_req_desc_e_axaddr_3_reg[31:0] = int_wr_req_desc_e_axaddr_3_addr;
   assign uc2rb_wr_req_desc_e_axid_0_reg[31:0] = int_wr_req_desc_e_axid_0_axid;
   assign uc2rb_wr_req_desc_e_axid_1_reg[31:0] = int_wr_req_desc_e_axid_1_axid;
   assign uc2rb_wr_req_desc_e_axid_2_reg[31:0] = int_wr_req_desc_e_axid_2_axid;
   assign uc2rb_wr_req_desc_e_axid_3_reg[31:0] = int_wr_req_desc_e_axid_3_axid;
   assign uc2rb_wr_req_desc_e_axuser_0_reg[31:0] = int_wr_req_desc_e_axuser_0_axuser;
   assign uc2rb_wr_req_desc_e_axuser_1_reg[31:0] = int_wr_req_desc_e_axuser_1_axuser;
   assign uc2rb_wr_req_desc_e_axuser_2_reg[31:0] = int_wr_req_desc_e_axuser_2_axuser;
   assign uc2rb_wr_req_desc_e_axuser_3_reg[31:0] = int_wr_req_desc_e_axuser_3_axuser;
   assign uc2rb_wr_req_desc_e_axuser_4_reg[31:0] = int_wr_req_desc_e_axuser_4_axuser;
   assign uc2rb_wr_req_desc_e_axuser_5_reg[31:0] = int_wr_req_desc_e_axuser_5_axuser;
   assign uc2rb_wr_req_desc_e_axuser_6_reg[31:0] = int_wr_req_desc_e_axuser_6_axuser;
   assign uc2rb_wr_req_desc_e_axuser_7_reg[31:0] = int_wr_req_desc_e_axuser_7_axuser;
   assign uc2rb_wr_req_desc_e_axuser_8_reg[31:0] = int_wr_req_desc_e_axuser_8_axuser;
   assign uc2rb_wr_req_desc_e_axuser_9_reg[31:0] = int_wr_req_desc_e_axuser_9_axuser;
   assign uc2rb_wr_req_desc_e_axuser_10_reg[31:0] = int_wr_req_desc_e_axuser_10_axuser;
   assign uc2rb_wr_req_desc_e_axuser_11_reg[31:0] = int_wr_req_desc_e_axuser_11_axuser;
   assign uc2rb_wr_req_desc_e_axuser_12_reg[31:0] = int_wr_req_desc_e_axuser_12_axuser;
   assign uc2rb_wr_req_desc_e_axuser_13_reg[31:0] = int_wr_req_desc_e_axuser_13_axuser;
   assign uc2rb_wr_req_desc_e_axuser_14_reg[31:0] = int_wr_req_desc_e_axuser_14_axuser;
   assign uc2rb_wr_req_desc_e_axuser_15_reg[31:0] = int_wr_req_desc_e_axuser_15_axuser;
   assign uc2rb_wr_req_desc_e_wuser_0_reg[31:0] = int_wr_req_desc_e_wuser_0_wuser;
   assign uc2rb_wr_req_desc_e_wuser_1_reg[31:0] = int_wr_req_desc_e_wuser_1_wuser;
   assign uc2rb_wr_req_desc_e_wuser_2_reg[31:0] = int_wr_req_desc_e_wuser_2_wuser;
   assign uc2rb_wr_req_desc_e_wuser_3_reg[31:0] = int_wr_req_desc_e_wuser_3_wuser;
   assign uc2rb_wr_req_desc_e_wuser_4_reg[31:0] = int_wr_req_desc_e_wuser_4_wuser;
   assign uc2rb_wr_req_desc_e_wuser_5_reg[31:0] = int_wr_req_desc_e_wuser_5_wuser;
   assign uc2rb_wr_req_desc_e_wuser_6_reg[31:0] = int_wr_req_desc_e_wuser_6_wuser;
   assign uc2rb_wr_req_desc_e_wuser_7_reg[31:0] = int_wr_req_desc_e_wuser_7_wuser;
   assign uc2rb_wr_req_desc_e_wuser_8_reg[31:0] = int_wr_req_desc_e_wuser_8_wuser;
   assign uc2rb_wr_req_desc_e_wuser_9_reg[31:0] = int_wr_req_desc_e_wuser_9_wuser;
   assign uc2rb_wr_req_desc_e_wuser_10_reg[31:0] = int_wr_req_desc_e_wuser_10_wuser;
   assign uc2rb_wr_req_desc_e_wuser_11_reg[31:0] = int_wr_req_desc_e_wuser_11_wuser;
   assign uc2rb_wr_req_desc_e_wuser_12_reg[31:0] = int_wr_req_desc_e_wuser_12_wuser;
   assign uc2rb_wr_req_desc_e_wuser_13_reg[31:0] = int_wr_req_desc_e_wuser_13_wuser;
   assign uc2rb_wr_req_desc_e_wuser_14_reg[31:0] = int_wr_req_desc_e_wuser_14_wuser;
   assign uc2rb_wr_req_desc_e_wuser_15_reg[31:0] = int_wr_req_desc_e_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_e_resp_reg[4:0] = int_sn_resp_desc_e_resp_resp;
   assign uc2rb_rd_req_desc_f_size_reg[31:0] = int_rd_req_desc_f_size_txn_size;
   assign uc2rb_rd_req_desc_f_axsize_reg[2:0] = int_rd_req_desc_f_axsize_axsize;
   assign uc2rb_rd_req_desc_f_attr_reg[27:24] = int_rd_req_desc_f_attr_axsnoop;
   assign uc2rb_rd_req_desc_f_attr_reg[23:22] = int_rd_req_desc_f_attr_axdomain;
   assign uc2rb_rd_req_desc_f_attr_reg[21:20] = int_rd_req_desc_f_attr_axbar;
   assign uc2rb_rd_req_desc_f_attr_reg[18:15] = int_rd_req_desc_f_attr_axregion;
   assign uc2rb_rd_req_desc_f_attr_reg[14:11] = int_rd_req_desc_f_attr_axqos;
   assign uc2rb_rd_req_desc_f_attr_reg[10:8] = int_rd_req_desc_f_attr_axprot;
   assign uc2rb_rd_req_desc_f_attr_reg[7:4] = int_rd_req_desc_f_attr_axcache;
   assign uc2rb_rd_req_desc_f_attr_reg[2] = int_rd_req_desc_f_attr_axlock;
   assign uc2rb_rd_req_desc_f_attr_reg[1:0] = int_rd_req_desc_f_attr_axburst;
   assign uc2rb_rd_req_desc_f_axaddr_0_reg[31:0] = int_rd_req_desc_f_axaddr_0_addr;
   assign uc2rb_rd_req_desc_f_axaddr_1_reg[31:0] = int_rd_req_desc_f_axaddr_1_addr;
   assign uc2rb_rd_req_desc_f_axaddr_2_reg[31:0] = int_rd_req_desc_f_axaddr_2_addr;
   assign uc2rb_rd_req_desc_f_axaddr_3_reg[31:0] = int_rd_req_desc_f_axaddr_3_addr;
   assign uc2rb_rd_req_desc_f_axid_0_reg[31:0] = int_rd_req_desc_f_axid_0_axid;
   assign uc2rb_rd_req_desc_f_axid_1_reg[31:0] = int_rd_req_desc_f_axid_1_axid;
   assign uc2rb_rd_req_desc_f_axid_2_reg[31:0] = int_rd_req_desc_f_axid_2_axid;
   assign uc2rb_rd_req_desc_f_axid_3_reg[31:0] = int_rd_req_desc_f_axid_3_axid;
   assign uc2rb_rd_req_desc_f_axuser_0_reg[31:0] = int_rd_req_desc_f_axuser_0_axuser;
   assign uc2rb_rd_req_desc_f_axuser_1_reg[31:0] = int_rd_req_desc_f_axuser_1_axuser;
   assign uc2rb_rd_req_desc_f_axuser_2_reg[31:0] = int_rd_req_desc_f_axuser_2_axuser;
   assign uc2rb_rd_req_desc_f_axuser_3_reg[31:0] = int_rd_req_desc_f_axuser_3_axuser;
   assign uc2rb_rd_req_desc_f_axuser_4_reg[31:0] = int_rd_req_desc_f_axuser_4_axuser;
   assign uc2rb_rd_req_desc_f_axuser_5_reg[31:0] = int_rd_req_desc_f_axuser_5_axuser;
   assign uc2rb_rd_req_desc_f_axuser_6_reg[31:0] = int_rd_req_desc_f_axuser_6_axuser;
   assign uc2rb_rd_req_desc_f_axuser_7_reg[31:0] = int_rd_req_desc_f_axuser_7_axuser;
   assign uc2rb_rd_req_desc_f_axuser_8_reg[31:0] = int_rd_req_desc_f_axuser_8_axuser;
   assign uc2rb_rd_req_desc_f_axuser_9_reg[31:0] = int_rd_req_desc_f_axuser_9_axuser;
   assign uc2rb_rd_req_desc_f_axuser_10_reg[31:0] = int_rd_req_desc_f_axuser_10_axuser;
   assign uc2rb_rd_req_desc_f_axuser_11_reg[31:0] = int_rd_req_desc_f_axuser_11_axuser;
   assign uc2rb_rd_req_desc_f_axuser_12_reg[31:0] = int_rd_req_desc_f_axuser_12_axuser;
   assign uc2rb_rd_req_desc_f_axuser_13_reg[31:0] = int_rd_req_desc_f_axuser_13_axuser;
   assign uc2rb_rd_req_desc_f_axuser_14_reg[31:0] = int_rd_req_desc_f_axuser_14_axuser;
   assign uc2rb_rd_req_desc_f_axuser_15_reg[31:0] = int_rd_req_desc_f_axuser_15_axuser;
   assign uc2rb_wr_req_desc_f_txn_type_reg[1] = int_wr_req_desc_f_txn_type_wr_strb;
   assign uc2rb_wr_req_desc_f_size_reg[31:0] = int_wr_req_desc_f_size_txn_size;
   assign uc2rb_wr_req_desc_f_data_offset_reg[13:0] = int_wr_req_desc_f_data_offset_addr;
   assign uc2rb_wr_req_desc_f_axsize_reg[2:0] = int_wr_req_desc_f_axsize_axsize;
   assign uc2rb_wr_req_desc_f_attr_reg[27:24] = int_wr_req_desc_f_attr_axsnoop;
   assign uc2rb_wr_req_desc_f_attr_reg[23:22] = int_wr_req_desc_f_attr_axdomain;
   assign uc2rb_wr_req_desc_f_attr_reg[21:20] = int_wr_req_desc_f_attr_axbar;
   assign uc2rb_wr_req_desc_f_attr_reg[19] = int_wr_req_desc_f_attr_awunique;
   assign uc2rb_wr_req_desc_f_attr_reg[18:15] = int_wr_req_desc_f_attr_axregion;
   assign uc2rb_wr_req_desc_f_attr_reg[14:11] = int_wr_req_desc_f_attr_axqos;
   assign uc2rb_wr_req_desc_f_attr_reg[10:8] = int_wr_req_desc_f_attr_axprot;
   assign uc2rb_wr_req_desc_f_attr_reg[7:4] = int_wr_req_desc_f_attr_axcache;
   assign uc2rb_wr_req_desc_f_attr_reg[2] = int_wr_req_desc_f_attr_axlock;
   assign uc2rb_wr_req_desc_f_attr_reg[1:0] = int_wr_req_desc_f_attr_axburst;
   assign uc2rb_wr_req_desc_f_axaddr_0_reg[31:0] = int_wr_req_desc_f_axaddr_0_addr;
   assign uc2rb_wr_req_desc_f_axaddr_1_reg[31:0] = int_wr_req_desc_f_axaddr_1_addr;
   assign uc2rb_wr_req_desc_f_axaddr_2_reg[31:0] = int_wr_req_desc_f_axaddr_2_addr;
   assign uc2rb_wr_req_desc_f_axaddr_3_reg[31:0] = int_wr_req_desc_f_axaddr_3_addr;
   assign uc2rb_wr_req_desc_f_axid_0_reg[31:0] = int_wr_req_desc_f_axid_0_axid;
   assign uc2rb_wr_req_desc_f_axid_1_reg[31:0] = int_wr_req_desc_f_axid_1_axid;
   assign uc2rb_wr_req_desc_f_axid_2_reg[31:0] = int_wr_req_desc_f_axid_2_axid;
   assign uc2rb_wr_req_desc_f_axid_3_reg[31:0] = int_wr_req_desc_f_axid_3_axid;
   assign uc2rb_wr_req_desc_f_axuser_0_reg[31:0] = int_wr_req_desc_f_axuser_0_axuser;
   assign uc2rb_wr_req_desc_f_axuser_1_reg[31:0] = int_wr_req_desc_f_axuser_1_axuser;
   assign uc2rb_wr_req_desc_f_axuser_2_reg[31:0] = int_wr_req_desc_f_axuser_2_axuser;
   assign uc2rb_wr_req_desc_f_axuser_3_reg[31:0] = int_wr_req_desc_f_axuser_3_axuser;
   assign uc2rb_wr_req_desc_f_axuser_4_reg[31:0] = int_wr_req_desc_f_axuser_4_axuser;
   assign uc2rb_wr_req_desc_f_axuser_5_reg[31:0] = int_wr_req_desc_f_axuser_5_axuser;
   assign uc2rb_wr_req_desc_f_axuser_6_reg[31:0] = int_wr_req_desc_f_axuser_6_axuser;
   assign uc2rb_wr_req_desc_f_axuser_7_reg[31:0] = int_wr_req_desc_f_axuser_7_axuser;
   assign uc2rb_wr_req_desc_f_axuser_8_reg[31:0] = int_wr_req_desc_f_axuser_8_axuser;
   assign uc2rb_wr_req_desc_f_axuser_9_reg[31:0] = int_wr_req_desc_f_axuser_9_axuser;
   assign uc2rb_wr_req_desc_f_axuser_10_reg[31:0] = int_wr_req_desc_f_axuser_10_axuser;
   assign uc2rb_wr_req_desc_f_axuser_11_reg[31:0] = int_wr_req_desc_f_axuser_11_axuser;
   assign uc2rb_wr_req_desc_f_axuser_12_reg[31:0] = int_wr_req_desc_f_axuser_12_axuser;
   assign uc2rb_wr_req_desc_f_axuser_13_reg[31:0] = int_wr_req_desc_f_axuser_13_axuser;
   assign uc2rb_wr_req_desc_f_axuser_14_reg[31:0] = int_wr_req_desc_f_axuser_14_axuser;
   assign uc2rb_wr_req_desc_f_axuser_15_reg[31:0] = int_wr_req_desc_f_axuser_15_axuser;
   assign uc2rb_wr_req_desc_f_wuser_0_reg[31:0] = int_wr_req_desc_f_wuser_0_wuser;
   assign uc2rb_wr_req_desc_f_wuser_1_reg[31:0] = int_wr_req_desc_f_wuser_1_wuser;
   assign uc2rb_wr_req_desc_f_wuser_2_reg[31:0] = int_wr_req_desc_f_wuser_2_wuser;
   assign uc2rb_wr_req_desc_f_wuser_3_reg[31:0] = int_wr_req_desc_f_wuser_3_wuser;
   assign uc2rb_wr_req_desc_f_wuser_4_reg[31:0] = int_wr_req_desc_f_wuser_4_wuser;
   assign uc2rb_wr_req_desc_f_wuser_5_reg[31:0] = int_wr_req_desc_f_wuser_5_wuser;
   assign uc2rb_wr_req_desc_f_wuser_6_reg[31:0] = int_wr_req_desc_f_wuser_6_wuser;
   assign uc2rb_wr_req_desc_f_wuser_7_reg[31:0] = int_wr_req_desc_f_wuser_7_wuser;
   assign uc2rb_wr_req_desc_f_wuser_8_reg[31:0] = int_wr_req_desc_f_wuser_8_wuser;
   assign uc2rb_wr_req_desc_f_wuser_9_reg[31:0] = int_wr_req_desc_f_wuser_9_wuser;
   assign uc2rb_wr_req_desc_f_wuser_10_reg[31:0] = int_wr_req_desc_f_wuser_10_wuser;
   assign uc2rb_wr_req_desc_f_wuser_11_reg[31:0] = int_wr_req_desc_f_wuser_11_wuser;
   assign uc2rb_wr_req_desc_f_wuser_12_reg[31:0] = int_wr_req_desc_f_wuser_12_wuser;
   assign uc2rb_wr_req_desc_f_wuser_13_reg[31:0] = int_wr_req_desc_f_wuser_13_wuser;
   assign uc2rb_wr_req_desc_f_wuser_14_reg[31:0] = int_wr_req_desc_f_wuser_14_wuser;
   assign uc2rb_wr_req_desc_f_wuser_15_reg[31:0] = int_wr_req_desc_f_wuser_15_wuser;
   assign uc2rb_sn_resp_desc_f_resp_reg[4:0] = int_sn_resp_desc_f_resp_resp;
   assign uc2rb_rd_req_fifo_pop_desc_reg[30:4] = 'h0;
   assign uc2rb_rd_req_fifo_fill_level_reg[31:5] = 'h0;
   assign uc2rb_rd_resp_fifo_free_level_reg[31:5] = 'h0;
   assign uc2rb_rd_resp_intr_comp_status_reg[31:16] = 'h0;
   assign uc2rb_wr_req_fifo_pop_desc_reg[30:4] = 'h0;
   assign uc2rb_wr_req_fifo_fill_level_reg[31:5] = 'h0;
   assign uc2rb_wr_resp_fifo_free_level_reg[31:5] = 'h0;
   assign uc2rb_wr_resp_intr_comp_status_reg[31:16] = 'h0;
   assign uc2rb_sn_req_fifo_free_level_reg[31:5] = 'h0;
   assign uc2rb_sn_req_intr_comp_status_reg[31:16] = 'h0;
   assign uc2rb_sn_resp_fifo_pop_desc_reg[30:4] = 'h0;
   assign uc2rb_sn_resp_fifo_fill_level_reg[31:5] = 'h0;
   assign uc2rb_sn_data_fifo_pop_desc_reg[30:4] = 'h0;
   assign uc2rb_sn_data_fifo_fill_level_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_0_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_0_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_0_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_0_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_0_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_0_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_0_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_0_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_0_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_0_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_0_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_0_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_0_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_0_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_1_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_1_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_1_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_1_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_1_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_1_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_1_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_1_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_1_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_1_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_1_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_1_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_1_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_1_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_2_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_2_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_2_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_2_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_2_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_2_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_2_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_2_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_2_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_2_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_2_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_2_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_2_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_2_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_3_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_3_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_3_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_3_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_3_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_3_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_3_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_3_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_3_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_3_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_3_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_3_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_3_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_3_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_4_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_4_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_4_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_4_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_4_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_4_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_4_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_4_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_4_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_4_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_4_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_4_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_4_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_4_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_5_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_5_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_5_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_5_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_5_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_5_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_5_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_5_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_5_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_5_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_5_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_5_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_5_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_5_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_6_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_6_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_6_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_6_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_6_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_6_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_6_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_6_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_6_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_6_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_6_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_6_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_6_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_6_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_7_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_7_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_7_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_7_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_7_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_7_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_7_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_7_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_7_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_7_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_7_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_7_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_7_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_7_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_8_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_8_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_8_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_8_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_8_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_8_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_8_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_8_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_8_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_8_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_8_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_8_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_8_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_8_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_9_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_9_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_9_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_9_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_9_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_9_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_9_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_9_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_9_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_9_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_9_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_9_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_9_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_9_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_a_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_a_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_a_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_a_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_a_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_a_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_a_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_a_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_a_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_a_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_a_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_a_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_a_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_a_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_b_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_b_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_b_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_b_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_b_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_b_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_b_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_b_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_b_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_b_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_b_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_b_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_b_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_b_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_c_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_c_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_c_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_c_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_c_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_c_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_c_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_c_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_c_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_c_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_c_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_c_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_c_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_c_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_d_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_d_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_d_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_d_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_d_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_d_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_d_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_d_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_d_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_d_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_d_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_d_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_d_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_d_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_e_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_e_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_e_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_e_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_e_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_e_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_e_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_e_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_e_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_e_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_e_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_e_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_e_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_e_resp_reg[31:5] = 'h0;
   assign uc2rb_rd_req_desc_f_txn_type_reg[31:2] = 'h0;
   assign uc2rb_rd_req_desc_f_txn_type_reg[1] = 'h0;
   assign uc2rb_rd_req_desc_f_txn_type_reg[0] = 'h0;
   assign uc2rb_rd_req_desc_f_axsize_reg[31:3] = 'h0;
   assign uc2rb_rd_req_desc_f_attr_reg[31:28] = 'h0;
   assign uc2rb_rd_req_desc_f_attr_reg[19] = 'h0;
   assign uc2rb_rd_req_desc_f_attr_reg[3] = 'h0;
   assign uc2rb_wr_req_desc_f_txn_type_reg[31:2] = 'h0;
   assign uc2rb_wr_req_desc_f_txn_type_reg[0] = 'h0;
   assign uc2rb_wr_req_desc_f_data_offset_reg[31:14] = 'h0;
   assign uc2rb_wr_req_desc_f_axsize_reg[31:3] = 'h0;
   assign uc2rb_wr_req_desc_f_attr_reg[31:28] = 'h0;
   assign uc2rb_wr_req_desc_f_attr_reg[3] = 'h0;
   assign uc2rb_sn_resp_desc_f_resp_reg[31:5] = 'h0;


   //Tie all uc2rb_<reg>_reg_we to high because current implementation of uc2rb_<reg>_reg

   //such that it will always hold intended correct value.

   assign uc2rb_intr_error_status_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_fifo_pop_desc_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_fifo_fill_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_resp_fifo_free_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_resp_intr_comp_status_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_fifo_pop_desc_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_fifo_fill_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_resp_fifo_free_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_resp_intr_comp_status_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_req_fifo_free_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_req_intr_comp_status_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_fifo_pop_desc_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_fifo_fill_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_data_fifo_pop_desc_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_data_fifo_fill_level_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_0_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_0_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_0_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_1_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_1_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_1_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_2_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_2_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_2_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_3_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_3_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_3_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_4_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_4_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_4_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_5_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_5_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_5_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_6_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_6_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_6_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_7_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_7_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_7_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_8_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_8_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_8_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_9_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_9_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_9_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_a_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_a_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_a_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_b_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_b_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_b_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_c_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_c_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_c_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_d_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_d_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_d_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_e_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_e_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_e_resp_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_rd_req_desc_f_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_txn_type_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_size_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_data_offset_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axsize_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_attr_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axaddr_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axaddr_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axaddr_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axaddr_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axid_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axid_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axid_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axid_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_axuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_0_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_1_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_2_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_3_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_4_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_5_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_6_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_7_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_8_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_9_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_10_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_11_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_12_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_13_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_14_reg_we = 32'hFFFFFFFF;
   assign uc2rb_wr_req_desc_f_wuser_15_reg_we = 32'hFFFFFFFF;
   assign uc2rb_sn_resp_desc_f_resp_reg_we = 32'hFFFFFFFF;





   //////////////////////
   //Instantiate ace_slv_inf 
   //////////////////////
   
   ace_slv_inf #(
		  /*AUTOINSTPARAM*/
		  // Parameters
		  .ACE_PROTOCOL            (ACE_PROTOCOL),
		  .ADDR_WIDTH              (ADDR_WIDTH),
		  .XX_DATA_WIDTH           (XX_DATA_WIDTH),
		  .SN_DATA_WIDTH           (SN_DATA_WIDTH),
		  .ID_WIDTH                (ID_WIDTH),
		  .AWUSER_WIDTH            (AWUSER_WIDTH),
		  .WUSER_WIDTH             (WUSER_WIDTH),
		  .BUSER_WIDTH             (BUSER_WIDTH),
		  .ARUSER_WIDTH            (ARUSER_WIDTH),
		  .RUSER_WIDTH             (RUSER_WIDTH),
		  .CACHE_LINE_SIZE         (CACHE_LINE_SIZE),
		  .XX_MAX_DESC             (XX_MAX_DESC),
		  .SN_MAX_DESC             (SN_MAX_DESC),
		  .XX_RAM_SIZE             (XX_RAM_SIZE),
		  .SN_RAM_SIZE             (SN_RAM_SIZE))
   i_ace_slv_inf (
		   /*AUTOINST*/
                   // Outputs
                   .s_ace_usr_awready      (s_ace_usr_awready),
                   .s_ace_usr_wready       (s_ace_usr_wready),
                   .s_ace_usr_bid          (s_ace_usr_bid),
                   .s_ace_usr_bresp        (s_ace_usr_bresp),
                   .s_ace_usr_buser        (s_ace_usr_buser),
                   .s_ace_usr_bvalid       (s_ace_usr_bvalid),
                   .s_ace_usr_arready      (s_ace_usr_arready),
                   .s_ace_usr_rid          (s_ace_usr_rid),
                   .s_ace_usr_rdata        (s_ace_usr_rdata),
                   .s_ace_usr_rresp        (s_ace_usr_rresp),
                   .s_ace_usr_rlast        (s_ace_usr_rlast),
                   .s_ace_usr_ruser        (s_ace_usr_ruser),
                   .s_ace_usr_rvalid       (s_ace_usr_rvalid),
                   .s_ace_usr_acaddr       (s_ace_usr_acaddr),
                   .s_ace_usr_acsnoop      (s_ace_usr_acsnoop),
                   .s_ace_usr_acprot       (s_ace_usr_acprot),
                   .s_ace_usr_acvalid      (s_ace_usr_acvalid),
                   .s_ace_usr_crready      (s_ace_usr_crready),
                   .s_ace_usr_cdready      (s_ace_usr_cdready),
                   .uc2rb_rd_addr          (uc2rb_rd_addr),
                   .uc2rb_wr_we            (uc2rb_wr_we),
                   .uc2rb_wr_bwe           (uc2rb_wr_bwe),
                   .uc2rb_wr_addr          (uc2rb_wr_addr),
                   .uc2rb_wr_data          (uc2rb_wr_data),
                   .uc2rb_wr_wstrb         (uc2rb_wr_wstrb),
                   .uc2rb_sn_we            (uc2rb_sn_we),
                   .uc2rb_sn_bwe           (uc2rb_sn_bwe),
                   .uc2rb_sn_addr          (uc2rb_sn_addr),
                   .uc2rb_sn_data          (uc2rb_sn_data),
                   .rd_uc2hm_trig          (rd_uc2hm_trig),
                   .wr_uc2hm_trig          (wr_uc2hm_trig),
                   .int_intr_error_status_err_0(int_intr_error_status_err_0),
                   .int_rd_req_fifo_pop_desc_valid(int_rd_req_fifo_pop_desc_valid),
                   .int_rd_req_fifo_pop_desc_desc_index(int_rd_req_fifo_pop_desc_desc_index),
                   .int_rd_req_fifo_fill_level_fill(int_rd_req_fifo_fill_level_fill),
                   .int_rd_resp_fifo_free_level_free(int_rd_resp_fifo_free_level_free),
                   .int_rd_resp_intr_comp_status_comp(int_rd_resp_intr_comp_status_comp),
                   .int_wr_req_fifo_pop_desc_valid(int_wr_req_fifo_pop_desc_valid),
                   .int_wr_req_fifo_pop_desc_desc_index(int_wr_req_fifo_pop_desc_desc_index),
                   .int_wr_req_fifo_fill_level_fill(int_wr_req_fifo_fill_level_fill),
                   .int_wr_resp_fifo_free_level_free(int_wr_resp_fifo_free_level_free),
                   .int_wr_resp_intr_comp_status_comp(int_wr_resp_intr_comp_status_comp),
                   .int_sn_req_fifo_free_level_free(int_sn_req_fifo_free_level_free),
                   .int_sn_req_intr_comp_status_comp(int_sn_req_intr_comp_status_comp),
                   .int_sn_resp_fifo_pop_desc_valid(int_sn_resp_fifo_pop_desc_valid),
                   .int_sn_resp_fifo_pop_desc_desc_index(int_sn_resp_fifo_pop_desc_desc_index),
                   .int_sn_resp_fifo_fill_level_fill(int_sn_resp_fifo_fill_level_fill),
                   .int_sn_data_fifo_pop_desc_valid(int_sn_data_fifo_pop_desc_valid),
                   .int_sn_data_fifo_pop_desc_desc_index(int_sn_data_fifo_pop_desc_desc_index),
                   .int_sn_data_fifo_fill_level_fill(int_sn_data_fifo_fill_level_fill),
                   .int_rd_req_desc_0_size_txn_size(int_rd_req_desc_0_size_txn_size),
                   .int_rd_req_desc_0_axsize_axsize(int_rd_req_desc_0_axsize_axsize),
                   .int_rd_req_desc_0_attr_axsnoop(int_rd_req_desc_0_attr_axsnoop),
                   .int_rd_req_desc_0_attr_axdomain(int_rd_req_desc_0_attr_axdomain),
                   .int_rd_req_desc_0_attr_axbar(int_rd_req_desc_0_attr_axbar),
                   .int_rd_req_desc_0_attr_axregion(int_rd_req_desc_0_attr_axregion),
                   .int_rd_req_desc_0_attr_axqos(int_rd_req_desc_0_attr_axqos),
                   .int_rd_req_desc_0_attr_axprot(int_rd_req_desc_0_attr_axprot),
                   .int_rd_req_desc_0_attr_axcache(int_rd_req_desc_0_attr_axcache),
                   .int_rd_req_desc_0_attr_axlock(int_rd_req_desc_0_attr_axlock),
                   .int_rd_req_desc_0_attr_axburst(int_rd_req_desc_0_attr_axburst),
                   .int_rd_req_desc_0_axaddr_0_addr(int_rd_req_desc_0_axaddr_0_addr),
                   .int_rd_req_desc_0_axaddr_1_addr(int_rd_req_desc_0_axaddr_1_addr),
                   .int_rd_req_desc_0_axaddr_2_addr(int_rd_req_desc_0_axaddr_2_addr),
                   .int_rd_req_desc_0_axaddr_3_addr(int_rd_req_desc_0_axaddr_3_addr),
                   .int_rd_req_desc_0_axid_0_axid(int_rd_req_desc_0_axid_0_axid),
                   .int_rd_req_desc_0_axid_1_axid(int_rd_req_desc_0_axid_1_axid),
                   .int_rd_req_desc_0_axid_2_axid(int_rd_req_desc_0_axid_2_axid),
                   .int_rd_req_desc_0_axid_3_axid(int_rd_req_desc_0_axid_3_axid),
                   .int_rd_req_desc_0_axuser_0_axuser(int_rd_req_desc_0_axuser_0_axuser),
                   .int_rd_req_desc_0_axuser_1_axuser(int_rd_req_desc_0_axuser_1_axuser),
                   .int_rd_req_desc_0_axuser_2_axuser(int_rd_req_desc_0_axuser_2_axuser),
                   .int_rd_req_desc_0_axuser_3_axuser(int_rd_req_desc_0_axuser_3_axuser),
                   .int_rd_req_desc_0_axuser_4_axuser(int_rd_req_desc_0_axuser_4_axuser),
                   .int_rd_req_desc_0_axuser_5_axuser(int_rd_req_desc_0_axuser_5_axuser),
                   .int_rd_req_desc_0_axuser_6_axuser(int_rd_req_desc_0_axuser_6_axuser),
                   .int_rd_req_desc_0_axuser_7_axuser(int_rd_req_desc_0_axuser_7_axuser),
                   .int_rd_req_desc_0_axuser_8_axuser(int_rd_req_desc_0_axuser_8_axuser),
                   .int_rd_req_desc_0_axuser_9_axuser(int_rd_req_desc_0_axuser_9_axuser),
                   .int_rd_req_desc_0_axuser_10_axuser(int_rd_req_desc_0_axuser_10_axuser),
                   .int_rd_req_desc_0_axuser_11_axuser(int_rd_req_desc_0_axuser_11_axuser),
                   .int_rd_req_desc_0_axuser_12_axuser(int_rd_req_desc_0_axuser_12_axuser),
                   .int_rd_req_desc_0_axuser_13_axuser(int_rd_req_desc_0_axuser_13_axuser),
                   .int_rd_req_desc_0_axuser_14_axuser(int_rd_req_desc_0_axuser_14_axuser),
                   .int_rd_req_desc_0_axuser_15_axuser(int_rd_req_desc_0_axuser_15_axuser),
                   .int_wr_req_desc_0_txn_type_wr_strb(int_wr_req_desc_0_txn_type_wr_strb),
                   .int_wr_req_desc_0_size_txn_size(int_wr_req_desc_0_size_txn_size),
                   .int_wr_req_desc_0_data_offset_addr(int_wr_req_desc_0_data_offset_addr),
                   .int_wr_req_desc_0_axsize_axsize(int_wr_req_desc_0_axsize_axsize),
                   .int_wr_req_desc_0_attr_axsnoop(int_wr_req_desc_0_attr_axsnoop),
                   .int_wr_req_desc_0_attr_axdomain(int_wr_req_desc_0_attr_axdomain),
                   .int_wr_req_desc_0_attr_axbar(int_wr_req_desc_0_attr_axbar),
                   .int_wr_req_desc_0_attr_awunique(int_wr_req_desc_0_attr_awunique),
                   .int_wr_req_desc_0_attr_axregion(int_wr_req_desc_0_attr_axregion),
                   .int_wr_req_desc_0_attr_axqos(int_wr_req_desc_0_attr_axqos),
                   .int_wr_req_desc_0_attr_axprot(int_wr_req_desc_0_attr_axprot),
                   .int_wr_req_desc_0_attr_axcache(int_wr_req_desc_0_attr_axcache),
                   .int_wr_req_desc_0_attr_axlock(int_wr_req_desc_0_attr_axlock),
                   .int_wr_req_desc_0_attr_axburst(int_wr_req_desc_0_attr_axburst),
                   .int_wr_req_desc_0_axaddr_0_addr(int_wr_req_desc_0_axaddr_0_addr),
                   .int_wr_req_desc_0_axaddr_1_addr(int_wr_req_desc_0_axaddr_1_addr),
                   .int_wr_req_desc_0_axaddr_2_addr(int_wr_req_desc_0_axaddr_2_addr),
                   .int_wr_req_desc_0_axaddr_3_addr(int_wr_req_desc_0_axaddr_3_addr),
                   .int_wr_req_desc_0_axid_0_axid(int_wr_req_desc_0_axid_0_axid),
                   .int_wr_req_desc_0_axid_1_axid(int_wr_req_desc_0_axid_1_axid),
                   .int_wr_req_desc_0_axid_2_axid(int_wr_req_desc_0_axid_2_axid),
                   .int_wr_req_desc_0_axid_3_axid(int_wr_req_desc_0_axid_3_axid),
                   .int_wr_req_desc_0_axuser_0_axuser(int_wr_req_desc_0_axuser_0_axuser),
                   .int_wr_req_desc_0_axuser_1_axuser(int_wr_req_desc_0_axuser_1_axuser),
                   .int_wr_req_desc_0_axuser_2_axuser(int_wr_req_desc_0_axuser_2_axuser),
                   .int_wr_req_desc_0_axuser_3_axuser(int_wr_req_desc_0_axuser_3_axuser),
                   .int_wr_req_desc_0_axuser_4_axuser(int_wr_req_desc_0_axuser_4_axuser),
                   .int_wr_req_desc_0_axuser_5_axuser(int_wr_req_desc_0_axuser_5_axuser),
                   .int_wr_req_desc_0_axuser_6_axuser(int_wr_req_desc_0_axuser_6_axuser),
                   .int_wr_req_desc_0_axuser_7_axuser(int_wr_req_desc_0_axuser_7_axuser),
                   .int_wr_req_desc_0_axuser_8_axuser(int_wr_req_desc_0_axuser_8_axuser),
                   .int_wr_req_desc_0_axuser_9_axuser(int_wr_req_desc_0_axuser_9_axuser),
                   .int_wr_req_desc_0_axuser_10_axuser(int_wr_req_desc_0_axuser_10_axuser),
                   .int_wr_req_desc_0_axuser_11_axuser(int_wr_req_desc_0_axuser_11_axuser),
                   .int_wr_req_desc_0_axuser_12_axuser(int_wr_req_desc_0_axuser_12_axuser),
                   .int_wr_req_desc_0_axuser_13_axuser(int_wr_req_desc_0_axuser_13_axuser),
                   .int_wr_req_desc_0_axuser_14_axuser(int_wr_req_desc_0_axuser_14_axuser),
                   .int_wr_req_desc_0_axuser_15_axuser(int_wr_req_desc_0_axuser_15_axuser),
                   .int_wr_req_desc_0_wuser_0_wuser(int_wr_req_desc_0_wuser_0_wuser),
                   .int_wr_req_desc_0_wuser_1_wuser(int_wr_req_desc_0_wuser_1_wuser),
                   .int_wr_req_desc_0_wuser_2_wuser(int_wr_req_desc_0_wuser_2_wuser),
                   .int_wr_req_desc_0_wuser_3_wuser(int_wr_req_desc_0_wuser_3_wuser),
                   .int_wr_req_desc_0_wuser_4_wuser(int_wr_req_desc_0_wuser_4_wuser),
                   .int_wr_req_desc_0_wuser_5_wuser(int_wr_req_desc_0_wuser_5_wuser),
                   .int_wr_req_desc_0_wuser_6_wuser(int_wr_req_desc_0_wuser_6_wuser),
                   .int_wr_req_desc_0_wuser_7_wuser(int_wr_req_desc_0_wuser_7_wuser),
                   .int_wr_req_desc_0_wuser_8_wuser(int_wr_req_desc_0_wuser_8_wuser),
                   .int_wr_req_desc_0_wuser_9_wuser(int_wr_req_desc_0_wuser_9_wuser),
                   .int_wr_req_desc_0_wuser_10_wuser(int_wr_req_desc_0_wuser_10_wuser),
                   .int_wr_req_desc_0_wuser_11_wuser(int_wr_req_desc_0_wuser_11_wuser),
                   .int_wr_req_desc_0_wuser_12_wuser(int_wr_req_desc_0_wuser_12_wuser),
                   .int_wr_req_desc_0_wuser_13_wuser(int_wr_req_desc_0_wuser_13_wuser),
                   .int_wr_req_desc_0_wuser_14_wuser(int_wr_req_desc_0_wuser_14_wuser),
                   .int_wr_req_desc_0_wuser_15_wuser(int_wr_req_desc_0_wuser_15_wuser),
                   .int_sn_resp_desc_0_resp_resp(int_sn_resp_desc_0_resp_resp),
                   .int_rd_req_desc_1_size_txn_size(int_rd_req_desc_1_size_txn_size),
                   .int_rd_req_desc_1_axsize_axsize(int_rd_req_desc_1_axsize_axsize),
                   .int_rd_req_desc_1_attr_axsnoop(int_rd_req_desc_1_attr_axsnoop),
                   .int_rd_req_desc_1_attr_axdomain(int_rd_req_desc_1_attr_axdomain),
                   .int_rd_req_desc_1_attr_axbar(int_rd_req_desc_1_attr_axbar),
                   .int_rd_req_desc_1_attr_axregion(int_rd_req_desc_1_attr_axregion),
                   .int_rd_req_desc_1_attr_axqos(int_rd_req_desc_1_attr_axqos),
                   .int_rd_req_desc_1_attr_axprot(int_rd_req_desc_1_attr_axprot),
                   .int_rd_req_desc_1_attr_axcache(int_rd_req_desc_1_attr_axcache),
                   .int_rd_req_desc_1_attr_axlock(int_rd_req_desc_1_attr_axlock),
                   .int_rd_req_desc_1_attr_axburst(int_rd_req_desc_1_attr_axburst),
                   .int_rd_req_desc_1_axaddr_0_addr(int_rd_req_desc_1_axaddr_0_addr),
                   .int_rd_req_desc_1_axaddr_1_addr(int_rd_req_desc_1_axaddr_1_addr),
                   .int_rd_req_desc_1_axaddr_2_addr(int_rd_req_desc_1_axaddr_2_addr),
                   .int_rd_req_desc_1_axaddr_3_addr(int_rd_req_desc_1_axaddr_3_addr),
                   .int_rd_req_desc_1_axid_0_axid(int_rd_req_desc_1_axid_0_axid),
                   .int_rd_req_desc_1_axid_1_axid(int_rd_req_desc_1_axid_1_axid),
                   .int_rd_req_desc_1_axid_2_axid(int_rd_req_desc_1_axid_2_axid),
                   .int_rd_req_desc_1_axid_3_axid(int_rd_req_desc_1_axid_3_axid),
                   .int_rd_req_desc_1_axuser_0_axuser(int_rd_req_desc_1_axuser_0_axuser),
                   .int_rd_req_desc_1_axuser_1_axuser(int_rd_req_desc_1_axuser_1_axuser),
                   .int_rd_req_desc_1_axuser_2_axuser(int_rd_req_desc_1_axuser_2_axuser),
                   .int_rd_req_desc_1_axuser_3_axuser(int_rd_req_desc_1_axuser_3_axuser),
                   .int_rd_req_desc_1_axuser_4_axuser(int_rd_req_desc_1_axuser_4_axuser),
                   .int_rd_req_desc_1_axuser_5_axuser(int_rd_req_desc_1_axuser_5_axuser),
                   .int_rd_req_desc_1_axuser_6_axuser(int_rd_req_desc_1_axuser_6_axuser),
                   .int_rd_req_desc_1_axuser_7_axuser(int_rd_req_desc_1_axuser_7_axuser),
                   .int_rd_req_desc_1_axuser_8_axuser(int_rd_req_desc_1_axuser_8_axuser),
                   .int_rd_req_desc_1_axuser_9_axuser(int_rd_req_desc_1_axuser_9_axuser),
                   .int_rd_req_desc_1_axuser_10_axuser(int_rd_req_desc_1_axuser_10_axuser),
                   .int_rd_req_desc_1_axuser_11_axuser(int_rd_req_desc_1_axuser_11_axuser),
                   .int_rd_req_desc_1_axuser_12_axuser(int_rd_req_desc_1_axuser_12_axuser),
                   .int_rd_req_desc_1_axuser_13_axuser(int_rd_req_desc_1_axuser_13_axuser),
                   .int_rd_req_desc_1_axuser_14_axuser(int_rd_req_desc_1_axuser_14_axuser),
                   .int_rd_req_desc_1_axuser_15_axuser(int_rd_req_desc_1_axuser_15_axuser),
                   .int_wr_req_desc_1_txn_type_wr_strb(int_wr_req_desc_1_txn_type_wr_strb),
                   .int_wr_req_desc_1_size_txn_size(int_wr_req_desc_1_size_txn_size),
                   .int_wr_req_desc_1_data_offset_addr(int_wr_req_desc_1_data_offset_addr),
                   .int_wr_req_desc_1_axsize_axsize(int_wr_req_desc_1_axsize_axsize),
                   .int_wr_req_desc_1_attr_axsnoop(int_wr_req_desc_1_attr_axsnoop),
                   .int_wr_req_desc_1_attr_axdomain(int_wr_req_desc_1_attr_axdomain),
                   .int_wr_req_desc_1_attr_axbar(int_wr_req_desc_1_attr_axbar),
                   .int_wr_req_desc_1_attr_awunique(int_wr_req_desc_1_attr_awunique),
                   .int_wr_req_desc_1_attr_axregion(int_wr_req_desc_1_attr_axregion),
                   .int_wr_req_desc_1_attr_axqos(int_wr_req_desc_1_attr_axqos),
                   .int_wr_req_desc_1_attr_axprot(int_wr_req_desc_1_attr_axprot),
                   .int_wr_req_desc_1_attr_axcache(int_wr_req_desc_1_attr_axcache),
                   .int_wr_req_desc_1_attr_axlock(int_wr_req_desc_1_attr_axlock),
                   .int_wr_req_desc_1_attr_axburst(int_wr_req_desc_1_attr_axburst),
                   .int_wr_req_desc_1_axaddr_0_addr(int_wr_req_desc_1_axaddr_0_addr),
                   .int_wr_req_desc_1_axaddr_1_addr(int_wr_req_desc_1_axaddr_1_addr),
                   .int_wr_req_desc_1_axaddr_2_addr(int_wr_req_desc_1_axaddr_2_addr),
                   .int_wr_req_desc_1_axaddr_3_addr(int_wr_req_desc_1_axaddr_3_addr),
                   .int_wr_req_desc_1_axid_0_axid(int_wr_req_desc_1_axid_0_axid),
                   .int_wr_req_desc_1_axid_1_axid(int_wr_req_desc_1_axid_1_axid),
                   .int_wr_req_desc_1_axid_2_axid(int_wr_req_desc_1_axid_2_axid),
                   .int_wr_req_desc_1_axid_3_axid(int_wr_req_desc_1_axid_3_axid),
                   .int_wr_req_desc_1_axuser_0_axuser(int_wr_req_desc_1_axuser_0_axuser),
                   .int_wr_req_desc_1_axuser_1_axuser(int_wr_req_desc_1_axuser_1_axuser),
                   .int_wr_req_desc_1_axuser_2_axuser(int_wr_req_desc_1_axuser_2_axuser),
                   .int_wr_req_desc_1_axuser_3_axuser(int_wr_req_desc_1_axuser_3_axuser),
                   .int_wr_req_desc_1_axuser_4_axuser(int_wr_req_desc_1_axuser_4_axuser),
                   .int_wr_req_desc_1_axuser_5_axuser(int_wr_req_desc_1_axuser_5_axuser),
                   .int_wr_req_desc_1_axuser_6_axuser(int_wr_req_desc_1_axuser_6_axuser),
                   .int_wr_req_desc_1_axuser_7_axuser(int_wr_req_desc_1_axuser_7_axuser),
                   .int_wr_req_desc_1_axuser_8_axuser(int_wr_req_desc_1_axuser_8_axuser),
                   .int_wr_req_desc_1_axuser_9_axuser(int_wr_req_desc_1_axuser_9_axuser),
                   .int_wr_req_desc_1_axuser_10_axuser(int_wr_req_desc_1_axuser_10_axuser),
                   .int_wr_req_desc_1_axuser_11_axuser(int_wr_req_desc_1_axuser_11_axuser),
                   .int_wr_req_desc_1_axuser_12_axuser(int_wr_req_desc_1_axuser_12_axuser),
                   .int_wr_req_desc_1_axuser_13_axuser(int_wr_req_desc_1_axuser_13_axuser),
                   .int_wr_req_desc_1_axuser_14_axuser(int_wr_req_desc_1_axuser_14_axuser),
                   .int_wr_req_desc_1_axuser_15_axuser(int_wr_req_desc_1_axuser_15_axuser),
                   .int_wr_req_desc_1_wuser_0_wuser(int_wr_req_desc_1_wuser_0_wuser),
                   .int_wr_req_desc_1_wuser_1_wuser(int_wr_req_desc_1_wuser_1_wuser),
                   .int_wr_req_desc_1_wuser_2_wuser(int_wr_req_desc_1_wuser_2_wuser),
                   .int_wr_req_desc_1_wuser_3_wuser(int_wr_req_desc_1_wuser_3_wuser),
                   .int_wr_req_desc_1_wuser_4_wuser(int_wr_req_desc_1_wuser_4_wuser),
                   .int_wr_req_desc_1_wuser_5_wuser(int_wr_req_desc_1_wuser_5_wuser),
                   .int_wr_req_desc_1_wuser_6_wuser(int_wr_req_desc_1_wuser_6_wuser),
                   .int_wr_req_desc_1_wuser_7_wuser(int_wr_req_desc_1_wuser_7_wuser),
                   .int_wr_req_desc_1_wuser_8_wuser(int_wr_req_desc_1_wuser_8_wuser),
                   .int_wr_req_desc_1_wuser_9_wuser(int_wr_req_desc_1_wuser_9_wuser),
                   .int_wr_req_desc_1_wuser_10_wuser(int_wr_req_desc_1_wuser_10_wuser),
                   .int_wr_req_desc_1_wuser_11_wuser(int_wr_req_desc_1_wuser_11_wuser),
                   .int_wr_req_desc_1_wuser_12_wuser(int_wr_req_desc_1_wuser_12_wuser),
                   .int_wr_req_desc_1_wuser_13_wuser(int_wr_req_desc_1_wuser_13_wuser),
                   .int_wr_req_desc_1_wuser_14_wuser(int_wr_req_desc_1_wuser_14_wuser),
                   .int_wr_req_desc_1_wuser_15_wuser(int_wr_req_desc_1_wuser_15_wuser),
                   .int_sn_resp_desc_1_resp_resp(int_sn_resp_desc_1_resp_resp),
                   .int_rd_req_desc_2_size_txn_size(int_rd_req_desc_2_size_txn_size),
                   .int_rd_req_desc_2_axsize_axsize(int_rd_req_desc_2_axsize_axsize),
                   .int_rd_req_desc_2_attr_axsnoop(int_rd_req_desc_2_attr_axsnoop),
                   .int_rd_req_desc_2_attr_axdomain(int_rd_req_desc_2_attr_axdomain),
                   .int_rd_req_desc_2_attr_axbar(int_rd_req_desc_2_attr_axbar),
                   .int_rd_req_desc_2_attr_axregion(int_rd_req_desc_2_attr_axregion),
                   .int_rd_req_desc_2_attr_axqos(int_rd_req_desc_2_attr_axqos),
                   .int_rd_req_desc_2_attr_axprot(int_rd_req_desc_2_attr_axprot),
                   .int_rd_req_desc_2_attr_axcache(int_rd_req_desc_2_attr_axcache),
                   .int_rd_req_desc_2_attr_axlock(int_rd_req_desc_2_attr_axlock),
                   .int_rd_req_desc_2_attr_axburst(int_rd_req_desc_2_attr_axburst),
                   .int_rd_req_desc_2_axaddr_0_addr(int_rd_req_desc_2_axaddr_0_addr),
                   .int_rd_req_desc_2_axaddr_1_addr(int_rd_req_desc_2_axaddr_1_addr),
                   .int_rd_req_desc_2_axaddr_2_addr(int_rd_req_desc_2_axaddr_2_addr),
                   .int_rd_req_desc_2_axaddr_3_addr(int_rd_req_desc_2_axaddr_3_addr),
                   .int_rd_req_desc_2_axid_0_axid(int_rd_req_desc_2_axid_0_axid),
                   .int_rd_req_desc_2_axid_1_axid(int_rd_req_desc_2_axid_1_axid),
                   .int_rd_req_desc_2_axid_2_axid(int_rd_req_desc_2_axid_2_axid),
                   .int_rd_req_desc_2_axid_3_axid(int_rd_req_desc_2_axid_3_axid),
                   .int_rd_req_desc_2_axuser_0_axuser(int_rd_req_desc_2_axuser_0_axuser),
                   .int_rd_req_desc_2_axuser_1_axuser(int_rd_req_desc_2_axuser_1_axuser),
                   .int_rd_req_desc_2_axuser_2_axuser(int_rd_req_desc_2_axuser_2_axuser),
                   .int_rd_req_desc_2_axuser_3_axuser(int_rd_req_desc_2_axuser_3_axuser),
                   .int_rd_req_desc_2_axuser_4_axuser(int_rd_req_desc_2_axuser_4_axuser),
                   .int_rd_req_desc_2_axuser_5_axuser(int_rd_req_desc_2_axuser_5_axuser),
                   .int_rd_req_desc_2_axuser_6_axuser(int_rd_req_desc_2_axuser_6_axuser),
                   .int_rd_req_desc_2_axuser_7_axuser(int_rd_req_desc_2_axuser_7_axuser),
                   .int_rd_req_desc_2_axuser_8_axuser(int_rd_req_desc_2_axuser_8_axuser),
                   .int_rd_req_desc_2_axuser_9_axuser(int_rd_req_desc_2_axuser_9_axuser),
                   .int_rd_req_desc_2_axuser_10_axuser(int_rd_req_desc_2_axuser_10_axuser),
                   .int_rd_req_desc_2_axuser_11_axuser(int_rd_req_desc_2_axuser_11_axuser),
                   .int_rd_req_desc_2_axuser_12_axuser(int_rd_req_desc_2_axuser_12_axuser),
                   .int_rd_req_desc_2_axuser_13_axuser(int_rd_req_desc_2_axuser_13_axuser),
                   .int_rd_req_desc_2_axuser_14_axuser(int_rd_req_desc_2_axuser_14_axuser),
                   .int_rd_req_desc_2_axuser_15_axuser(int_rd_req_desc_2_axuser_15_axuser),
                   .int_wr_req_desc_2_txn_type_wr_strb(int_wr_req_desc_2_txn_type_wr_strb),
                   .int_wr_req_desc_2_size_txn_size(int_wr_req_desc_2_size_txn_size),
                   .int_wr_req_desc_2_data_offset_addr(int_wr_req_desc_2_data_offset_addr),
                   .int_wr_req_desc_2_axsize_axsize(int_wr_req_desc_2_axsize_axsize),
                   .int_wr_req_desc_2_attr_axsnoop(int_wr_req_desc_2_attr_axsnoop),
                   .int_wr_req_desc_2_attr_axdomain(int_wr_req_desc_2_attr_axdomain),
                   .int_wr_req_desc_2_attr_axbar(int_wr_req_desc_2_attr_axbar),
                   .int_wr_req_desc_2_attr_awunique(int_wr_req_desc_2_attr_awunique),
                   .int_wr_req_desc_2_attr_axregion(int_wr_req_desc_2_attr_axregion),
                   .int_wr_req_desc_2_attr_axqos(int_wr_req_desc_2_attr_axqos),
                   .int_wr_req_desc_2_attr_axprot(int_wr_req_desc_2_attr_axprot),
                   .int_wr_req_desc_2_attr_axcache(int_wr_req_desc_2_attr_axcache),
                   .int_wr_req_desc_2_attr_axlock(int_wr_req_desc_2_attr_axlock),
                   .int_wr_req_desc_2_attr_axburst(int_wr_req_desc_2_attr_axburst),
                   .int_wr_req_desc_2_axaddr_0_addr(int_wr_req_desc_2_axaddr_0_addr),
                   .int_wr_req_desc_2_axaddr_1_addr(int_wr_req_desc_2_axaddr_1_addr),
                   .int_wr_req_desc_2_axaddr_2_addr(int_wr_req_desc_2_axaddr_2_addr),
                   .int_wr_req_desc_2_axaddr_3_addr(int_wr_req_desc_2_axaddr_3_addr),
                   .int_wr_req_desc_2_axid_0_axid(int_wr_req_desc_2_axid_0_axid),
                   .int_wr_req_desc_2_axid_1_axid(int_wr_req_desc_2_axid_1_axid),
                   .int_wr_req_desc_2_axid_2_axid(int_wr_req_desc_2_axid_2_axid),
                   .int_wr_req_desc_2_axid_3_axid(int_wr_req_desc_2_axid_3_axid),
                   .int_wr_req_desc_2_axuser_0_axuser(int_wr_req_desc_2_axuser_0_axuser),
                   .int_wr_req_desc_2_axuser_1_axuser(int_wr_req_desc_2_axuser_1_axuser),
                   .int_wr_req_desc_2_axuser_2_axuser(int_wr_req_desc_2_axuser_2_axuser),
                   .int_wr_req_desc_2_axuser_3_axuser(int_wr_req_desc_2_axuser_3_axuser),
                   .int_wr_req_desc_2_axuser_4_axuser(int_wr_req_desc_2_axuser_4_axuser),
                   .int_wr_req_desc_2_axuser_5_axuser(int_wr_req_desc_2_axuser_5_axuser),
                   .int_wr_req_desc_2_axuser_6_axuser(int_wr_req_desc_2_axuser_6_axuser),
                   .int_wr_req_desc_2_axuser_7_axuser(int_wr_req_desc_2_axuser_7_axuser),
                   .int_wr_req_desc_2_axuser_8_axuser(int_wr_req_desc_2_axuser_8_axuser),
                   .int_wr_req_desc_2_axuser_9_axuser(int_wr_req_desc_2_axuser_9_axuser),
                   .int_wr_req_desc_2_axuser_10_axuser(int_wr_req_desc_2_axuser_10_axuser),
                   .int_wr_req_desc_2_axuser_11_axuser(int_wr_req_desc_2_axuser_11_axuser),
                   .int_wr_req_desc_2_axuser_12_axuser(int_wr_req_desc_2_axuser_12_axuser),
                   .int_wr_req_desc_2_axuser_13_axuser(int_wr_req_desc_2_axuser_13_axuser),
                   .int_wr_req_desc_2_axuser_14_axuser(int_wr_req_desc_2_axuser_14_axuser),
                   .int_wr_req_desc_2_axuser_15_axuser(int_wr_req_desc_2_axuser_15_axuser),
                   .int_wr_req_desc_2_wuser_0_wuser(int_wr_req_desc_2_wuser_0_wuser),
                   .int_wr_req_desc_2_wuser_1_wuser(int_wr_req_desc_2_wuser_1_wuser),
                   .int_wr_req_desc_2_wuser_2_wuser(int_wr_req_desc_2_wuser_2_wuser),
                   .int_wr_req_desc_2_wuser_3_wuser(int_wr_req_desc_2_wuser_3_wuser),
                   .int_wr_req_desc_2_wuser_4_wuser(int_wr_req_desc_2_wuser_4_wuser),
                   .int_wr_req_desc_2_wuser_5_wuser(int_wr_req_desc_2_wuser_5_wuser),
                   .int_wr_req_desc_2_wuser_6_wuser(int_wr_req_desc_2_wuser_6_wuser),
                   .int_wr_req_desc_2_wuser_7_wuser(int_wr_req_desc_2_wuser_7_wuser),
                   .int_wr_req_desc_2_wuser_8_wuser(int_wr_req_desc_2_wuser_8_wuser),
                   .int_wr_req_desc_2_wuser_9_wuser(int_wr_req_desc_2_wuser_9_wuser),
                   .int_wr_req_desc_2_wuser_10_wuser(int_wr_req_desc_2_wuser_10_wuser),
                   .int_wr_req_desc_2_wuser_11_wuser(int_wr_req_desc_2_wuser_11_wuser),
                   .int_wr_req_desc_2_wuser_12_wuser(int_wr_req_desc_2_wuser_12_wuser),
                   .int_wr_req_desc_2_wuser_13_wuser(int_wr_req_desc_2_wuser_13_wuser),
                   .int_wr_req_desc_2_wuser_14_wuser(int_wr_req_desc_2_wuser_14_wuser),
                   .int_wr_req_desc_2_wuser_15_wuser(int_wr_req_desc_2_wuser_15_wuser),
                   .int_sn_resp_desc_2_resp_resp(int_sn_resp_desc_2_resp_resp),
                   .int_rd_req_desc_3_size_txn_size(int_rd_req_desc_3_size_txn_size),
                   .int_rd_req_desc_3_axsize_axsize(int_rd_req_desc_3_axsize_axsize),
                   .int_rd_req_desc_3_attr_axsnoop(int_rd_req_desc_3_attr_axsnoop),
                   .int_rd_req_desc_3_attr_axdomain(int_rd_req_desc_3_attr_axdomain),
                   .int_rd_req_desc_3_attr_axbar(int_rd_req_desc_3_attr_axbar),
                   .int_rd_req_desc_3_attr_axregion(int_rd_req_desc_3_attr_axregion),
                   .int_rd_req_desc_3_attr_axqos(int_rd_req_desc_3_attr_axqos),
                   .int_rd_req_desc_3_attr_axprot(int_rd_req_desc_3_attr_axprot),
                   .int_rd_req_desc_3_attr_axcache(int_rd_req_desc_3_attr_axcache),
                   .int_rd_req_desc_3_attr_axlock(int_rd_req_desc_3_attr_axlock),
                   .int_rd_req_desc_3_attr_axburst(int_rd_req_desc_3_attr_axburst),
                   .int_rd_req_desc_3_axaddr_0_addr(int_rd_req_desc_3_axaddr_0_addr),
                   .int_rd_req_desc_3_axaddr_1_addr(int_rd_req_desc_3_axaddr_1_addr),
                   .int_rd_req_desc_3_axaddr_2_addr(int_rd_req_desc_3_axaddr_2_addr),
                   .int_rd_req_desc_3_axaddr_3_addr(int_rd_req_desc_3_axaddr_3_addr),
                   .int_rd_req_desc_3_axid_0_axid(int_rd_req_desc_3_axid_0_axid),
                   .int_rd_req_desc_3_axid_1_axid(int_rd_req_desc_3_axid_1_axid),
                   .int_rd_req_desc_3_axid_2_axid(int_rd_req_desc_3_axid_2_axid),
                   .int_rd_req_desc_3_axid_3_axid(int_rd_req_desc_3_axid_3_axid),
                   .int_rd_req_desc_3_axuser_0_axuser(int_rd_req_desc_3_axuser_0_axuser),
                   .int_rd_req_desc_3_axuser_1_axuser(int_rd_req_desc_3_axuser_1_axuser),
                   .int_rd_req_desc_3_axuser_2_axuser(int_rd_req_desc_3_axuser_2_axuser),
                   .int_rd_req_desc_3_axuser_3_axuser(int_rd_req_desc_3_axuser_3_axuser),
                   .int_rd_req_desc_3_axuser_4_axuser(int_rd_req_desc_3_axuser_4_axuser),
                   .int_rd_req_desc_3_axuser_5_axuser(int_rd_req_desc_3_axuser_5_axuser),
                   .int_rd_req_desc_3_axuser_6_axuser(int_rd_req_desc_3_axuser_6_axuser),
                   .int_rd_req_desc_3_axuser_7_axuser(int_rd_req_desc_3_axuser_7_axuser),
                   .int_rd_req_desc_3_axuser_8_axuser(int_rd_req_desc_3_axuser_8_axuser),
                   .int_rd_req_desc_3_axuser_9_axuser(int_rd_req_desc_3_axuser_9_axuser),
                   .int_rd_req_desc_3_axuser_10_axuser(int_rd_req_desc_3_axuser_10_axuser),
                   .int_rd_req_desc_3_axuser_11_axuser(int_rd_req_desc_3_axuser_11_axuser),
                   .int_rd_req_desc_3_axuser_12_axuser(int_rd_req_desc_3_axuser_12_axuser),
                   .int_rd_req_desc_3_axuser_13_axuser(int_rd_req_desc_3_axuser_13_axuser),
                   .int_rd_req_desc_3_axuser_14_axuser(int_rd_req_desc_3_axuser_14_axuser),
                   .int_rd_req_desc_3_axuser_15_axuser(int_rd_req_desc_3_axuser_15_axuser),
                   .int_wr_req_desc_3_txn_type_wr_strb(int_wr_req_desc_3_txn_type_wr_strb),
                   .int_wr_req_desc_3_size_txn_size(int_wr_req_desc_3_size_txn_size),
                   .int_wr_req_desc_3_data_offset_addr(int_wr_req_desc_3_data_offset_addr),
                   .int_wr_req_desc_3_axsize_axsize(int_wr_req_desc_3_axsize_axsize),
                   .int_wr_req_desc_3_attr_axsnoop(int_wr_req_desc_3_attr_axsnoop),
                   .int_wr_req_desc_3_attr_axdomain(int_wr_req_desc_3_attr_axdomain),
                   .int_wr_req_desc_3_attr_axbar(int_wr_req_desc_3_attr_axbar),
                   .int_wr_req_desc_3_attr_awunique(int_wr_req_desc_3_attr_awunique),
                   .int_wr_req_desc_3_attr_axregion(int_wr_req_desc_3_attr_axregion),
                   .int_wr_req_desc_3_attr_axqos(int_wr_req_desc_3_attr_axqos),
                   .int_wr_req_desc_3_attr_axprot(int_wr_req_desc_3_attr_axprot),
                   .int_wr_req_desc_3_attr_axcache(int_wr_req_desc_3_attr_axcache),
                   .int_wr_req_desc_3_attr_axlock(int_wr_req_desc_3_attr_axlock),
                   .int_wr_req_desc_3_attr_axburst(int_wr_req_desc_3_attr_axburst),
                   .int_wr_req_desc_3_axaddr_0_addr(int_wr_req_desc_3_axaddr_0_addr),
                   .int_wr_req_desc_3_axaddr_1_addr(int_wr_req_desc_3_axaddr_1_addr),
                   .int_wr_req_desc_3_axaddr_2_addr(int_wr_req_desc_3_axaddr_2_addr),
                   .int_wr_req_desc_3_axaddr_3_addr(int_wr_req_desc_3_axaddr_3_addr),
                   .int_wr_req_desc_3_axid_0_axid(int_wr_req_desc_3_axid_0_axid),
                   .int_wr_req_desc_3_axid_1_axid(int_wr_req_desc_3_axid_1_axid),
                   .int_wr_req_desc_3_axid_2_axid(int_wr_req_desc_3_axid_2_axid),
                   .int_wr_req_desc_3_axid_3_axid(int_wr_req_desc_3_axid_3_axid),
                   .int_wr_req_desc_3_axuser_0_axuser(int_wr_req_desc_3_axuser_0_axuser),
                   .int_wr_req_desc_3_axuser_1_axuser(int_wr_req_desc_3_axuser_1_axuser),
                   .int_wr_req_desc_3_axuser_2_axuser(int_wr_req_desc_3_axuser_2_axuser),
                   .int_wr_req_desc_3_axuser_3_axuser(int_wr_req_desc_3_axuser_3_axuser),
                   .int_wr_req_desc_3_axuser_4_axuser(int_wr_req_desc_3_axuser_4_axuser),
                   .int_wr_req_desc_3_axuser_5_axuser(int_wr_req_desc_3_axuser_5_axuser),
                   .int_wr_req_desc_3_axuser_6_axuser(int_wr_req_desc_3_axuser_6_axuser),
                   .int_wr_req_desc_3_axuser_7_axuser(int_wr_req_desc_3_axuser_7_axuser),
                   .int_wr_req_desc_3_axuser_8_axuser(int_wr_req_desc_3_axuser_8_axuser),
                   .int_wr_req_desc_3_axuser_9_axuser(int_wr_req_desc_3_axuser_9_axuser),
                   .int_wr_req_desc_3_axuser_10_axuser(int_wr_req_desc_3_axuser_10_axuser),
                   .int_wr_req_desc_3_axuser_11_axuser(int_wr_req_desc_3_axuser_11_axuser),
                   .int_wr_req_desc_3_axuser_12_axuser(int_wr_req_desc_3_axuser_12_axuser),
                   .int_wr_req_desc_3_axuser_13_axuser(int_wr_req_desc_3_axuser_13_axuser),
                   .int_wr_req_desc_3_axuser_14_axuser(int_wr_req_desc_3_axuser_14_axuser),
                   .int_wr_req_desc_3_axuser_15_axuser(int_wr_req_desc_3_axuser_15_axuser),
                   .int_wr_req_desc_3_wuser_0_wuser(int_wr_req_desc_3_wuser_0_wuser),
                   .int_wr_req_desc_3_wuser_1_wuser(int_wr_req_desc_3_wuser_1_wuser),
                   .int_wr_req_desc_3_wuser_2_wuser(int_wr_req_desc_3_wuser_2_wuser),
                   .int_wr_req_desc_3_wuser_3_wuser(int_wr_req_desc_3_wuser_3_wuser),
                   .int_wr_req_desc_3_wuser_4_wuser(int_wr_req_desc_3_wuser_4_wuser),
                   .int_wr_req_desc_3_wuser_5_wuser(int_wr_req_desc_3_wuser_5_wuser),
                   .int_wr_req_desc_3_wuser_6_wuser(int_wr_req_desc_3_wuser_6_wuser),
                   .int_wr_req_desc_3_wuser_7_wuser(int_wr_req_desc_3_wuser_7_wuser),
                   .int_wr_req_desc_3_wuser_8_wuser(int_wr_req_desc_3_wuser_8_wuser),
                   .int_wr_req_desc_3_wuser_9_wuser(int_wr_req_desc_3_wuser_9_wuser),
                   .int_wr_req_desc_3_wuser_10_wuser(int_wr_req_desc_3_wuser_10_wuser),
                   .int_wr_req_desc_3_wuser_11_wuser(int_wr_req_desc_3_wuser_11_wuser),
                   .int_wr_req_desc_3_wuser_12_wuser(int_wr_req_desc_3_wuser_12_wuser),
                   .int_wr_req_desc_3_wuser_13_wuser(int_wr_req_desc_3_wuser_13_wuser),
                   .int_wr_req_desc_3_wuser_14_wuser(int_wr_req_desc_3_wuser_14_wuser),
                   .int_wr_req_desc_3_wuser_15_wuser(int_wr_req_desc_3_wuser_15_wuser),
                   .int_sn_resp_desc_3_resp_resp(int_sn_resp_desc_3_resp_resp),
                   .int_rd_req_desc_4_size_txn_size(int_rd_req_desc_4_size_txn_size),
                   .int_rd_req_desc_4_axsize_axsize(int_rd_req_desc_4_axsize_axsize),
                   .int_rd_req_desc_4_attr_axsnoop(int_rd_req_desc_4_attr_axsnoop),
                   .int_rd_req_desc_4_attr_axdomain(int_rd_req_desc_4_attr_axdomain),
                   .int_rd_req_desc_4_attr_axbar(int_rd_req_desc_4_attr_axbar),
                   .int_rd_req_desc_4_attr_axregion(int_rd_req_desc_4_attr_axregion),
                   .int_rd_req_desc_4_attr_axqos(int_rd_req_desc_4_attr_axqos),
                   .int_rd_req_desc_4_attr_axprot(int_rd_req_desc_4_attr_axprot),
                   .int_rd_req_desc_4_attr_axcache(int_rd_req_desc_4_attr_axcache),
                   .int_rd_req_desc_4_attr_axlock(int_rd_req_desc_4_attr_axlock),
                   .int_rd_req_desc_4_attr_axburst(int_rd_req_desc_4_attr_axburst),
                   .int_rd_req_desc_4_axaddr_0_addr(int_rd_req_desc_4_axaddr_0_addr),
                   .int_rd_req_desc_4_axaddr_1_addr(int_rd_req_desc_4_axaddr_1_addr),
                   .int_rd_req_desc_4_axaddr_2_addr(int_rd_req_desc_4_axaddr_2_addr),
                   .int_rd_req_desc_4_axaddr_3_addr(int_rd_req_desc_4_axaddr_3_addr),
                   .int_rd_req_desc_4_axid_0_axid(int_rd_req_desc_4_axid_0_axid),
                   .int_rd_req_desc_4_axid_1_axid(int_rd_req_desc_4_axid_1_axid),
                   .int_rd_req_desc_4_axid_2_axid(int_rd_req_desc_4_axid_2_axid),
                   .int_rd_req_desc_4_axid_3_axid(int_rd_req_desc_4_axid_3_axid),
                   .int_rd_req_desc_4_axuser_0_axuser(int_rd_req_desc_4_axuser_0_axuser),
                   .int_rd_req_desc_4_axuser_1_axuser(int_rd_req_desc_4_axuser_1_axuser),
                   .int_rd_req_desc_4_axuser_2_axuser(int_rd_req_desc_4_axuser_2_axuser),
                   .int_rd_req_desc_4_axuser_3_axuser(int_rd_req_desc_4_axuser_3_axuser),
                   .int_rd_req_desc_4_axuser_4_axuser(int_rd_req_desc_4_axuser_4_axuser),
                   .int_rd_req_desc_4_axuser_5_axuser(int_rd_req_desc_4_axuser_5_axuser),
                   .int_rd_req_desc_4_axuser_6_axuser(int_rd_req_desc_4_axuser_6_axuser),
                   .int_rd_req_desc_4_axuser_7_axuser(int_rd_req_desc_4_axuser_7_axuser),
                   .int_rd_req_desc_4_axuser_8_axuser(int_rd_req_desc_4_axuser_8_axuser),
                   .int_rd_req_desc_4_axuser_9_axuser(int_rd_req_desc_4_axuser_9_axuser),
                   .int_rd_req_desc_4_axuser_10_axuser(int_rd_req_desc_4_axuser_10_axuser),
                   .int_rd_req_desc_4_axuser_11_axuser(int_rd_req_desc_4_axuser_11_axuser),
                   .int_rd_req_desc_4_axuser_12_axuser(int_rd_req_desc_4_axuser_12_axuser),
                   .int_rd_req_desc_4_axuser_13_axuser(int_rd_req_desc_4_axuser_13_axuser),
                   .int_rd_req_desc_4_axuser_14_axuser(int_rd_req_desc_4_axuser_14_axuser),
                   .int_rd_req_desc_4_axuser_15_axuser(int_rd_req_desc_4_axuser_15_axuser),
                   .int_wr_req_desc_4_txn_type_wr_strb(int_wr_req_desc_4_txn_type_wr_strb),
                   .int_wr_req_desc_4_size_txn_size(int_wr_req_desc_4_size_txn_size),
                   .int_wr_req_desc_4_data_offset_addr(int_wr_req_desc_4_data_offset_addr),
                   .int_wr_req_desc_4_axsize_axsize(int_wr_req_desc_4_axsize_axsize),
                   .int_wr_req_desc_4_attr_axsnoop(int_wr_req_desc_4_attr_axsnoop),
                   .int_wr_req_desc_4_attr_axdomain(int_wr_req_desc_4_attr_axdomain),
                   .int_wr_req_desc_4_attr_axbar(int_wr_req_desc_4_attr_axbar),
                   .int_wr_req_desc_4_attr_awunique(int_wr_req_desc_4_attr_awunique),
                   .int_wr_req_desc_4_attr_axregion(int_wr_req_desc_4_attr_axregion),
                   .int_wr_req_desc_4_attr_axqos(int_wr_req_desc_4_attr_axqos),
                   .int_wr_req_desc_4_attr_axprot(int_wr_req_desc_4_attr_axprot),
                   .int_wr_req_desc_4_attr_axcache(int_wr_req_desc_4_attr_axcache),
                   .int_wr_req_desc_4_attr_axlock(int_wr_req_desc_4_attr_axlock),
                   .int_wr_req_desc_4_attr_axburst(int_wr_req_desc_4_attr_axburst),
                   .int_wr_req_desc_4_axaddr_0_addr(int_wr_req_desc_4_axaddr_0_addr),
                   .int_wr_req_desc_4_axaddr_1_addr(int_wr_req_desc_4_axaddr_1_addr),
                   .int_wr_req_desc_4_axaddr_2_addr(int_wr_req_desc_4_axaddr_2_addr),
                   .int_wr_req_desc_4_axaddr_3_addr(int_wr_req_desc_4_axaddr_3_addr),
                   .int_wr_req_desc_4_axid_0_axid(int_wr_req_desc_4_axid_0_axid),
                   .int_wr_req_desc_4_axid_1_axid(int_wr_req_desc_4_axid_1_axid),
                   .int_wr_req_desc_4_axid_2_axid(int_wr_req_desc_4_axid_2_axid),
                   .int_wr_req_desc_4_axid_3_axid(int_wr_req_desc_4_axid_3_axid),
                   .int_wr_req_desc_4_axuser_0_axuser(int_wr_req_desc_4_axuser_0_axuser),
                   .int_wr_req_desc_4_axuser_1_axuser(int_wr_req_desc_4_axuser_1_axuser),
                   .int_wr_req_desc_4_axuser_2_axuser(int_wr_req_desc_4_axuser_2_axuser),
                   .int_wr_req_desc_4_axuser_3_axuser(int_wr_req_desc_4_axuser_3_axuser),
                   .int_wr_req_desc_4_axuser_4_axuser(int_wr_req_desc_4_axuser_4_axuser),
                   .int_wr_req_desc_4_axuser_5_axuser(int_wr_req_desc_4_axuser_5_axuser),
                   .int_wr_req_desc_4_axuser_6_axuser(int_wr_req_desc_4_axuser_6_axuser),
                   .int_wr_req_desc_4_axuser_7_axuser(int_wr_req_desc_4_axuser_7_axuser),
                   .int_wr_req_desc_4_axuser_8_axuser(int_wr_req_desc_4_axuser_8_axuser),
                   .int_wr_req_desc_4_axuser_9_axuser(int_wr_req_desc_4_axuser_9_axuser),
                   .int_wr_req_desc_4_axuser_10_axuser(int_wr_req_desc_4_axuser_10_axuser),
                   .int_wr_req_desc_4_axuser_11_axuser(int_wr_req_desc_4_axuser_11_axuser),
                   .int_wr_req_desc_4_axuser_12_axuser(int_wr_req_desc_4_axuser_12_axuser),
                   .int_wr_req_desc_4_axuser_13_axuser(int_wr_req_desc_4_axuser_13_axuser),
                   .int_wr_req_desc_4_axuser_14_axuser(int_wr_req_desc_4_axuser_14_axuser),
                   .int_wr_req_desc_4_axuser_15_axuser(int_wr_req_desc_4_axuser_15_axuser),
                   .int_wr_req_desc_4_wuser_0_wuser(int_wr_req_desc_4_wuser_0_wuser),
                   .int_wr_req_desc_4_wuser_1_wuser(int_wr_req_desc_4_wuser_1_wuser),
                   .int_wr_req_desc_4_wuser_2_wuser(int_wr_req_desc_4_wuser_2_wuser),
                   .int_wr_req_desc_4_wuser_3_wuser(int_wr_req_desc_4_wuser_3_wuser),
                   .int_wr_req_desc_4_wuser_4_wuser(int_wr_req_desc_4_wuser_4_wuser),
                   .int_wr_req_desc_4_wuser_5_wuser(int_wr_req_desc_4_wuser_5_wuser),
                   .int_wr_req_desc_4_wuser_6_wuser(int_wr_req_desc_4_wuser_6_wuser),
                   .int_wr_req_desc_4_wuser_7_wuser(int_wr_req_desc_4_wuser_7_wuser),
                   .int_wr_req_desc_4_wuser_8_wuser(int_wr_req_desc_4_wuser_8_wuser),
                   .int_wr_req_desc_4_wuser_9_wuser(int_wr_req_desc_4_wuser_9_wuser),
                   .int_wr_req_desc_4_wuser_10_wuser(int_wr_req_desc_4_wuser_10_wuser),
                   .int_wr_req_desc_4_wuser_11_wuser(int_wr_req_desc_4_wuser_11_wuser),
                   .int_wr_req_desc_4_wuser_12_wuser(int_wr_req_desc_4_wuser_12_wuser),
                   .int_wr_req_desc_4_wuser_13_wuser(int_wr_req_desc_4_wuser_13_wuser),
                   .int_wr_req_desc_4_wuser_14_wuser(int_wr_req_desc_4_wuser_14_wuser),
                   .int_wr_req_desc_4_wuser_15_wuser(int_wr_req_desc_4_wuser_15_wuser),
                   .int_sn_resp_desc_4_resp_resp(int_sn_resp_desc_4_resp_resp),
                   .int_rd_req_desc_5_size_txn_size(int_rd_req_desc_5_size_txn_size),
                   .int_rd_req_desc_5_axsize_axsize(int_rd_req_desc_5_axsize_axsize),
                   .int_rd_req_desc_5_attr_axsnoop(int_rd_req_desc_5_attr_axsnoop),
                   .int_rd_req_desc_5_attr_axdomain(int_rd_req_desc_5_attr_axdomain),
                   .int_rd_req_desc_5_attr_axbar(int_rd_req_desc_5_attr_axbar),
                   .int_rd_req_desc_5_attr_axregion(int_rd_req_desc_5_attr_axregion),
                   .int_rd_req_desc_5_attr_axqos(int_rd_req_desc_5_attr_axqos),
                   .int_rd_req_desc_5_attr_axprot(int_rd_req_desc_5_attr_axprot),
                   .int_rd_req_desc_5_attr_axcache(int_rd_req_desc_5_attr_axcache),
                   .int_rd_req_desc_5_attr_axlock(int_rd_req_desc_5_attr_axlock),
                   .int_rd_req_desc_5_attr_axburst(int_rd_req_desc_5_attr_axburst),
                   .int_rd_req_desc_5_axaddr_0_addr(int_rd_req_desc_5_axaddr_0_addr),
                   .int_rd_req_desc_5_axaddr_1_addr(int_rd_req_desc_5_axaddr_1_addr),
                   .int_rd_req_desc_5_axaddr_2_addr(int_rd_req_desc_5_axaddr_2_addr),
                   .int_rd_req_desc_5_axaddr_3_addr(int_rd_req_desc_5_axaddr_3_addr),
                   .int_rd_req_desc_5_axid_0_axid(int_rd_req_desc_5_axid_0_axid),
                   .int_rd_req_desc_5_axid_1_axid(int_rd_req_desc_5_axid_1_axid),
                   .int_rd_req_desc_5_axid_2_axid(int_rd_req_desc_5_axid_2_axid),
                   .int_rd_req_desc_5_axid_3_axid(int_rd_req_desc_5_axid_3_axid),
                   .int_rd_req_desc_5_axuser_0_axuser(int_rd_req_desc_5_axuser_0_axuser),
                   .int_rd_req_desc_5_axuser_1_axuser(int_rd_req_desc_5_axuser_1_axuser),
                   .int_rd_req_desc_5_axuser_2_axuser(int_rd_req_desc_5_axuser_2_axuser),
                   .int_rd_req_desc_5_axuser_3_axuser(int_rd_req_desc_5_axuser_3_axuser),
                   .int_rd_req_desc_5_axuser_4_axuser(int_rd_req_desc_5_axuser_4_axuser),
                   .int_rd_req_desc_5_axuser_5_axuser(int_rd_req_desc_5_axuser_5_axuser),
                   .int_rd_req_desc_5_axuser_6_axuser(int_rd_req_desc_5_axuser_6_axuser),
                   .int_rd_req_desc_5_axuser_7_axuser(int_rd_req_desc_5_axuser_7_axuser),
                   .int_rd_req_desc_5_axuser_8_axuser(int_rd_req_desc_5_axuser_8_axuser),
                   .int_rd_req_desc_5_axuser_9_axuser(int_rd_req_desc_5_axuser_9_axuser),
                   .int_rd_req_desc_5_axuser_10_axuser(int_rd_req_desc_5_axuser_10_axuser),
                   .int_rd_req_desc_5_axuser_11_axuser(int_rd_req_desc_5_axuser_11_axuser),
                   .int_rd_req_desc_5_axuser_12_axuser(int_rd_req_desc_5_axuser_12_axuser),
                   .int_rd_req_desc_5_axuser_13_axuser(int_rd_req_desc_5_axuser_13_axuser),
                   .int_rd_req_desc_5_axuser_14_axuser(int_rd_req_desc_5_axuser_14_axuser),
                   .int_rd_req_desc_5_axuser_15_axuser(int_rd_req_desc_5_axuser_15_axuser),
                   .int_wr_req_desc_5_txn_type_wr_strb(int_wr_req_desc_5_txn_type_wr_strb),
                   .int_wr_req_desc_5_size_txn_size(int_wr_req_desc_5_size_txn_size),
                   .int_wr_req_desc_5_data_offset_addr(int_wr_req_desc_5_data_offset_addr),
                   .int_wr_req_desc_5_axsize_axsize(int_wr_req_desc_5_axsize_axsize),
                   .int_wr_req_desc_5_attr_axsnoop(int_wr_req_desc_5_attr_axsnoop),
                   .int_wr_req_desc_5_attr_axdomain(int_wr_req_desc_5_attr_axdomain),
                   .int_wr_req_desc_5_attr_axbar(int_wr_req_desc_5_attr_axbar),
                   .int_wr_req_desc_5_attr_awunique(int_wr_req_desc_5_attr_awunique),
                   .int_wr_req_desc_5_attr_axregion(int_wr_req_desc_5_attr_axregion),
                   .int_wr_req_desc_5_attr_axqos(int_wr_req_desc_5_attr_axqos),
                   .int_wr_req_desc_5_attr_axprot(int_wr_req_desc_5_attr_axprot),
                   .int_wr_req_desc_5_attr_axcache(int_wr_req_desc_5_attr_axcache),
                   .int_wr_req_desc_5_attr_axlock(int_wr_req_desc_5_attr_axlock),
                   .int_wr_req_desc_5_attr_axburst(int_wr_req_desc_5_attr_axburst),
                   .int_wr_req_desc_5_axaddr_0_addr(int_wr_req_desc_5_axaddr_0_addr),
                   .int_wr_req_desc_5_axaddr_1_addr(int_wr_req_desc_5_axaddr_1_addr),
                   .int_wr_req_desc_5_axaddr_2_addr(int_wr_req_desc_5_axaddr_2_addr),
                   .int_wr_req_desc_5_axaddr_3_addr(int_wr_req_desc_5_axaddr_3_addr),
                   .int_wr_req_desc_5_axid_0_axid(int_wr_req_desc_5_axid_0_axid),
                   .int_wr_req_desc_5_axid_1_axid(int_wr_req_desc_5_axid_1_axid),
                   .int_wr_req_desc_5_axid_2_axid(int_wr_req_desc_5_axid_2_axid),
                   .int_wr_req_desc_5_axid_3_axid(int_wr_req_desc_5_axid_3_axid),
                   .int_wr_req_desc_5_axuser_0_axuser(int_wr_req_desc_5_axuser_0_axuser),
                   .int_wr_req_desc_5_axuser_1_axuser(int_wr_req_desc_5_axuser_1_axuser),
                   .int_wr_req_desc_5_axuser_2_axuser(int_wr_req_desc_5_axuser_2_axuser),
                   .int_wr_req_desc_5_axuser_3_axuser(int_wr_req_desc_5_axuser_3_axuser),
                   .int_wr_req_desc_5_axuser_4_axuser(int_wr_req_desc_5_axuser_4_axuser),
                   .int_wr_req_desc_5_axuser_5_axuser(int_wr_req_desc_5_axuser_5_axuser),
                   .int_wr_req_desc_5_axuser_6_axuser(int_wr_req_desc_5_axuser_6_axuser),
                   .int_wr_req_desc_5_axuser_7_axuser(int_wr_req_desc_5_axuser_7_axuser),
                   .int_wr_req_desc_5_axuser_8_axuser(int_wr_req_desc_5_axuser_8_axuser),
                   .int_wr_req_desc_5_axuser_9_axuser(int_wr_req_desc_5_axuser_9_axuser),
                   .int_wr_req_desc_5_axuser_10_axuser(int_wr_req_desc_5_axuser_10_axuser),
                   .int_wr_req_desc_5_axuser_11_axuser(int_wr_req_desc_5_axuser_11_axuser),
                   .int_wr_req_desc_5_axuser_12_axuser(int_wr_req_desc_5_axuser_12_axuser),
                   .int_wr_req_desc_5_axuser_13_axuser(int_wr_req_desc_5_axuser_13_axuser),
                   .int_wr_req_desc_5_axuser_14_axuser(int_wr_req_desc_5_axuser_14_axuser),
                   .int_wr_req_desc_5_axuser_15_axuser(int_wr_req_desc_5_axuser_15_axuser),
                   .int_wr_req_desc_5_wuser_0_wuser(int_wr_req_desc_5_wuser_0_wuser),
                   .int_wr_req_desc_5_wuser_1_wuser(int_wr_req_desc_5_wuser_1_wuser),
                   .int_wr_req_desc_5_wuser_2_wuser(int_wr_req_desc_5_wuser_2_wuser),
                   .int_wr_req_desc_5_wuser_3_wuser(int_wr_req_desc_5_wuser_3_wuser),
                   .int_wr_req_desc_5_wuser_4_wuser(int_wr_req_desc_5_wuser_4_wuser),
                   .int_wr_req_desc_5_wuser_5_wuser(int_wr_req_desc_5_wuser_5_wuser),
                   .int_wr_req_desc_5_wuser_6_wuser(int_wr_req_desc_5_wuser_6_wuser),
                   .int_wr_req_desc_5_wuser_7_wuser(int_wr_req_desc_5_wuser_7_wuser),
                   .int_wr_req_desc_5_wuser_8_wuser(int_wr_req_desc_5_wuser_8_wuser),
                   .int_wr_req_desc_5_wuser_9_wuser(int_wr_req_desc_5_wuser_9_wuser),
                   .int_wr_req_desc_5_wuser_10_wuser(int_wr_req_desc_5_wuser_10_wuser),
                   .int_wr_req_desc_5_wuser_11_wuser(int_wr_req_desc_5_wuser_11_wuser),
                   .int_wr_req_desc_5_wuser_12_wuser(int_wr_req_desc_5_wuser_12_wuser),
                   .int_wr_req_desc_5_wuser_13_wuser(int_wr_req_desc_5_wuser_13_wuser),
                   .int_wr_req_desc_5_wuser_14_wuser(int_wr_req_desc_5_wuser_14_wuser),
                   .int_wr_req_desc_5_wuser_15_wuser(int_wr_req_desc_5_wuser_15_wuser),
                   .int_sn_resp_desc_5_resp_resp(int_sn_resp_desc_5_resp_resp),
                   .int_rd_req_desc_6_size_txn_size(int_rd_req_desc_6_size_txn_size),
                   .int_rd_req_desc_6_axsize_axsize(int_rd_req_desc_6_axsize_axsize),
                   .int_rd_req_desc_6_attr_axsnoop(int_rd_req_desc_6_attr_axsnoop),
                   .int_rd_req_desc_6_attr_axdomain(int_rd_req_desc_6_attr_axdomain),
                   .int_rd_req_desc_6_attr_axbar(int_rd_req_desc_6_attr_axbar),
                   .int_rd_req_desc_6_attr_axregion(int_rd_req_desc_6_attr_axregion),
                   .int_rd_req_desc_6_attr_axqos(int_rd_req_desc_6_attr_axqos),
                   .int_rd_req_desc_6_attr_axprot(int_rd_req_desc_6_attr_axprot),
                   .int_rd_req_desc_6_attr_axcache(int_rd_req_desc_6_attr_axcache),
                   .int_rd_req_desc_6_attr_axlock(int_rd_req_desc_6_attr_axlock),
                   .int_rd_req_desc_6_attr_axburst(int_rd_req_desc_6_attr_axburst),
                   .int_rd_req_desc_6_axaddr_0_addr(int_rd_req_desc_6_axaddr_0_addr),
                   .int_rd_req_desc_6_axaddr_1_addr(int_rd_req_desc_6_axaddr_1_addr),
                   .int_rd_req_desc_6_axaddr_2_addr(int_rd_req_desc_6_axaddr_2_addr),
                   .int_rd_req_desc_6_axaddr_3_addr(int_rd_req_desc_6_axaddr_3_addr),
                   .int_rd_req_desc_6_axid_0_axid(int_rd_req_desc_6_axid_0_axid),
                   .int_rd_req_desc_6_axid_1_axid(int_rd_req_desc_6_axid_1_axid),
                   .int_rd_req_desc_6_axid_2_axid(int_rd_req_desc_6_axid_2_axid),
                   .int_rd_req_desc_6_axid_3_axid(int_rd_req_desc_6_axid_3_axid),
                   .int_rd_req_desc_6_axuser_0_axuser(int_rd_req_desc_6_axuser_0_axuser),
                   .int_rd_req_desc_6_axuser_1_axuser(int_rd_req_desc_6_axuser_1_axuser),
                   .int_rd_req_desc_6_axuser_2_axuser(int_rd_req_desc_6_axuser_2_axuser),
                   .int_rd_req_desc_6_axuser_3_axuser(int_rd_req_desc_6_axuser_3_axuser),
                   .int_rd_req_desc_6_axuser_4_axuser(int_rd_req_desc_6_axuser_4_axuser),
                   .int_rd_req_desc_6_axuser_5_axuser(int_rd_req_desc_6_axuser_5_axuser),
                   .int_rd_req_desc_6_axuser_6_axuser(int_rd_req_desc_6_axuser_6_axuser),
                   .int_rd_req_desc_6_axuser_7_axuser(int_rd_req_desc_6_axuser_7_axuser),
                   .int_rd_req_desc_6_axuser_8_axuser(int_rd_req_desc_6_axuser_8_axuser),
                   .int_rd_req_desc_6_axuser_9_axuser(int_rd_req_desc_6_axuser_9_axuser),
                   .int_rd_req_desc_6_axuser_10_axuser(int_rd_req_desc_6_axuser_10_axuser),
                   .int_rd_req_desc_6_axuser_11_axuser(int_rd_req_desc_6_axuser_11_axuser),
                   .int_rd_req_desc_6_axuser_12_axuser(int_rd_req_desc_6_axuser_12_axuser),
                   .int_rd_req_desc_6_axuser_13_axuser(int_rd_req_desc_6_axuser_13_axuser),
                   .int_rd_req_desc_6_axuser_14_axuser(int_rd_req_desc_6_axuser_14_axuser),
                   .int_rd_req_desc_6_axuser_15_axuser(int_rd_req_desc_6_axuser_15_axuser),
                   .int_wr_req_desc_6_txn_type_wr_strb(int_wr_req_desc_6_txn_type_wr_strb),
                   .int_wr_req_desc_6_size_txn_size(int_wr_req_desc_6_size_txn_size),
                   .int_wr_req_desc_6_data_offset_addr(int_wr_req_desc_6_data_offset_addr),
                   .int_wr_req_desc_6_axsize_axsize(int_wr_req_desc_6_axsize_axsize),
                   .int_wr_req_desc_6_attr_axsnoop(int_wr_req_desc_6_attr_axsnoop),
                   .int_wr_req_desc_6_attr_axdomain(int_wr_req_desc_6_attr_axdomain),
                   .int_wr_req_desc_6_attr_axbar(int_wr_req_desc_6_attr_axbar),
                   .int_wr_req_desc_6_attr_awunique(int_wr_req_desc_6_attr_awunique),
                   .int_wr_req_desc_6_attr_axregion(int_wr_req_desc_6_attr_axregion),
                   .int_wr_req_desc_6_attr_axqos(int_wr_req_desc_6_attr_axqos),
                   .int_wr_req_desc_6_attr_axprot(int_wr_req_desc_6_attr_axprot),
                   .int_wr_req_desc_6_attr_axcache(int_wr_req_desc_6_attr_axcache),
                   .int_wr_req_desc_6_attr_axlock(int_wr_req_desc_6_attr_axlock),
                   .int_wr_req_desc_6_attr_axburst(int_wr_req_desc_6_attr_axburst),
                   .int_wr_req_desc_6_axaddr_0_addr(int_wr_req_desc_6_axaddr_0_addr),
                   .int_wr_req_desc_6_axaddr_1_addr(int_wr_req_desc_6_axaddr_1_addr),
                   .int_wr_req_desc_6_axaddr_2_addr(int_wr_req_desc_6_axaddr_2_addr),
                   .int_wr_req_desc_6_axaddr_3_addr(int_wr_req_desc_6_axaddr_3_addr),
                   .int_wr_req_desc_6_axid_0_axid(int_wr_req_desc_6_axid_0_axid),
                   .int_wr_req_desc_6_axid_1_axid(int_wr_req_desc_6_axid_1_axid),
                   .int_wr_req_desc_6_axid_2_axid(int_wr_req_desc_6_axid_2_axid),
                   .int_wr_req_desc_6_axid_3_axid(int_wr_req_desc_6_axid_3_axid),
                   .int_wr_req_desc_6_axuser_0_axuser(int_wr_req_desc_6_axuser_0_axuser),
                   .int_wr_req_desc_6_axuser_1_axuser(int_wr_req_desc_6_axuser_1_axuser),
                   .int_wr_req_desc_6_axuser_2_axuser(int_wr_req_desc_6_axuser_2_axuser),
                   .int_wr_req_desc_6_axuser_3_axuser(int_wr_req_desc_6_axuser_3_axuser),
                   .int_wr_req_desc_6_axuser_4_axuser(int_wr_req_desc_6_axuser_4_axuser),
                   .int_wr_req_desc_6_axuser_5_axuser(int_wr_req_desc_6_axuser_5_axuser),
                   .int_wr_req_desc_6_axuser_6_axuser(int_wr_req_desc_6_axuser_6_axuser),
                   .int_wr_req_desc_6_axuser_7_axuser(int_wr_req_desc_6_axuser_7_axuser),
                   .int_wr_req_desc_6_axuser_8_axuser(int_wr_req_desc_6_axuser_8_axuser),
                   .int_wr_req_desc_6_axuser_9_axuser(int_wr_req_desc_6_axuser_9_axuser),
                   .int_wr_req_desc_6_axuser_10_axuser(int_wr_req_desc_6_axuser_10_axuser),
                   .int_wr_req_desc_6_axuser_11_axuser(int_wr_req_desc_6_axuser_11_axuser),
                   .int_wr_req_desc_6_axuser_12_axuser(int_wr_req_desc_6_axuser_12_axuser),
                   .int_wr_req_desc_6_axuser_13_axuser(int_wr_req_desc_6_axuser_13_axuser),
                   .int_wr_req_desc_6_axuser_14_axuser(int_wr_req_desc_6_axuser_14_axuser),
                   .int_wr_req_desc_6_axuser_15_axuser(int_wr_req_desc_6_axuser_15_axuser),
                   .int_wr_req_desc_6_wuser_0_wuser(int_wr_req_desc_6_wuser_0_wuser),
                   .int_wr_req_desc_6_wuser_1_wuser(int_wr_req_desc_6_wuser_1_wuser),
                   .int_wr_req_desc_6_wuser_2_wuser(int_wr_req_desc_6_wuser_2_wuser),
                   .int_wr_req_desc_6_wuser_3_wuser(int_wr_req_desc_6_wuser_3_wuser),
                   .int_wr_req_desc_6_wuser_4_wuser(int_wr_req_desc_6_wuser_4_wuser),
                   .int_wr_req_desc_6_wuser_5_wuser(int_wr_req_desc_6_wuser_5_wuser),
                   .int_wr_req_desc_6_wuser_6_wuser(int_wr_req_desc_6_wuser_6_wuser),
                   .int_wr_req_desc_6_wuser_7_wuser(int_wr_req_desc_6_wuser_7_wuser),
                   .int_wr_req_desc_6_wuser_8_wuser(int_wr_req_desc_6_wuser_8_wuser),
                   .int_wr_req_desc_6_wuser_9_wuser(int_wr_req_desc_6_wuser_9_wuser),
                   .int_wr_req_desc_6_wuser_10_wuser(int_wr_req_desc_6_wuser_10_wuser),
                   .int_wr_req_desc_6_wuser_11_wuser(int_wr_req_desc_6_wuser_11_wuser),
                   .int_wr_req_desc_6_wuser_12_wuser(int_wr_req_desc_6_wuser_12_wuser),
                   .int_wr_req_desc_6_wuser_13_wuser(int_wr_req_desc_6_wuser_13_wuser),
                   .int_wr_req_desc_6_wuser_14_wuser(int_wr_req_desc_6_wuser_14_wuser),
                   .int_wr_req_desc_6_wuser_15_wuser(int_wr_req_desc_6_wuser_15_wuser),
                   .int_sn_resp_desc_6_resp_resp(int_sn_resp_desc_6_resp_resp),
                   .int_rd_req_desc_7_size_txn_size(int_rd_req_desc_7_size_txn_size),
                   .int_rd_req_desc_7_axsize_axsize(int_rd_req_desc_7_axsize_axsize),
                   .int_rd_req_desc_7_attr_axsnoop(int_rd_req_desc_7_attr_axsnoop),
                   .int_rd_req_desc_7_attr_axdomain(int_rd_req_desc_7_attr_axdomain),
                   .int_rd_req_desc_7_attr_axbar(int_rd_req_desc_7_attr_axbar),
                   .int_rd_req_desc_7_attr_axregion(int_rd_req_desc_7_attr_axregion),
                   .int_rd_req_desc_7_attr_axqos(int_rd_req_desc_7_attr_axqos),
                   .int_rd_req_desc_7_attr_axprot(int_rd_req_desc_7_attr_axprot),
                   .int_rd_req_desc_7_attr_axcache(int_rd_req_desc_7_attr_axcache),
                   .int_rd_req_desc_7_attr_axlock(int_rd_req_desc_7_attr_axlock),
                   .int_rd_req_desc_7_attr_axburst(int_rd_req_desc_7_attr_axburst),
                   .int_rd_req_desc_7_axaddr_0_addr(int_rd_req_desc_7_axaddr_0_addr),
                   .int_rd_req_desc_7_axaddr_1_addr(int_rd_req_desc_7_axaddr_1_addr),
                   .int_rd_req_desc_7_axaddr_2_addr(int_rd_req_desc_7_axaddr_2_addr),
                   .int_rd_req_desc_7_axaddr_3_addr(int_rd_req_desc_7_axaddr_3_addr),
                   .int_rd_req_desc_7_axid_0_axid(int_rd_req_desc_7_axid_0_axid),
                   .int_rd_req_desc_7_axid_1_axid(int_rd_req_desc_7_axid_1_axid),
                   .int_rd_req_desc_7_axid_2_axid(int_rd_req_desc_7_axid_2_axid),
                   .int_rd_req_desc_7_axid_3_axid(int_rd_req_desc_7_axid_3_axid),
                   .int_rd_req_desc_7_axuser_0_axuser(int_rd_req_desc_7_axuser_0_axuser),
                   .int_rd_req_desc_7_axuser_1_axuser(int_rd_req_desc_7_axuser_1_axuser),
                   .int_rd_req_desc_7_axuser_2_axuser(int_rd_req_desc_7_axuser_2_axuser),
                   .int_rd_req_desc_7_axuser_3_axuser(int_rd_req_desc_7_axuser_3_axuser),
                   .int_rd_req_desc_7_axuser_4_axuser(int_rd_req_desc_7_axuser_4_axuser),
                   .int_rd_req_desc_7_axuser_5_axuser(int_rd_req_desc_7_axuser_5_axuser),
                   .int_rd_req_desc_7_axuser_6_axuser(int_rd_req_desc_7_axuser_6_axuser),
                   .int_rd_req_desc_7_axuser_7_axuser(int_rd_req_desc_7_axuser_7_axuser),
                   .int_rd_req_desc_7_axuser_8_axuser(int_rd_req_desc_7_axuser_8_axuser),
                   .int_rd_req_desc_7_axuser_9_axuser(int_rd_req_desc_7_axuser_9_axuser),
                   .int_rd_req_desc_7_axuser_10_axuser(int_rd_req_desc_7_axuser_10_axuser),
                   .int_rd_req_desc_7_axuser_11_axuser(int_rd_req_desc_7_axuser_11_axuser),
                   .int_rd_req_desc_7_axuser_12_axuser(int_rd_req_desc_7_axuser_12_axuser),
                   .int_rd_req_desc_7_axuser_13_axuser(int_rd_req_desc_7_axuser_13_axuser),
                   .int_rd_req_desc_7_axuser_14_axuser(int_rd_req_desc_7_axuser_14_axuser),
                   .int_rd_req_desc_7_axuser_15_axuser(int_rd_req_desc_7_axuser_15_axuser),
                   .int_wr_req_desc_7_txn_type_wr_strb(int_wr_req_desc_7_txn_type_wr_strb),
                   .int_wr_req_desc_7_size_txn_size(int_wr_req_desc_7_size_txn_size),
                   .int_wr_req_desc_7_data_offset_addr(int_wr_req_desc_7_data_offset_addr),
                   .int_wr_req_desc_7_axsize_axsize(int_wr_req_desc_7_axsize_axsize),
                   .int_wr_req_desc_7_attr_axsnoop(int_wr_req_desc_7_attr_axsnoop),
                   .int_wr_req_desc_7_attr_axdomain(int_wr_req_desc_7_attr_axdomain),
                   .int_wr_req_desc_7_attr_axbar(int_wr_req_desc_7_attr_axbar),
                   .int_wr_req_desc_7_attr_awunique(int_wr_req_desc_7_attr_awunique),
                   .int_wr_req_desc_7_attr_axregion(int_wr_req_desc_7_attr_axregion),
                   .int_wr_req_desc_7_attr_axqos(int_wr_req_desc_7_attr_axqos),
                   .int_wr_req_desc_7_attr_axprot(int_wr_req_desc_7_attr_axprot),
                   .int_wr_req_desc_7_attr_axcache(int_wr_req_desc_7_attr_axcache),
                   .int_wr_req_desc_7_attr_axlock(int_wr_req_desc_7_attr_axlock),
                   .int_wr_req_desc_7_attr_axburst(int_wr_req_desc_7_attr_axburst),
                   .int_wr_req_desc_7_axaddr_0_addr(int_wr_req_desc_7_axaddr_0_addr),
                   .int_wr_req_desc_7_axaddr_1_addr(int_wr_req_desc_7_axaddr_1_addr),
                   .int_wr_req_desc_7_axaddr_2_addr(int_wr_req_desc_7_axaddr_2_addr),
                   .int_wr_req_desc_7_axaddr_3_addr(int_wr_req_desc_7_axaddr_3_addr),
                   .int_wr_req_desc_7_axid_0_axid(int_wr_req_desc_7_axid_0_axid),
                   .int_wr_req_desc_7_axid_1_axid(int_wr_req_desc_7_axid_1_axid),
                   .int_wr_req_desc_7_axid_2_axid(int_wr_req_desc_7_axid_2_axid),
                   .int_wr_req_desc_7_axid_3_axid(int_wr_req_desc_7_axid_3_axid),
                   .int_wr_req_desc_7_axuser_0_axuser(int_wr_req_desc_7_axuser_0_axuser),
                   .int_wr_req_desc_7_axuser_1_axuser(int_wr_req_desc_7_axuser_1_axuser),
                   .int_wr_req_desc_7_axuser_2_axuser(int_wr_req_desc_7_axuser_2_axuser),
                   .int_wr_req_desc_7_axuser_3_axuser(int_wr_req_desc_7_axuser_3_axuser),
                   .int_wr_req_desc_7_axuser_4_axuser(int_wr_req_desc_7_axuser_4_axuser),
                   .int_wr_req_desc_7_axuser_5_axuser(int_wr_req_desc_7_axuser_5_axuser),
                   .int_wr_req_desc_7_axuser_6_axuser(int_wr_req_desc_7_axuser_6_axuser),
                   .int_wr_req_desc_7_axuser_7_axuser(int_wr_req_desc_7_axuser_7_axuser),
                   .int_wr_req_desc_7_axuser_8_axuser(int_wr_req_desc_7_axuser_8_axuser),
                   .int_wr_req_desc_7_axuser_9_axuser(int_wr_req_desc_7_axuser_9_axuser),
                   .int_wr_req_desc_7_axuser_10_axuser(int_wr_req_desc_7_axuser_10_axuser),
                   .int_wr_req_desc_7_axuser_11_axuser(int_wr_req_desc_7_axuser_11_axuser),
                   .int_wr_req_desc_7_axuser_12_axuser(int_wr_req_desc_7_axuser_12_axuser),
                   .int_wr_req_desc_7_axuser_13_axuser(int_wr_req_desc_7_axuser_13_axuser),
                   .int_wr_req_desc_7_axuser_14_axuser(int_wr_req_desc_7_axuser_14_axuser),
                   .int_wr_req_desc_7_axuser_15_axuser(int_wr_req_desc_7_axuser_15_axuser),
                   .int_wr_req_desc_7_wuser_0_wuser(int_wr_req_desc_7_wuser_0_wuser),
                   .int_wr_req_desc_7_wuser_1_wuser(int_wr_req_desc_7_wuser_1_wuser),
                   .int_wr_req_desc_7_wuser_2_wuser(int_wr_req_desc_7_wuser_2_wuser),
                   .int_wr_req_desc_7_wuser_3_wuser(int_wr_req_desc_7_wuser_3_wuser),
                   .int_wr_req_desc_7_wuser_4_wuser(int_wr_req_desc_7_wuser_4_wuser),
                   .int_wr_req_desc_7_wuser_5_wuser(int_wr_req_desc_7_wuser_5_wuser),
                   .int_wr_req_desc_7_wuser_6_wuser(int_wr_req_desc_7_wuser_6_wuser),
                   .int_wr_req_desc_7_wuser_7_wuser(int_wr_req_desc_7_wuser_7_wuser),
                   .int_wr_req_desc_7_wuser_8_wuser(int_wr_req_desc_7_wuser_8_wuser),
                   .int_wr_req_desc_7_wuser_9_wuser(int_wr_req_desc_7_wuser_9_wuser),
                   .int_wr_req_desc_7_wuser_10_wuser(int_wr_req_desc_7_wuser_10_wuser),
                   .int_wr_req_desc_7_wuser_11_wuser(int_wr_req_desc_7_wuser_11_wuser),
                   .int_wr_req_desc_7_wuser_12_wuser(int_wr_req_desc_7_wuser_12_wuser),
                   .int_wr_req_desc_7_wuser_13_wuser(int_wr_req_desc_7_wuser_13_wuser),
                   .int_wr_req_desc_7_wuser_14_wuser(int_wr_req_desc_7_wuser_14_wuser),
                   .int_wr_req_desc_7_wuser_15_wuser(int_wr_req_desc_7_wuser_15_wuser),
                   .int_sn_resp_desc_7_resp_resp(int_sn_resp_desc_7_resp_resp),
                   .int_rd_req_desc_8_size_txn_size(int_rd_req_desc_8_size_txn_size),
                   .int_rd_req_desc_8_axsize_axsize(int_rd_req_desc_8_axsize_axsize),
                   .int_rd_req_desc_8_attr_axsnoop(int_rd_req_desc_8_attr_axsnoop),
                   .int_rd_req_desc_8_attr_axdomain(int_rd_req_desc_8_attr_axdomain),
                   .int_rd_req_desc_8_attr_axbar(int_rd_req_desc_8_attr_axbar),
                   .int_rd_req_desc_8_attr_axregion(int_rd_req_desc_8_attr_axregion),
                   .int_rd_req_desc_8_attr_axqos(int_rd_req_desc_8_attr_axqos),
                   .int_rd_req_desc_8_attr_axprot(int_rd_req_desc_8_attr_axprot),
                   .int_rd_req_desc_8_attr_axcache(int_rd_req_desc_8_attr_axcache),
                   .int_rd_req_desc_8_attr_axlock(int_rd_req_desc_8_attr_axlock),
                   .int_rd_req_desc_8_attr_axburst(int_rd_req_desc_8_attr_axburst),
                   .int_rd_req_desc_8_axaddr_0_addr(int_rd_req_desc_8_axaddr_0_addr),
                   .int_rd_req_desc_8_axaddr_1_addr(int_rd_req_desc_8_axaddr_1_addr),
                   .int_rd_req_desc_8_axaddr_2_addr(int_rd_req_desc_8_axaddr_2_addr),
                   .int_rd_req_desc_8_axaddr_3_addr(int_rd_req_desc_8_axaddr_3_addr),
                   .int_rd_req_desc_8_axid_0_axid(int_rd_req_desc_8_axid_0_axid),
                   .int_rd_req_desc_8_axid_1_axid(int_rd_req_desc_8_axid_1_axid),
                   .int_rd_req_desc_8_axid_2_axid(int_rd_req_desc_8_axid_2_axid),
                   .int_rd_req_desc_8_axid_3_axid(int_rd_req_desc_8_axid_3_axid),
                   .int_rd_req_desc_8_axuser_0_axuser(int_rd_req_desc_8_axuser_0_axuser),
                   .int_rd_req_desc_8_axuser_1_axuser(int_rd_req_desc_8_axuser_1_axuser),
                   .int_rd_req_desc_8_axuser_2_axuser(int_rd_req_desc_8_axuser_2_axuser),
                   .int_rd_req_desc_8_axuser_3_axuser(int_rd_req_desc_8_axuser_3_axuser),
                   .int_rd_req_desc_8_axuser_4_axuser(int_rd_req_desc_8_axuser_4_axuser),
                   .int_rd_req_desc_8_axuser_5_axuser(int_rd_req_desc_8_axuser_5_axuser),
                   .int_rd_req_desc_8_axuser_6_axuser(int_rd_req_desc_8_axuser_6_axuser),
                   .int_rd_req_desc_8_axuser_7_axuser(int_rd_req_desc_8_axuser_7_axuser),
                   .int_rd_req_desc_8_axuser_8_axuser(int_rd_req_desc_8_axuser_8_axuser),
                   .int_rd_req_desc_8_axuser_9_axuser(int_rd_req_desc_8_axuser_9_axuser),
                   .int_rd_req_desc_8_axuser_10_axuser(int_rd_req_desc_8_axuser_10_axuser),
                   .int_rd_req_desc_8_axuser_11_axuser(int_rd_req_desc_8_axuser_11_axuser),
                   .int_rd_req_desc_8_axuser_12_axuser(int_rd_req_desc_8_axuser_12_axuser),
                   .int_rd_req_desc_8_axuser_13_axuser(int_rd_req_desc_8_axuser_13_axuser),
                   .int_rd_req_desc_8_axuser_14_axuser(int_rd_req_desc_8_axuser_14_axuser),
                   .int_rd_req_desc_8_axuser_15_axuser(int_rd_req_desc_8_axuser_15_axuser),
                   .int_wr_req_desc_8_txn_type_wr_strb(int_wr_req_desc_8_txn_type_wr_strb),
                   .int_wr_req_desc_8_size_txn_size(int_wr_req_desc_8_size_txn_size),
                   .int_wr_req_desc_8_data_offset_addr(int_wr_req_desc_8_data_offset_addr),
                   .int_wr_req_desc_8_axsize_axsize(int_wr_req_desc_8_axsize_axsize),
                   .int_wr_req_desc_8_attr_axsnoop(int_wr_req_desc_8_attr_axsnoop),
                   .int_wr_req_desc_8_attr_axdomain(int_wr_req_desc_8_attr_axdomain),
                   .int_wr_req_desc_8_attr_axbar(int_wr_req_desc_8_attr_axbar),
                   .int_wr_req_desc_8_attr_awunique(int_wr_req_desc_8_attr_awunique),
                   .int_wr_req_desc_8_attr_axregion(int_wr_req_desc_8_attr_axregion),
                   .int_wr_req_desc_8_attr_axqos(int_wr_req_desc_8_attr_axqos),
                   .int_wr_req_desc_8_attr_axprot(int_wr_req_desc_8_attr_axprot),
                   .int_wr_req_desc_8_attr_axcache(int_wr_req_desc_8_attr_axcache),
                   .int_wr_req_desc_8_attr_axlock(int_wr_req_desc_8_attr_axlock),
                   .int_wr_req_desc_8_attr_axburst(int_wr_req_desc_8_attr_axburst),
                   .int_wr_req_desc_8_axaddr_0_addr(int_wr_req_desc_8_axaddr_0_addr),
                   .int_wr_req_desc_8_axaddr_1_addr(int_wr_req_desc_8_axaddr_1_addr),
                   .int_wr_req_desc_8_axaddr_2_addr(int_wr_req_desc_8_axaddr_2_addr),
                   .int_wr_req_desc_8_axaddr_3_addr(int_wr_req_desc_8_axaddr_3_addr),
                   .int_wr_req_desc_8_axid_0_axid(int_wr_req_desc_8_axid_0_axid),
                   .int_wr_req_desc_8_axid_1_axid(int_wr_req_desc_8_axid_1_axid),
                   .int_wr_req_desc_8_axid_2_axid(int_wr_req_desc_8_axid_2_axid),
                   .int_wr_req_desc_8_axid_3_axid(int_wr_req_desc_8_axid_3_axid),
                   .int_wr_req_desc_8_axuser_0_axuser(int_wr_req_desc_8_axuser_0_axuser),
                   .int_wr_req_desc_8_axuser_1_axuser(int_wr_req_desc_8_axuser_1_axuser),
                   .int_wr_req_desc_8_axuser_2_axuser(int_wr_req_desc_8_axuser_2_axuser),
                   .int_wr_req_desc_8_axuser_3_axuser(int_wr_req_desc_8_axuser_3_axuser),
                   .int_wr_req_desc_8_axuser_4_axuser(int_wr_req_desc_8_axuser_4_axuser),
                   .int_wr_req_desc_8_axuser_5_axuser(int_wr_req_desc_8_axuser_5_axuser),
                   .int_wr_req_desc_8_axuser_6_axuser(int_wr_req_desc_8_axuser_6_axuser),
                   .int_wr_req_desc_8_axuser_7_axuser(int_wr_req_desc_8_axuser_7_axuser),
                   .int_wr_req_desc_8_axuser_8_axuser(int_wr_req_desc_8_axuser_8_axuser),
                   .int_wr_req_desc_8_axuser_9_axuser(int_wr_req_desc_8_axuser_9_axuser),
                   .int_wr_req_desc_8_axuser_10_axuser(int_wr_req_desc_8_axuser_10_axuser),
                   .int_wr_req_desc_8_axuser_11_axuser(int_wr_req_desc_8_axuser_11_axuser),
                   .int_wr_req_desc_8_axuser_12_axuser(int_wr_req_desc_8_axuser_12_axuser),
                   .int_wr_req_desc_8_axuser_13_axuser(int_wr_req_desc_8_axuser_13_axuser),
                   .int_wr_req_desc_8_axuser_14_axuser(int_wr_req_desc_8_axuser_14_axuser),
                   .int_wr_req_desc_8_axuser_15_axuser(int_wr_req_desc_8_axuser_15_axuser),
                   .int_wr_req_desc_8_wuser_0_wuser(int_wr_req_desc_8_wuser_0_wuser),
                   .int_wr_req_desc_8_wuser_1_wuser(int_wr_req_desc_8_wuser_1_wuser),
                   .int_wr_req_desc_8_wuser_2_wuser(int_wr_req_desc_8_wuser_2_wuser),
                   .int_wr_req_desc_8_wuser_3_wuser(int_wr_req_desc_8_wuser_3_wuser),
                   .int_wr_req_desc_8_wuser_4_wuser(int_wr_req_desc_8_wuser_4_wuser),
                   .int_wr_req_desc_8_wuser_5_wuser(int_wr_req_desc_8_wuser_5_wuser),
                   .int_wr_req_desc_8_wuser_6_wuser(int_wr_req_desc_8_wuser_6_wuser),
                   .int_wr_req_desc_8_wuser_7_wuser(int_wr_req_desc_8_wuser_7_wuser),
                   .int_wr_req_desc_8_wuser_8_wuser(int_wr_req_desc_8_wuser_8_wuser),
                   .int_wr_req_desc_8_wuser_9_wuser(int_wr_req_desc_8_wuser_9_wuser),
                   .int_wr_req_desc_8_wuser_10_wuser(int_wr_req_desc_8_wuser_10_wuser),
                   .int_wr_req_desc_8_wuser_11_wuser(int_wr_req_desc_8_wuser_11_wuser),
                   .int_wr_req_desc_8_wuser_12_wuser(int_wr_req_desc_8_wuser_12_wuser),
                   .int_wr_req_desc_8_wuser_13_wuser(int_wr_req_desc_8_wuser_13_wuser),
                   .int_wr_req_desc_8_wuser_14_wuser(int_wr_req_desc_8_wuser_14_wuser),
                   .int_wr_req_desc_8_wuser_15_wuser(int_wr_req_desc_8_wuser_15_wuser),
                   .int_sn_resp_desc_8_resp_resp(int_sn_resp_desc_8_resp_resp),
                   .int_rd_req_desc_9_size_txn_size(int_rd_req_desc_9_size_txn_size),
                   .int_rd_req_desc_9_axsize_axsize(int_rd_req_desc_9_axsize_axsize),
                   .int_rd_req_desc_9_attr_axsnoop(int_rd_req_desc_9_attr_axsnoop),
                   .int_rd_req_desc_9_attr_axdomain(int_rd_req_desc_9_attr_axdomain),
                   .int_rd_req_desc_9_attr_axbar(int_rd_req_desc_9_attr_axbar),
                   .int_rd_req_desc_9_attr_axregion(int_rd_req_desc_9_attr_axregion),
                   .int_rd_req_desc_9_attr_axqos(int_rd_req_desc_9_attr_axqos),
                   .int_rd_req_desc_9_attr_axprot(int_rd_req_desc_9_attr_axprot),
                   .int_rd_req_desc_9_attr_axcache(int_rd_req_desc_9_attr_axcache),
                   .int_rd_req_desc_9_attr_axlock(int_rd_req_desc_9_attr_axlock),
                   .int_rd_req_desc_9_attr_axburst(int_rd_req_desc_9_attr_axburst),
                   .int_rd_req_desc_9_axaddr_0_addr(int_rd_req_desc_9_axaddr_0_addr),
                   .int_rd_req_desc_9_axaddr_1_addr(int_rd_req_desc_9_axaddr_1_addr),
                   .int_rd_req_desc_9_axaddr_2_addr(int_rd_req_desc_9_axaddr_2_addr),
                   .int_rd_req_desc_9_axaddr_3_addr(int_rd_req_desc_9_axaddr_3_addr),
                   .int_rd_req_desc_9_axid_0_axid(int_rd_req_desc_9_axid_0_axid),
                   .int_rd_req_desc_9_axid_1_axid(int_rd_req_desc_9_axid_1_axid),
                   .int_rd_req_desc_9_axid_2_axid(int_rd_req_desc_9_axid_2_axid),
                   .int_rd_req_desc_9_axid_3_axid(int_rd_req_desc_9_axid_3_axid),
                   .int_rd_req_desc_9_axuser_0_axuser(int_rd_req_desc_9_axuser_0_axuser),
                   .int_rd_req_desc_9_axuser_1_axuser(int_rd_req_desc_9_axuser_1_axuser),
                   .int_rd_req_desc_9_axuser_2_axuser(int_rd_req_desc_9_axuser_2_axuser),
                   .int_rd_req_desc_9_axuser_3_axuser(int_rd_req_desc_9_axuser_3_axuser),
                   .int_rd_req_desc_9_axuser_4_axuser(int_rd_req_desc_9_axuser_4_axuser),
                   .int_rd_req_desc_9_axuser_5_axuser(int_rd_req_desc_9_axuser_5_axuser),
                   .int_rd_req_desc_9_axuser_6_axuser(int_rd_req_desc_9_axuser_6_axuser),
                   .int_rd_req_desc_9_axuser_7_axuser(int_rd_req_desc_9_axuser_7_axuser),
                   .int_rd_req_desc_9_axuser_8_axuser(int_rd_req_desc_9_axuser_8_axuser),
                   .int_rd_req_desc_9_axuser_9_axuser(int_rd_req_desc_9_axuser_9_axuser),
                   .int_rd_req_desc_9_axuser_10_axuser(int_rd_req_desc_9_axuser_10_axuser),
                   .int_rd_req_desc_9_axuser_11_axuser(int_rd_req_desc_9_axuser_11_axuser),
                   .int_rd_req_desc_9_axuser_12_axuser(int_rd_req_desc_9_axuser_12_axuser),
                   .int_rd_req_desc_9_axuser_13_axuser(int_rd_req_desc_9_axuser_13_axuser),
                   .int_rd_req_desc_9_axuser_14_axuser(int_rd_req_desc_9_axuser_14_axuser),
                   .int_rd_req_desc_9_axuser_15_axuser(int_rd_req_desc_9_axuser_15_axuser),
                   .int_wr_req_desc_9_txn_type_wr_strb(int_wr_req_desc_9_txn_type_wr_strb),
                   .int_wr_req_desc_9_size_txn_size(int_wr_req_desc_9_size_txn_size),
                   .int_wr_req_desc_9_data_offset_addr(int_wr_req_desc_9_data_offset_addr),
                   .int_wr_req_desc_9_axsize_axsize(int_wr_req_desc_9_axsize_axsize),
                   .int_wr_req_desc_9_attr_axsnoop(int_wr_req_desc_9_attr_axsnoop),
                   .int_wr_req_desc_9_attr_axdomain(int_wr_req_desc_9_attr_axdomain),
                   .int_wr_req_desc_9_attr_axbar(int_wr_req_desc_9_attr_axbar),
                   .int_wr_req_desc_9_attr_awunique(int_wr_req_desc_9_attr_awunique),
                   .int_wr_req_desc_9_attr_axregion(int_wr_req_desc_9_attr_axregion),
                   .int_wr_req_desc_9_attr_axqos(int_wr_req_desc_9_attr_axqos),
                   .int_wr_req_desc_9_attr_axprot(int_wr_req_desc_9_attr_axprot),
                   .int_wr_req_desc_9_attr_axcache(int_wr_req_desc_9_attr_axcache),
                   .int_wr_req_desc_9_attr_axlock(int_wr_req_desc_9_attr_axlock),
                   .int_wr_req_desc_9_attr_axburst(int_wr_req_desc_9_attr_axburst),
                   .int_wr_req_desc_9_axaddr_0_addr(int_wr_req_desc_9_axaddr_0_addr),
                   .int_wr_req_desc_9_axaddr_1_addr(int_wr_req_desc_9_axaddr_1_addr),
                   .int_wr_req_desc_9_axaddr_2_addr(int_wr_req_desc_9_axaddr_2_addr),
                   .int_wr_req_desc_9_axaddr_3_addr(int_wr_req_desc_9_axaddr_3_addr),
                   .int_wr_req_desc_9_axid_0_axid(int_wr_req_desc_9_axid_0_axid),
                   .int_wr_req_desc_9_axid_1_axid(int_wr_req_desc_9_axid_1_axid),
                   .int_wr_req_desc_9_axid_2_axid(int_wr_req_desc_9_axid_2_axid),
                   .int_wr_req_desc_9_axid_3_axid(int_wr_req_desc_9_axid_3_axid),
                   .int_wr_req_desc_9_axuser_0_axuser(int_wr_req_desc_9_axuser_0_axuser),
                   .int_wr_req_desc_9_axuser_1_axuser(int_wr_req_desc_9_axuser_1_axuser),
                   .int_wr_req_desc_9_axuser_2_axuser(int_wr_req_desc_9_axuser_2_axuser),
                   .int_wr_req_desc_9_axuser_3_axuser(int_wr_req_desc_9_axuser_3_axuser),
                   .int_wr_req_desc_9_axuser_4_axuser(int_wr_req_desc_9_axuser_4_axuser),
                   .int_wr_req_desc_9_axuser_5_axuser(int_wr_req_desc_9_axuser_5_axuser),
                   .int_wr_req_desc_9_axuser_6_axuser(int_wr_req_desc_9_axuser_6_axuser),
                   .int_wr_req_desc_9_axuser_7_axuser(int_wr_req_desc_9_axuser_7_axuser),
                   .int_wr_req_desc_9_axuser_8_axuser(int_wr_req_desc_9_axuser_8_axuser),
                   .int_wr_req_desc_9_axuser_9_axuser(int_wr_req_desc_9_axuser_9_axuser),
                   .int_wr_req_desc_9_axuser_10_axuser(int_wr_req_desc_9_axuser_10_axuser),
                   .int_wr_req_desc_9_axuser_11_axuser(int_wr_req_desc_9_axuser_11_axuser),
                   .int_wr_req_desc_9_axuser_12_axuser(int_wr_req_desc_9_axuser_12_axuser),
                   .int_wr_req_desc_9_axuser_13_axuser(int_wr_req_desc_9_axuser_13_axuser),
                   .int_wr_req_desc_9_axuser_14_axuser(int_wr_req_desc_9_axuser_14_axuser),
                   .int_wr_req_desc_9_axuser_15_axuser(int_wr_req_desc_9_axuser_15_axuser),
                   .int_wr_req_desc_9_wuser_0_wuser(int_wr_req_desc_9_wuser_0_wuser),
                   .int_wr_req_desc_9_wuser_1_wuser(int_wr_req_desc_9_wuser_1_wuser),
                   .int_wr_req_desc_9_wuser_2_wuser(int_wr_req_desc_9_wuser_2_wuser),
                   .int_wr_req_desc_9_wuser_3_wuser(int_wr_req_desc_9_wuser_3_wuser),
                   .int_wr_req_desc_9_wuser_4_wuser(int_wr_req_desc_9_wuser_4_wuser),
                   .int_wr_req_desc_9_wuser_5_wuser(int_wr_req_desc_9_wuser_5_wuser),
                   .int_wr_req_desc_9_wuser_6_wuser(int_wr_req_desc_9_wuser_6_wuser),
                   .int_wr_req_desc_9_wuser_7_wuser(int_wr_req_desc_9_wuser_7_wuser),
                   .int_wr_req_desc_9_wuser_8_wuser(int_wr_req_desc_9_wuser_8_wuser),
                   .int_wr_req_desc_9_wuser_9_wuser(int_wr_req_desc_9_wuser_9_wuser),
                   .int_wr_req_desc_9_wuser_10_wuser(int_wr_req_desc_9_wuser_10_wuser),
                   .int_wr_req_desc_9_wuser_11_wuser(int_wr_req_desc_9_wuser_11_wuser),
                   .int_wr_req_desc_9_wuser_12_wuser(int_wr_req_desc_9_wuser_12_wuser),
                   .int_wr_req_desc_9_wuser_13_wuser(int_wr_req_desc_9_wuser_13_wuser),
                   .int_wr_req_desc_9_wuser_14_wuser(int_wr_req_desc_9_wuser_14_wuser),
                   .int_wr_req_desc_9_wuser_15_wuser(int_wr_req_desc_9_wuser_15_wuser),
                   .int_sn_resp_desc_9_resp_resp(int_sn_resp_desc_9_resp_resp),
                   .int_rd_req_desc_a_size_txn_size(int_rd_req_desc_a_size_txn_size),
                   .int_rd_req_desc_a_axsize_axsize(int_rd_req_desc_a_axsize_axsize),
                   .int_rd_req_desc_a_attr_axsnoop(int_rd_req_desc_a_attr_axsnoop),
                   .int_rd_req_desc_a_attr_axdomain(int_rd_req_desc_a_attr_axdomain),
                   .int_rd_req_desc_a_attr_axbar(int_rd_req_desc_a_attr_axbar),
                   .int_rd_req_desc_a_attr_axregion(int_rd_req_desc_a_attr_axregion),
                   .int_rd_req_desc_a_attr_axqos(int_rd_req_desc_a_attr_axqos),
                   .int_rd_req_desc_a_attr_axprot(int_rd_req_desc_a_attr_axprot),
                   .int_rd_req_desc_a_attr_axcache(int_rd_req_desc_a_attr_axcache),
                   .int_rd_req_desc_a_attr_axlock(int_rd_req_desc_a_attr_axlock),
                   .int_rd_req_desc_a_attr_axburst(int_rd_req_desc_a_attr_axburst),
                   .int_rd_req_desc_a_axaddr_0_addr(int_rd_req_desc_a_axaddr_0_addr),
                   .int_rd_req_desc_a_axaddr_1_addr(int_rd_req_desc_a_axaddr_1_addr),
                   .int_rd_req_desc_a_axaddr_2_addr(int_rd_req_desc_a_axaddr_2_addr),
                   .int_rd_req_desc_a_axaddr_3_addr(int_rd_req_desc_a_axaddr_3_addr),
                   .int_rd_req_desc_a_axid_0_axid(int_rd_req_desc_a_axid_0_axid),
                   .int_rd_req_desc_a_axid_1_axid(int_rd_req_desc_a_axid_1_axid),
                   .int_rd_req_desc_a_axid_2_axid(int_rd_req_desc_a_axid_2_axid),
                   .int_rd_req_desc_a_axid_3_axid(int_rd_req_desc_a_axid_3_axid),
                   .int_rd_req_desc_a_axuser_0_axuser(int_rd_req_desc_a_axuser_0_axuser),
                   .int_rd_req_desc_a_axuser_1_axuser(int_rd_req_desc_a_axuser_1_axuser),
                   .int_rd_req_desc_a_axuser_2_axuser(int_rd_req_desc_a_axuser_2_axuser),
                   .int_rd_req_desc_a_axuser_3_axuser(int_rd_req_desc_a_axuser_3_axuser),
                   .int_rd_req_desc_a_axuser_4_axuser(int_rd_req_desc_a_axuser_4_axuser),
                   .int_rd_req_desc_a_axuser_5_axuser(int_rd_req_desc_a_axuser_5_axuser),
                   .int_rd_req_desc_a_axuser_6_axuser(int_rd_req_desc_a_axuser_6_axuser),
                   .int_rd_req_desc_a_axuser_7_axuser(int_rd_req_desc_a_axuser_7_axuser),
                   .int_rd_req_desc_a_axuser_8_axuser(int_rd_req_desc_a_axuser_8_axuser),
                   .int_rd_req_desc_a_axuser_9_axuser(int_rd_req_desc_a_axuser_9_axuser),
                   .int_rd_req_desc_a_axuser_10_axuser(int_rd_req_desc_a_axuser_10_axuser),
                   .int_rd_req_desc_a_axuser_11_axuser(int_rd_req_desc_a_axuser_11_axuser),
                   .int_rd_req_desc_a_axuser_12_axuser(int_rd_req_desc_a_axuser_12_axuser),
                   .int_rd_req_desc_a_axuser_13_axuser(int_rd_req_desc_a_axuser_13_axuser),
                   .int_rd_req_desc_a_axuser_14_axuser(int_rd_req_desc_a_axuser_14_axuser),
                   .int_rd_req_desc_a_axuser_15_axuser(int_rd_req_desc_a_axuser_15_axuser),
                   .int_wr_req_desc_a_txn_type_wr_strb(int_wr_req_desc_a_txn_type_wr_strb),
                   .int_wr_req_desc_a_size_txn_size(int_wr_req_desc_a_size_txn_size),
                   .int_wr_req_desc_a_data_offset_addr(int_wr_req_desc_a_data_offset_addr),
                   .int_wr_req_desc_a_axsize_axsize(int_wr_req_desc_a_axsize_axsize),
                   .int_wr_req_desc_a_attr_axsnoop(int_wr_req_desc_a_attr_axsnoop),
                   .int_wr_req_desc_a_attr_axdomain(int_wr_req_desc_a_attr_axdomain),
                   .int_wr_req_desc_a_attr_axbar(int_wr_req_desc_a_attr_axbar),
                   .int_wr_req_desc_a_attr_awunique(int_wr_req_desc_a_attr_awunique),
                   .int_wr_req_desc_a_attr_axregion(int_wr_req_desc_a_attr_axregion),
                   .int_wr_req_desc_a_attr_axqos(int_wr_req_desc_a_attr_axqos),
                   .int_wr_req_desc_a_attr_axprot(int_wr_req_desc_a_attr_axprot),
                   .int_wr_req_desc_a_attr_axcache(int_wr_req_desc_a_attr_axcache),
                   .int_wr_req_desc_a_attr_axlock(int_wr_req_desc_a_attr_axlock),
                   .int_wr_req_desc_a_attr_axburst(int_wr_req_desc_a_attr_axburst),
                   .int_wr_req_desc_a_axaddr_0_addr(int_wr_req_desc_a_axaddr_0_addr),
                   .int_wr_req_desc_a_axaddr_1_addr(int_wr_req_desc_a_axaddr_1_addr),
                   .int_wr_req_desc_a_axaddr_2_addr(int_wr_req_desc_a_axaddr_2_addr),
                   .int_wr_req_desc_a_axaddr_3_addr(int_wr_req_desc_a_axaddr_3_addr),
                   .int_wr_req_desc_a_axid_0_axid(int_wr_req_desc_a_axid_0_axid),
                   .int_wr_req_desc_a_axid_1_axid(int_wr_req_desc_a_axid_1_axid),
                   .int_wr_req_desc_a_axid_2_axid(int_wr_req_desc_a_axid_2_axid),
                   .int_wr_req_desc_a_axid_3_axid(int_wr_req_desc_a_axid_3_axid),
                   .int_wr_req_desc_a_axuser_0_axuser(int_wr_req_desc_a_axuser_0_axuser),
                   .int_wr_req_desc_a_axuser_1_axuser(int_wr_req_desc_a_axuser_1_axuser),
                   .int_wr_req_desc_a_axuser_2_axuser(int_wr_req_desc_a_axuser_2_axuser),
                   .int_wr_req_desc_a_axuser_3_axuser(int_wr_req_desc_a_axuser_3_axuser),
                   .int_wr_req_desc_a_axuser_4_axuser(int_wr_req_desc_a_axuser_4_axuser),
                   .int_wr_req_desc_a_axuser_5_axuser(int_wr_req_desc_a_axuser_5_axuser),
                   .int_wr_req_desc_a_axuser_6_axuser(int_wr_req_desc_a_axuser_6_axuser),
                   .int_wr_req_desc_a_axuser_7_axuser(int_wr_req_desc_a_axuser_7_axuser),
                   .int_wr_req_desc_a_axuser_8_axuser(int_wr_req_desc_a_axuser_8_axuser),
                   .int_wr_req_desc_a_axuser_9_axuser(int_wr_req_desc_a_axuser_9_axuser),
                   .int_wr_req_desc_a_axuser_10_axuser(int_wr_req_desc_a_axuser_10_axuser),
                   .int_wr_req_desc_a_axuser_11_axuser(int_wr_req_desc_a_axuser_11_axuser),
                   .int_wr_req_desc_a_axuser_12_axuser(int_wr_req_desc_a_axuser_12_axuser),
                   .int_wr_req_desc_a_axuser_13_axuser(int_wr_req_desc_a_axuser_13_axuser),
                   .int_wr_req_desc_a_axuser_14_axuser(int_wr_req_desc_a_axuser_14_axuser),
                   .int_wr_req_desc_a_axuser_15_axuser(int_wr_req_desc_a_axuser_15_axuser),
                   .int_wr_req_desc_a_wuser_0_wuser(int_wr_req_desc_a_wuser_0_wuser),
                   .int_wr_req_desc_a_wuser_1_wuser(int_wr_req_desc_a_wuser_1_wuser),
                   .int_wr_req_desc_a_wuser_2_wuser(int_wr_req_desc_a_wuser_2_wuser),
                   .int_wr_req_desc_a_wuser_3_wuser(int_wr_req_desc_a_wuser_3_wuser),
                   .int_wr_req_desc_a_wuser_4_wuser(int_wr_req_desc_a_wuser_4_wuser),
                   .int_wr_req_desc_a_wuser_5_wuser(int_wr_req_desc_a_wuser_5_wuser),
                   .int_wr_req_desc_a_wuser_6_wuser(int_wr_req_desc_a_wuser_6_wuser),
                   .int_wr_req_desc_a_wuser_7_wuser(int_wr_req_desc_a_wuser_7_wuser),
                   .int_wr_req_desc_a_wuser_8_wuser(int_wr_req_desc_a_wuser_8_wuser),
                   .int_wr_req_desc_a_wuser_9_wuser(int_wr_req_desc_a_wuser_9_wuser),
                   .int_wr_req_desc_a_wuser_10_wuser(int_wr_req_desc_a_wuser_10_wuser),
                   .int_wr_req_desc_a_wuser_11_wuser(int_wr_req_desc_a_wuser_11_wuser),
                   .int_wr_req_desc_a_wuser_12_wuser(int_wr_req_desc_a_wuser_12_wuser),
                   .int_wr_req_desc_a_wuser_13_wuser(int_wr_req_desc_a_wuser_13_wuser),
                   .int_wr_req_desc_a_wuser_14_wuser(int_wr_req_desc_a_wuser_14_wuser),
                   .int_wr_req_desc_a_wuser_15_wuser(int_wr_req_desc_a_wuser_15_wuser),
                   .int_sn_resp_desc_a_resp_resp(int_sn_resp_desc_a_resp_resp),
                   .int_rd_req_desc_b_size_txn_size(int_rd_req_desc_b_size_txn_size),
                   .int_rd_req_desc_b_axsize_axsize(int_rd_req_desc_b_axsize_axsize),
                   .int_rd_req_desc_b_attr_axsnoop(int_rd_req_desc_b_attr_axsnoop),
                   .int_rd_req_desc_b_attr_axdomain(int_rd_req_desc_b_attr_axdomain),
                   .int_rd_req_desc_b_attr_axbar(int_rd_req_desc_b_attr_axbar),
                   .int_rd_req_desc_b_attr_axregion(int_rd_req_desc_b_attr_axregion),
                   .int_rd_req_desc_b_attr_axqos(int_rd_req_desc_b_attr_axqos),
                   .int_rd_req_desc_b_attr_axprot(int_rd_req_desc_b_attr_axprot),
                   .int_rd_req_desc_b_attr_axcache(int_rd_req_desc_b_attr_axcache),
                   .int_rd_req_desc_b_attr_axlock(int_rd_req_desc_b_attr_axlock),
                   .int_rd_req_desc_b_attr_axburst(int_rd_req_desc_b_attr_axburst),
                   .int_rd_req_desc_b_axaddr_0_addr(int_rd_req_desc_b_axaddr_0_addr),
                   .int_rd_req_desc_b_axaddr_1_addr(int_rd_req_desc_b_axaddr_1_addr),
                   .int_rd_req_desc_b_axaddr_2_addr(int_rd_req_desc_b_axaddr_2_addr),
                   .int_rd_req_desc_b_axaddr_3_addr(int_rd_req_desc_b_axaddr_3_addr),
                   .int_rd_req_desc_b_axid_0_axid(int_rd_req_desc_b_axid_0_axid),
                   .int_rd_req_desc_b_axid_1_axid(int_rd_req_desc_b_axid_1_axid),
                   .int_rd_req_desc_b_axid_2_axid(int_rd_req_desc_b_axid_2_axid),
                   .int_rd_req_desc_b_axid_3_axid(int_rd_req_desc_b_axid_3_axid),
                   .int_rd_req_desc_b_axuser_0_axuser(int_rd_req_desc_b_axuser_0_axuser),
                   .int_rd_req_desc_b_axuser_1_axuser(int_rd_req_desc_b_axuser_1_axuser),
                   .int_rd_req_desc_b_axuser_2_axuser(int_rd_req_desc_b_axuser_2_axuser),
                   .int_rd_req_desc_b_axuser_3_axuser(int_rd_req_desc_b_axuser_3_axuser),
                   .int_rd_req_desc_b_axuser_4_axuser(int_rd_req_desc_b_axuser_4_axuser),
                   .int_rd_req_desc_b_axuser_5_axuser(int_rd_req_desc_b_axuser_5_axuser),
                   .int_rd_req_desc_b_axuser_6_axuser(int_rd_req_desc_b_axuser_6_axuser),
                   .int_rd_req_desc_b_axuser_7_axuser(int_rd_req_desc_b_axuser_7_axuser),
                   .int_rd_req_desc_b_axuser_8_axuser(int_rd_req_desc_b_axuser_8_axuser),
                   .int_rd_req_desc_b_axuser_9_axuser(int_rd_req_desc_b_axuser_9_axuser),
                   .int_rd_req_desc_b_axuser_10_axuser(int_rd_req_desc_b_axuser_10_axuser),
                   .int_rd_req_desc_b_axuser_11_axuser(int_rd_req_desc_b_axuser_11_axuser),
                   .int_rd_req_desc_b_axuser_12_axuser(int_rd_req_desc_b_axuser_12_axuser),
                   .int_rd_req_desc_b_axuser_13_axuser(int_rd_req_desc_b_axuser_13_axuser),
                   .int_rd_req_desc_b_axuser_14_axuser(int_rd_req_desc_b_axuser_14_axuser),
                   .int_rd_req_desc_b_axuser_15_axuser(int_rd_req_desc_b_axuser_15_axuser),
                   .int_wr_req_desc_b_txn_type_wr_strb(int_wr_req_desc_b_txn_type_wr_strb),
                   .int_wr_req_desc_b_size_txn_size(int_wr_req_desc_b_size_txn_size),
                   .int_wr_req_desc_b_data_offset_addr(int_wr_req_desc_b_data_offset_addr),
                   .int_wr_req_desc_b_axsize_axsize(int_wr_req_desc_b_axsize_axsize),
                   .int_wr_req_desc_b_attr_axsnoop(int_wr_req_desc_b_attr_axsnoop),
                   .int_wr_req_desc_b_attr_axdomain(int_wr_req_desc_b_attr_axdomain),
                   .int_wr_req_desc_b_attr_axbar(int_wr_req_desc_b_attr_axbar),
                   .int_wr_req_desc_b_attr_awunique(int_wr_req_desc_b_attr_awunique),
                   .int_wr_req_desc_b_attr_axregion(int_wr_req_desc_b_attr_axregion),
                   .int_wr_req_desc_b_attr_axqos(int_wr_req_desc_b_attr_axqos),
                   .int_wr_req_desc_b_attr_axprot(int_wr_req_desc_b_attr_axprot),
                   .int_wr_req_desc_b_attr_axcache(int_wr_req_desc_b_attr_axcache),
                   .int_wr_req_desc_b_attr_axlock(int_wr_req_desc_b_attr_axlock),
                   .int_wr_req_desc_b_attr_axburst(int_wr_req_desc_b_attr_axburst),
                   .int_wr_req_desc_b_axaddr_0_addr(int_wr_req_desc_b_axaddr_0_addr),
                   .int_wr_req_desc_b_axaddr_1_addr(int_wr_req_desc_b_axaddr_1_addr),
                   .int_wr_req_desc_b_axaddr_2_addr(int_wr_req_desc_b_axaddr_2_addr),
                   .int_wr_req_desc_b_axaddr_3_addr(int_wr_req_desc_b_axaddr_3_addr),
                   .int_wr_req_desc_b_axid_0_axid(int_wr_req_desc_b_axid_0_axid),
                   .int_wr_req_desc_b_axid_1_axid(int_wr_req_desc_b_axid_1_axid),
                   .int_wr_req_desc_b_axid_2_axid(int_wr_req_desc_b_axid_2_axid),
                   .int_wr_req_desc_b_axid_3_axid(int_wr_req_desc_b_axid_3_axid),
                   .int_wr_req_desc_b_axuser_0_axuser(int_wr_req_desc_b_axuser_0_axuser),
                   .int_wr_req_desc_b_axuser_1_axuser(int_wr_req_desc_b_axuser_1_axuser),
                   .int_wr_req_desc_b_axuser_2_axuser(int_wr_req_desc_b_axuser_2_axuser),
                   .int_wr_req_desc_b_axuser_3_axuser(int_wr_req_desc_b_axuser_3_axuser),
                   .int_wr_req_desc_b_axuser_4_axuser(int_wr_req_desc_b_axuser_4_axuser),
                   .int_wr_req_desc_b_axuser_5_axuser(int_wr_req_desc_b_axuser_5_axuser),
                   .int_wr_req_desc_b_axuser_6_axuser(int_wr_req_desc_b_axuser_6_axuser),
                   .int_wr_req_desc_b_axuser_7_axuser(int_wr_req_desc_b_axuser_7_axuser),
                   .int_wr_req_desc_b_axuser_8_axuser(int_wr_req_desc_b_axuser_8_axuser),
                   .int_wr_req_desc_b_axuser_9_axuser(int_wr_req_desc_b_axuser_9_axuser),
                   .int_wr_req_desc_b_axuser_10_axuser(int_wr_req_desc_b_axuser_10_axuser),
                   .int_wr_req_desc_b_axuser_11_axuser(int_wr_req_desc_b_axuser_11_axuser),
                   .int_wr_req_desc_b_axuser_12_axuser(int_wr_req_desc_b_axuser_12_axuser),
                   .int_wr_req_desc_b_axuser_13_axuser(int_wr_req_desc_b_axuser_13_axuser),
                   .int_wr_req_desc_b_axuser_14_axuser(int_wr_req_desc_b_axuser_14_axuser),
                   .int_wr_req_desc_b_axuser_15_axuser(int_wr_req_desc_b_axuser_15_axuser),
                   .int_wr_req_desc_b_wuser_0_wuser(int_wr_req_desc_b_wuser_0_wuser),
                   .int_wr_req_desc_b_wuser_1_wuser(int_wr_req_desc_b_wuser_1_wuser),
                   .int_wr_req_desc_b_wuser_2_wuser(int_wr_req_desc_b_wuser_2_wuser),
                   .int_wr_req_desc_b_wuser_3_wuser(int_wr_req_desc_b_wuser_3_wuser),
                   .int_wr_req_desc_b_wuser_4_wuser(int_wr_req_desc_b_wuser_4_wuser),
                   .int_wr_req_desc_b_wuser_5_wuser(int_wr_req_desc_b_wuser_5_wuser),
                   .int_wr_req_desc_b_wuser_6_wuser(int_wr_req_desc_b_wuser_6_wuser),
                   .int_wr_req_desc_b_wuser_7_wuser(int_wr_req_desc_b_wuser_7_wuser),
                   .int_wr_req_desc_b_wuser_8_wuser(int_wr_req_desc_b_wuser_8_wuser),
                   .int_wr_req_desc_b_wuser_9_wuser(int_wr_req_desc_b_wuser_9_wuser),
                   .int_wr_req_desc_b_wuser_10_wuser(int_wr_req_desc_b_wuser_10_wuser),
                   .int_wr_req_desc_b_wuser_11_wuser(int_wr_req_desc_b_wuser_11_wuser),
                   .int_wr_req_desc_b_wuser_12_wuser(int_wr_req_desc_b_wuser_12_wuser),
                   .int_wr_req_desc_b_wuser_13_wuser(int_wr_req_desc_b_wuser_13_wuser),
                   .int_wr_req_desc_b_wuser_14_wuser(int_wr_req_desc_b_wuser_14_wuser),
                   .int_wr_req_desc_b_wuser_15_wuser(int_wr_req_desc_b_wuser_15_wuser),
                   .int_sn_resp_desc_b_resp_resp(int_sn_resp_desc_b_resp_resp),
                   .int_rd_req_desc_c_size_txn_size(int_rd_req_desc_c_size_txn_size),
                   .int_rd_req_desc_c_axsize_axsize(int_rd_req_desc_c_axsize_axsize),
                   .int_rd_req_desc_c_attr_axsnoop(int_rd_req_desc_c_attr_axsnoop),
                   .int_rd_req_desc_c_attr_axdomain(int_rd_req_desc_c_attr_axdomain),
                   .int_rd_req_desc_c_attr_axbar(int_rd_req_desc_c_attr_axbar),
                   .int_rd_req_desc_c_attr_axregion(int_rd_req_desc_c_attr_axregion),
                   .int_rd_req_desc_c_attr_axqos(int_rd_req_desc_c_attr_axqos),
                   .int_rd_req_desc_c_attr_axprot(int_rd_req_desc_c_attr_axprot),
                   .int_rd_req_desc_c_attr_axcache(int_rd_req_desc_c_attr_axcache),
                   .int_rd_req_desc_c_attr_axlock(int_rd_req_desc_c_attr_axlock),
                   .int_rd_req_desc_c_attr_axburst(int_rd_req_desc_c_attr_axburst),
                   .int_rd_req_desc_c_axaddr_0_addr(int_rd_req_desc_c_axaddr_0_addr),
                   .int_rd_req_desc_c_axaddr_1_addr(int_rd_req_desc_c_axaddr_1_addr),
                   .int_rd_req_desc_c_axaddr_2_addr(int_rd_req_desc_c_axaddr_2_addr),
                   .int_rd_req_desc_c_axaddr_3_addr(int_rd_req_desc_c_axaddr_3_addr),
                   .int_rd_req_desc_c_axid_0_axid(int_rd_req_desc_c_axid_0_axid),
                   .int_rd_req_desc_c_axid_1_axid(int_rd_req_desc_c_axid_1_axid),
                   .int_rd_req_desc_c_axid_2_axid(int_rd_req_desc_c_axid_2_axid),
                   .int_rd_req_desc_c_axid_3_axid(int_rd_req_desc_c_axid_3_axid),
                   .int_rd_req_desc_c_axuser_0_axuser(int_rd_req_desc_c_axuser_0_axuser),
                   .int_rd_req_desc_c_axuser_1_axuser(int_rd_req_desc_c_axuser_1_axuser),
                   .int_rd_req_desc_c_axuser_2_axuser(int_rd_req_desc_c_axuser_2_axuser),
                   .int_rd_req_desc_c_axuser_3_axuser(int_rd_req_desc_c_axuser_3_axuser),
                   .int_rd_req_desc_c_axuser_4_axuser(int_rd_req_desc_c_axuser_4_axuser),
                   .int_rd_req_desc_c_axuser_5_axuser(int_rd_req_desc_c_axuser_5_axuser),
                   .int_rd_req_desc_c_axuser_6_axuser(int_rd_req_desc_c_axuser_6_axuser),
                   .int_rd_req_desc_c_axuser_7_axuser(int_rd_req_desc_c_axuser_7_axuser),
                   .int_rd_req_desc_c_axuser_8_axuser(int_rd_req_desc_c_axuser_8_axuser),
                   .int_rd_req_desc_c_axuser_9_axuser(int_rd_req_desc_c_axuser_9_axuser),
                   .int_rd_req_desc_c_axuser_10_axuser(int_rd_req_desc_c_axuser_10_axuser),
                   .int_rd_req_desc_c_axuser_11_axuser(int_rd_req_desc_c_axuser_11_axuser),
                   .int_rd_req_desc_c_axuser_12_axuser(int_rd_req_desc_c_axuser_12_axuser),
                   .int_rd_req_desc_c_axuser_13_axuser(int_rd_req_desc_c_axuser_13_axuser),
                   .int_rd_req_desc_c_axuser_14_axuser(int_rd_req_desc_c_axuser_14_axuser),
                   .int_rd_req_desc_c_axuser_15_axuser(int_rd_req_desc_c_axuser_15_axuser),
                   .int_wr_req_desc_c_txn_type_wr_strb(int_wr_req_desc_c_txn_type_wr_strb),
                   .int_wr_req_desc_c_size_txn_size(int_wr_req_desc_c_size_txn_size),
                   .int_wr_req_desc_c_data_offset_addr(int_wr_req_desc_c_data_offset_addr),
                   .int_wr_req_desc_c_axsize_axsize(int_wr_req_desc_c_axsize_axsize),
                   .int_wr_req_desc_c_attr_axsnoop(int_wr_req_desc_c_attr_axsnoop),
                   .int_wr_req_desc_c_attr_axdomain(int_wr_req_desc_c_attr_axdomain),
                   .int_wr_req_desc_c_attr_axbar(int_wr_req_desc_c_attr_axbar),
                   .int_wr_req_desc_c_attr_awunique(int_wr_req_desc_c_attr_awunique),
                   .int_wr_req_desc_c_attr_axregion(int_wr_req_desc_c_attr_axregion),
                   .int_wr_req_desc_c_attr_axqos(int_wr_req_desc_c_attr_axqos),
                   .int_wr_req_desc_c_attr_axprot(int_wr_req_desc_c_attr_axprot),
                   .int_wr_req_desc_c_attr_axcache(int_wr_req_desc_c_attr_axcache),
                   .int_wr_req_desc_c_attr_axlock(int_wr_req_desc_c_attr_axlock),
                   .int_wr_req_desc_c_attr_axburst(int_wr_req_desc_c_attr_axburst),
                   .int_wr_req_desc_c_axaddr_0_addr(int_wr_req_desc_c_axaddr_0_addr),
                   .int_wr_req_desc_c_axaddr_1_addr(int_wr_req_desc_c_axaddr_1_addr),
                   .int_wr_req_desc_c_axaddr_2_addr(int_wr_req_desc_c_axaddr_2_addr),
                   .int_wr_req_desc_c_axaddr_3_addr(int_wr_req_desc_c_axaddr_3_addr),
                   .int_wr_req_desc_c_axid_0_axid(int_wr_req_desc_c_axid_0_axid),
                   .int_wr_req_desc_c_axid_1_axid(int_wr_req_desc_c_axid_1_axid),
                   .int_wr_req_desc_c_axid_2_axid(int_wr_req_desc_c_axid_2_axid),
                   .int_wr_req_desc_c_axid_3_axid(int_wr_req_desc_c_axid_3_axid),
                   .int_wr_req_desc_c_axuser_0_axuser(int_wr_req_desc_c_axuser_0_axuser),
                   .int_wr_req_desc_c_axuser_1_axuser(int_wr_req_desc_c_axuser_1_axuser),
                   .int_wr_req_desc_c_axuser_2_axuser(int_wr_req_desc_c_axuser_2_axuser),
                   .int_wr_req_desc_c_axuser_3_axuser(int_wr_req_desc_c_axuser_3_axuser),
                   .int_wr_req_desc_c_axuser_4_axuser(int_wr_req_desc_c_axuser_4_axuser),
                   .int_wr_req_desc_c_axuser_5_axuser(int_wr_req_desc_c_axuser_5_axuser),
                   .int_wr_req_desc_c_axuser_6_axuser(int_wr_req_desc_c_axuser_6_axuser),
                   .int_wr_req_desc_c_axuser_7_axuser(int_wr_req_desc_c_axuser_7_axuser),
                   .int_wr_req_desc_c_axuser_8_axuser(int_wr_req_desc_c_axuser_8_axuser),
                   .int_wr_req_desc_c_axuser_9_axuser(int_wr_req_desc_c_axuser_9_axuser),
                   .int_wr_req_desc_c_axuser_10_axuser(int_wr_req_desc_c_axuser_10_axuser),
                   .int_wr_req_desc_c_axuser_11_axuser(int_wr_req_desc_c_axuser_11_axuser),
                   .int_wr_req_desc_c_axuser_12_axuser(int_wr_req_desc_c_axuser_12_axuser),
                   .int_wr_req_desc_c_axuser_13_axuser(int_wr_req_desc_c_axuser_13_axuser),
                   .int_wr_req_desc_c_axuser_14_axuser(int_wr_req_desc_c_axuser_14_axuser),
                   .int_wr_req_desc_c_axuser_15_axuser(int_wr_req_desc_c_axuser_15_axuser),
                   .int_wr_req_desc_c_wuser_0_wuser(int_wr_req_desc_c_wuser_0_wuser),
                   .int_wr_req_desc_c_wuser_1_wuser(int_wr_req_desc_c_wuser_1_wuser),
                   .int_wr_req_desc_c_wuser_2_wuser(int_wr_req_desc_c_wuser_2_wuser),
                   .int_wr_req_desc_c_wuser_3_wuser(int_wr_req_desc_c_wuser_3_wuser),
                   .int_wr_req_desc_c_wuser_4_wuser(int_wr_req_desc_c_wuser_4_wuser),
                   .int_wr_req_desc_c_wuser_5_wuser(int_wr_req_desc_c_wuser_5_wuser),
                   .int_wr_req_desc_c_wuser_6_wuser(int_wr_req_desc_c_wuser_6_wuser),
                   .int_wr_req_desc_c_wuser_7_wuser(int_wr_req_desc_c_wuser_7_wuser),
                   .int_wr_req_desc_c_wuser_8_wuser(int_wr_req_desc_c_wuser_8_wuser),
                   .int_wr_req_desc_c_wuser_9_wuser(int_wr_req_desc_c_wuser_9_wuser),
                   .int_wr_req_desc_c_wuser_10_wuser(int_wr_req_desc_c_wuser_10_wuser),
                   .int_wr_req_desc_c_wuser_11_wuser(int_wr_req_desc_c_wuser_11_wuser),
                   .int_wr_req_desc_c_wuser_12_wuser(int_wr_req_desc_c_wuser_12_wuser),
                   .int_wr_req_desc_c_wuser_13_wuser(int_wr_req_desc_c_wuser_13_wuser),
                   .int_wr_req_desc_c_wuser_14_wuser(int_wr_req_desc_c_wuser_14_wuser),
                   .int_wr_req_desc_c_wuser_15_wuser(int_wr_req_desc_c_wuser_15_wuser),
                   .int_sn_resp_desc_c_resp_resp(int_sn_resp_desc_c_resp_resp),
                   .int_rd_req_desc_d_size_txn_size(int_rd_req_desc_d_size_txn_size),
                   .int_rd_req_desc_d_axsize_axsize(int_rd_req_desc_d_axsize_axsize),
                   .int_rd_req_desc_d_attr_axsnoop(int_rd_req_desc_d_attr_axsnoop),
                   .int_rd_req_desc_d_attr_axdomain(int_rd_req_desc_d_attr_axdomain),
                   .int_rd_req_desc_d_attr_axbar(int_rd_req_desc_d_attr_axbar),
                   .int_rd_req_desc_d_attr_axregion(int_rd_req_desc_d_attr_axregion),
                   .int_rd_req_desc_d_attr_axqos(int_rd_req_desc_d_attr_axqos),
                   .int_rd_req_desc_d_attr_axprot(int_rd_req_desc_d_attr_axprot),
                   .int_rd_req_desc_d_attr_axcache(int_rd_req_desc_d_attr_axcache),
                   .int_rd_req_desc_d_attr_axlock(int_rd_req_desc_d_attr_axlock),
                   .int_rd_req_desc_d_attr_axburst(int_rd_req_desc_d_attr_axburst),
                   .int_rd_req_desc_d_axaddr_0_addr(int_rd_req_desc_d_axaddr_0_addr),
                   .int_rd_req_desc_d_axaddr_1_addr(int_rd_req_desc_d_axaddr_1_addr),
                   .int_rd_req_desc_d_axaddr_2_addr(int_rd_req_desc_d_axaddr_2_addr),
                   .int_rd_req_desc_d_axaddr_3_addr(int_rd_req_desc_d_axaddr_3_addr),
                   .int_rd_req_desc_d_axid_0_axid(int_rd_req_desc_d_axid_0_axid),
                   .int_rd_req_desc_d_axid_1_axid(int_rd_req_desc_d_axid_1_axid),
                   .int_rd_req_desc_d_axid_2_axid(int_rd_req_desc_d_axid_2_axid),
                   .int_rd_req_desc_d_axid_3_axid(int_rd_req_desc_d_axid_3_axid),
                   .int_rd_req_desc_d_axuser_0_axuser(int_rd_req_desc_d_axuser_0_axuser),
                   .int_rd_req_desc_d_axuser_1_axuser(int_rd_req_desc_d_axuser_1_axuser),
                   .int_rd_req_desc_d_axuser_2_axuser(int_rd_req_desc_d_axuser_2_axuser),
                   .int_rd_req_desc_d_axuser_3_axuser(int_rd_req_desc_d_axuser_3_axuser),
                   .int_rd_req_desc_d_axuser_4_axuser(int_rd_req_desc_d_axuser_4_axuser),
                   .int_rd_req_desc_d_axuser_5_axuser(int_rd_req_desc_d_axuser_5_axuser),
                   .int_rd_req_desc_d_axuser_6_axuser(int_rd_req_desc_d_axuser_6_axuser),
                   .int_rd_req_desc_d_axuser_7_axuser(int_rd_req_desc_d_axuser_7_axuser),
                   .int_rd_req_desc_d_axuser_8_axuser(int_rd_req_desc_d_axuser_8_axuser),
                   .int_rd_req_desc_d_axuser_9_axuser(int_rd_req_desc_d_axuser_9_axuser),
                   .int_rd_req_desc_d_axuser_10_axuser(int_rd_req_desc_d_axuser_10_axuser),
                   .int_rd_req_desc_d_axuser_11_axuser(int_rd_req_desc_d_axuser_11_axuser),
                   .int_rd_req_desc_d_axuser_12_axuser(int_rd_req_desc_d_axuser_12_axuser),
                   .int_rd_req_desc_d_axuser_13_axuser(int_rd_req_desc_d_axuser_13_axuser),
                   .int_rd_req_desc_d_axuser_14_axuser(int_rd_req_desc_d_axuser_14_axuser),
                   .int_rd_req_desc_d_axuser_15_axuser(int_rd_req_desc_d_axuser_15_axuser),
                   .int_wr_req_desc_d_txn_type_wr_strb(int_wr_req_desc_d_txn_type_wr_strb),
                   .int_wr_req_desc_d_size_txn_size(int_wr_req_desc_d_size_txn_size),
                   .int_wr_req_desc_d_data_offset_addr(int_wr_req_desc_d_data_offset_addr),
                   .int_wr_req_desc_d_axsize_axsize(int_wr_req_desc_d_axsize_axsize),
                   .int_wr_req_desc_d_attr_axsnoop(int_wr_req_desc_d_attr_axsnoop),
                   .int_wr_req_desc_d_attr_axdomain(int_wr_req_desc_d_attr_axdomain),
                   .int_wr_req_desc_d_attr_axbar(int_wr_req_desc_d_attr_axbar),
                   .int_wr_req_desc_d_attr_awunique(int_wr_req_desc_d_attr_awunique),
                   .int_wr_req_desc_d_attr_axregion(int_wr_req_desc_d_attr_axregion),
                   .int_wr_req_desc_d_attr_axqos(int_wr_req_desc_d_attr_axqos),
                   .int_wr_req_desc_d_attr_axprot(int_wr_req_desc_d_attr_axprot),
                   .int_wr_req_desc_d_attr_axcache(int_wr_req_desc_d_attr_axcache),
                   .int_wr_req_desc_d_attr_axlock(int_wr_req_desc_d_attr_axlock),
                   .int_wr_req_desc_d_attr_axburst(int_wr_req_desc_d_attr_axburst),
                   .int_wr_req_desc_d_axaddr_0_addr(int_wr_req_desc_d_axaddr_0_addr),
                   .int_wr_req_desc_d_axaddr_1_addr(int_wr_req_desc_d_axaddr_1_addr),
                   .int_wr_req_desc_d_axaddr_2_addr(int_wr_req_desc_d_axaddr_2_addr),
                   .int_wr_req_desc_d_axaddr_3_addr(int_wr_req_desc_d_axaddr_3_addr),
                   .int_wr_req_desc_d_axid_0_axid(int_wr_req_desc_d_axid_0_axid),
                   .int_wr_req_desc_d_axid_1_axid(int_wr_req_desc_d_axid_1_axid),
                   .int_wr_req_desc_d_axid_2_axid(int_wr_req_desc_d_axid_2_axid),
                   .int_wr_req_desc_d_axid_3_axid(int_wr_req_desc_d_axid_3_axid),
                   .int_wr_req_desc_d_axuser_0_axuser(int_wr_req_desc_d_axuser_0_axuser),
                   .int_wr_req_desc_d_axuser_1_axuser(int_wr_req_desc_d_axuser_1_axuser),
                   .int_wr_req_desc_d_axuser_2_axuser(int_wr_req_desc_d_axuser_2_axuser),
                   .int_wr_req_desc_d_axuser_3_axuser(int_wr_req_desc_d_axuser_3_axuser),
                   .int_wr_req_desc_d_axuser_4_axuser(int_wr_req_desc_d_axuser_4_axuser),
                   .int_wr_req_desc_d_axuser_5_axuser(int_wr_req_desc_d_axuser_5_axuser),
                   .int_wr_req_desc_d_axuser_6_axuser(int_wr_req_desc_d_axuser_6_axuser),
                   .int_wr_req_desc_d_axuser_7_axuser(int_wr_req_desc_d_axuser_7_axuser),
                   .int_wr_req_desc_d_axuser_8_axuser(int_wr_req_desc_d_axuser_8_axuser),
                   .int_wr_req_desc_d_axuser_9_axuser(int_wr_req_desc_d_axuser_9_axuser),
                   .int_wr_req_desc_d_axuser_10_axuser(int_wr_req_desc_d_axuser_10_axuser),
                   .int_wr_req_desc_d_axuser_11_axuser(int_wr_req_desc_d_axuser_11_axuser),
                   .int_wr_req_desc_d_axuser_12_axuser(int_wr_req_desc_d_axuser_12_axuser),
                   .int_wr_req_desc_d_axuser_13_axuser(int_wr_req_desc_d_axuser_13_axuser),
                   .int_wr_req_desc_d_axuser_14_axuser(int_wr_req_desc_d_axuser_14_axuser),
                   .int_wr_req_desc_d_axuser_15_axuser(int_wr_req_desc_d_axuser_15_axuser),
                   .int_wr_req_desc_d_wuser_0_wuser(int_wr_req_desc_d_wuser_0_wuser),
                   .int_wr_req_desc_d_wuser_1_wuser(int_wr_req_desc_d_wuser_1_wuser),
                   .int_wr_req_desc_d_wuser_2_wuser(int_wr_req_desc_d_wuser_2_wuser),
                   .int_wr_req_desc_d_wuser_3_wuser(int_wr_req_desc_d_wuser_3_wuser),
                   .int_wr_req_desc_d_wuser_4_wuser(int_wr_req_desc_d_wuser_4_wuser),
                   .int_wr_req_desc_d_wuser_5_wuser(int_wr_req_desc_d_wuser_5_wuser),
                   .int_wr_req_desc_d_wuser_6_wuser(int_wr_req_desc_d_wuser_6_wuser),
                   .int_wr_req_desc_d_wuser_7_wuser(int_wr_req_desc_d_wuser_7_wuser),
                   .int_wr_req_desc_d_wuser_8_wuser(int_wr_req_desc_d_wuser_8_wuser),
                   .int_wr_req_desc_d_wuser_9_wuser(int_wr_req_desc_d_wuser_9_wuser),
                   .int_wr_req_desc_d_wuser_10_wuser(int_wr_req_desc_d_wuser_10_wuser),
                   .int_wr_req_desc_d_wuser_11_wuser(int_wr_req_desc_d_wuser_11_wuser),
                   .int_wr_req_desc_d_wuser_12_wuser(int_wr_req_desc_d_wuser_12_wuser),
                   .int_wr_req_desc_d_wuser_13_wuser(int_wr_req_desc_d_wuser_13_wuser),
                   .int_wr_req_desc_d_wuser_14_wuser(int_wr_req_desc_d_wuser_14_wuser),
                   .int_wr_req_desc_d_wuser_15_wuser(int_wr_req_desc_d_wuser_15_wuser),
                   .int_sn_resp_desc_d_resp_resp(int_sn_resp_desc_d_resp_resp),
                   .int_rd_req_desc_e_size_txn_size(int_rd_req_desc_e_size_txn_size),
                   .int_rd_req_desc_e_axsize_axsize(int_rd_req_desc_e_axsize_axsize),
                   .int_rd_req_desc_e_attr_axsnoop(int_rd_req_desc_e_attr_axsnoop),
                   .int_rd_req_desc_e_attr_axdomain(int_rd_req_desc_e_attr_axdomain),
                   .int_rd_req_desc_e_attr_axbar(int_rd_req_desc_e_attr_axbar),
                   .int_rd_req_desc_e_attr_axregion(int_rd_req_desc_e_attr_axregion),
                   .int_rd_req_desc_e_attr_axqos(int_rd_req_desc_e_attr_axqos),
                   .int_rd_req_desc_e_attr_axprot(int_rd_req_desc_e_attr_axprot),
                   .int_rd_req_desc_e_attr_axcache(int_rd_req_desc_e_attr_axcache),
                   .int_rd_req_desc_e_attr_axlock(int_rd_req_desc_e_attr_axlock),
                   .int_rd_req_desc_e_attr_axburst(int_rd_req_desc_e_attr_axburst),
                   .int_rd_req_desc_e_axaddr_0_addr(int_rd_req_desc_e_axaddr_0_addr),
                   .int_rd_req_desc_e_axaddr_1_addr(int_rd_req_desc_e_axaddr_1_addr),
                   .int_rd_req_desc_e_axaddr_2_addr(int_rd_req_desc_e_axaddr_2_addr),
                   .int_rd_req_desc_e_axaddr_3_addr(int_rd_req_desc_e_axaddr_3_addr),
                   .int_rd_req_desc_e_axid_0_axid(int_rd_req_desc_e_axid_0_axid),
                   .int_rd_req_desc_e_axid_1_axid(int_rd_req_desc_e_axid_1_axid),
                   .int_rd_req_desc_e_axid_2_axid(int_rd_req_desc_e_axid_2_axid),
                   .int_rd_req_desc_e_axid_3_axid(int_rd_req_desc_e_axid_3_axid),
                   .int_rd_req_desc_e_axuser_0_axuser(int_rd_req_desc_e_axuser_0_axuser),
                   .int_rd_req_desc_e_axuser_1_axuser(int_rd_req_desc_e_axuser_1_axuser),
                   .int_rd_req_desc_e_axuser_2_axuser(int_rd_req_desc_e_axuser_2_axuser),
                   .int_rd_req_desc_e_axuser_3_axuser(int_rd_req_desc_e_axuser_3_axuser),
                   .int_rd_req_desc_e_axuser_4_axuser(int_rd_req_desc_e_axuser_4_axuser),
                   .int_rd_req_desc_e_axuser_5_axuser(int_rd_req_desc_e_axuser_5_axuser),
                   .int_rd_req_desc_e_axuser_6_axuser(int_rd_req_desc_e_axuser_6_axuser),
                   .int_rd_req_desc_e_axuser_7_axuser(int_rd_req_desc_e_axuser_7_axuser),
                   .int_rd_req_desc_e_axuser_8_axuser(int_rd_req_desc_e_axuser_8_axuser),
                   .int_rd_req_desc_e_axuser_9_axuser(int_rd_req_desc_e_axuser_9_axuser),
                   .int_rd_req_desc_e_axuser_10_axuser(int_rd_req_desc_e_axuser_10_axuser),
                   .int_rd_req_desc_e_axuser_11_axuser(int_rd_req_desc_e_axuser_11_axuser),
                   .int_rd_req_desc_e_axuser_12_axuser(int_rd_req_desc_e_axuser_12_axuser),
                   .int_rd_req_desc_e_axuser_13_axuser(int_rd_req_desc_e_axuser_13_axuser),
                   .int_rd_req_desc_e_axuser_14_axuser(int_rd_req_desc_e_axuser_14_axuser),
                   .int_rd_req_desc_e_axuser_15_axuser(int_rd_req_desc_e_axuser_15_axuser),
                   .int_wr_req_desc_e_txn_type_wr_strb(int_wr_req_desc_e_txn_type_wr_strb),
                   .int_wr_req_desc_e_size_txn_size(int_wr_req_desc_e_size_txn_size),
                   .int_wr_req_desc_e_data_offset_addr(int_wr_req_desc_e_data_offset_addr),
                   .int_wr_req_desc_e_axsize_axsize(int_wr_req_desc_e_axsize_axsize),
                   .int_wr_req_desc_e_attr_axsnoop(int_wr_req_desc_e_attr_axsnoop),
                   .int_wr_req_desc_e_attr_axdomain(int_wr_req_desc_e_attr_axdomain),
                   .int_wr_req_desc_e_attr_axbar(int_wr_req_desc_e_attr_axbar),
                   .int_wr_req_desc_e_attr_awunique(int_wr_req_desc_e_attr_awunique),
                   .int_wr_req_desc_e_attr_axregion(int_wr_req_desc_e_attr_axregion),
                   .int_wr_req_desc_e_attr_axqos(int_wr_req_desc_e_attr_axqos),
                   .int_wr_req_desc_e_attr_axprot(int_wr_req_desc_e_attr_axprot),
                   .int_wr_req_desc_e_attr_axcache(int_wr_req_desc_e_attr_axcache),
                   .int_wr_req_desc_e_attr_axlock(int_wr_req_desc_e_attr_axlock),
                   .int_wr_req_desc_e_attr_axburst(int_wr_req_desc_e_attr_axburst),
                   .int_wr_req_desc_e_axaddr_0_addr(int_wr_req_desc_e_axaddr_0_addr),
                   .int_wr_req_desc_e_axaddr_1_addr(int_wr_req_desc_e_axaddr_1_addr),
                   .int_wr_req_desc_e_axaddr_2_addr(int_wr_req_desc_e_axaddr_2_addr),
                   .int_wr_req_desc_e_axaddr_3_addr(int_wr_req_desc_e_axaddr_3_addr),
                   .int_wr_req_desc_e_axid_0_axid(int_wr_req_desc_e_axid_0_axid),
                   .int_wr_req_desc_e_axid_1_axid(int_wr_req_desc_e_axid_1_axid),
                   .int_wr_req_desc_e_axid_2_axid(int_wr_req_desc_e_axid_2_axid),
                   .int_wr_req_desc_e_axid_3_axid(int_wr_req_desc_e_axid_3_axid),
                   .int_wr_req_desc_e_axuser_0_axuser(int_wr_req_desc_e_axuser_0_axuser),
                   .int_wr_req_desc_e_axuser_1_axuser(int_wr_req_desc_e_axuser_1_axuser),
                   .int_wr_req_desc_e_axuser_2_axuser(int_wr_req_desc_e_axuser_2_axuser),
                   .int_wr_req_desc_e_axuser_3_axuser(int_wr_req_desc_e_axuser_3_axuser),
                   .int_wr_req_desc_e_axuser_4_axuser(int_wr_req_desc_e_axuser_4_axuser),
                   .int_wr_req_desc_e_axuser_5_axuser(int_wr_req_desc_e_axuser_5_axuser),
                   .int_wr_req_desc_e_axuser_6_axuser(int_wr_req_desc_e_axuser_6_axuser),
                   .int_wr_req_desc_e_axuser_7_axuser(int_wr_req_desc_e_axuser_7_axuser),
                   .int_wr_req_desc_e_axuser_8_axuser(int_wr_req_desc_e_axuser_8_axuser),
                   .int_wr_req_desc_e_axuser_9_axuser(int_wr_req_desc_e_axuser_9_axuser),
                   .int_wr_req_desc_e_axuser_10_axuser(int_wr_req_desc_e_axuser_10_axuser),
                   .int_wr_req_desc_e_axuser_11_axuser(int_wr_req_desc_e_axuser_11_axuser),
                   .int_wr_req_desc_e_axuser_12_axuser(int_wr_req_desc_e_axuser_12_axuser),
                   .int_wr_req_desc_e_axuser_13_axuser(int_wr_req_desc_e_axuser_13_axuser),
                   .int_wr_req_desc_e_axuser_14_axuser(int_wr_req_desc_e_axuser_14_axuser),
                   .int_wr_req_desc_e_axuser_15_axuser(int_wr_req_desc_e_axuser_15_axuser),
                   .int_wr_req_desc_e_wuser_0_wuser(int_wr_req_desc_e_wuser_0_wuser),
                   .int_wr_req_desc_e_wuser_1_wuser(int_wr_req_desc_e_wuser_1_wuser),
                   .int_wr_req_desc_e_wuser_2_wuser(int_wr_req_desc_e_wuser_2_wuser),
                   .int_wr_req_desc_e_wuser_3_wuser(int_wr_req_desc_e_wuser_3_wuser),
                   .int_wr_req_desc_e_wuser_4_wuser(int_wr_req_desc_e_wuser_4_wuser),
                   .int_wr_req_desc_e_wuser_5_wuser(int_wr_req_desc_e_wuser_5_wuser),
                   .int_wr_req_desc_e_wuser_6_wuser(int_wr_req_desc_e_wuser_6_wuser),
                   .int_wr_req_desc_e_wuser_7_wuser(int_wr_req_desc_e_wuser_7_wuser),
                   .int_wr_req_desc_e_wuser_8_wuser(int_wr_req_desc_e_wuser_8_wuser),
                   .int_wr_req_desc_e_wuser_9_wuser(int_wr_req_desc_e_wuser_9_wuser),
                   .int_wr_req_desc_e_wuser_10_wuser(int_wr_req_desc_e_wuser_10_wuser),
                   .int_wr_req_desc_e_wuser_11_wuser(int_wr_req_desc_e_wuser_11_wuser),
                   .int_wr_req_desc_e_wuser_12_wuser(int_wr_req_desc_e_wuser_12_wuser),
                   .int_wr_req_desc_e_wuser_13_wuser(int_wr_req_desc_e_wuser_13_wuser),
                   .int_wr_req_desc_e_wuser_14_wuser(int_wr_req_desc_e_wuser_14_wuser),
                   .int_wr_req_desc_e_wuser_15_wuser(int_wr_req_desc_e_wuser_15_wuser),
                   .int_sn_resp_desc_e_resp_resp(int_sn_resp_desc_e_resp_resp),
                   .int_rd_req_desc_f_size_txn_size(int_rd_req_desc_f_size_txn_size),
                   .int_rd_req_desc_f_axsize_axsize(int_rd_req_desc_f_axsize_axsize),
                   .int_rd_req_desc_f_attr_axsnoop(int_rd_req_desc_f_attr_axsnoop),
                   .int_rd_req_desc_f_attr_axdomain(int_rd_req_desc_f_attr_axdomain),
                   .int_rd_req_desc_f_attr_axbar(int_rd_req_desc_f_attr_axbar),
                   .int_rd_req_desc_f_attr_axregion(int_rd_req_desc_f_attr_axregion),
                   .int_rd_req_desc_f_attr_axqos(int_rd_req_desc_f_attr_axqos),
                   .int_rd_req_desc_f_attr_axprot(int_rd_req_desc_f_attr_axprot),
                   .int_rd_req_desc_f_attr_axcache(int_rd_req_desc_f_attr_axcache),
                   .int_rd_req_desc_f_attr_axlock(int_rd_req_desc_f_attr_axlock),
                   .int_rd_req_desc_f_attr_axburst(int_rd_req_desc_f_attr_axburst),
                   .int_rd_req_desc_f_axaddr_0_addr(int_rd_req_desc_f_axaddr_0_addr),
                   .int_rd_req_desc_f_axaddr_1_addr(int_rd_req_desc_f_axaddr_1_addr),
                   .int_rd_req_desc_f_axaddr_2_addr(int_rd_req_desc_f_axaddr_2_addr),
                   .int_rd_req_desc_f_axaddr_3_addr(int_rd_req_desc_f_axaddr_3_addr),
                   .int_rd_req_desc_f_axid_0_axid(int_rd_req_desc_f_axid_0_axid),
                   .int_rd_req_desc_f_axid_1_axid(int_rd_req_desc_f_axid_1_axid),
                   .int_rd_req_desc_f_axid_2_axid(int_rd_req_desc_f_axid_2_axid),
                   .int_rd_req_desc_f_axid_3_axid(int_rd_req_desc_f_axid_3_axid),
                   .int_rd_req_desc_f_axuser_0_axuser(int_rd_req_desc_f_axuser_0_axuser),
                   .int_rd_req_desc_f_axuser_1_axuser(int_rd_req_desc_f_axuser_1_axuser),
                   .int_rd_req_desc_f_axuser_2_axuser(int_rd_req_desc_f_axuser_2_axuser),
                   .int_rd_req_desc_f_axuser_3_axuser(int_rd_req_desc_f_axuser_3_axuser),
                   .int_rd_req_desc_f_axuser_4_axuser(int_rd_req_desc_f_axuser_4_axuser),
                   .int_rd_req_desc_f_axuser_5_axuser(int_rd_req_desc_f_axuser_5_axuser),
                   .int_rd_req_desc_f_axuser_6_axuser(int_rd_req_desc_f_axuser_6_axuser),
                   .int_rd_req_desc_f_axuser_7_axuser(int_rd_req_desc_f_axuser_7_axuser),
                   .int_rd_req_desc_f_axuser_8_axuser(int_rd_req_desc_f_axuser_8_axuser),
                   .int_rd_req_desc_f_axuser_9_axuser(int_rd_req_desc_f_axuser_9_axuser),
                   .int_rd_req_desc_f_axuser_10_axuser(int_rd_req_desc_f_axuser_10_axuser),
                   .int_rd_req_desc_f_axuser_11_axuser(int_rd_req_desc_f_axuser_11_axuser),
                   .int_rd_req_desc_f_axuser_12_axuser(int_rd_req_desc_f_axuser_12_axuser),
                   .int_rd_req_desc_f_axuser_13_axuser(int_rd_req_desc_f_axuser_13_axuser),
                   .int_rd_req_desc_f_axuser_14_axuser(int_rd_req_desc_f_axuser_14_axuser),
                   .int_rd_req_desc_f_axuser_15_axuser(int_rd_req_desc_f_axuser_15_axuser),
                   .int_wr_req_desc_f_txn_type_wr_strb(int_wr_req_desc_f_txn_type_wr_strb),
                   .int_wr_req_desc_f_size_txn_size(int_wr_req_desc_f_size_txn_size),
                   .int_wr_req_desc_f_data_offset_addr(int_wr_req_desc_f_data_offset_addr),
                   .int_wr_req_desc_f_axsize_axsize(int_wr_req_desc_f_axsize_axsize),
                   .int_wr_req_desc_f_attr_axsnoop(int_wr_req_desc_f_attr_axsnoop),
                   .int_wr_req_desc_f_attr_axdomain(int_wr_req_desc_f_attr_axdomain),
                   .int_wr_req_desc_f_attr_axbar(int_wr_req_desc_f_attr_axbar),
                   .int_wr_req_desc_f_attr_awunique(int_wr_req_desc_f_attr_awunique),
                   .int_wr_req_desc_f_attr_axregion(int_wr_req_desc_f_attr_axregion),
                   .int_wr_req_desc_f_attr_axqos(int_wr_req_desc_f_attr_axqos),
                   .int_wr_req_desc_f_attr_axprot(int_wr_req_desc_f_attr_axprot),
                   .int_wr_req_desc_f_attr_axcache(int_wr_req_desc_f_attr_axcache),
                   .int_wr_req_desc_f_attr_axlock(int_wr_req_desc_f_attr_axlock),
                   .int_wr_req_desc_f_attr_axburst(int_wr_req_desc_f_attr_axburst),
                   .int_wr_req_desc_f_axaddr_0_addr(int_wr_req_desc_f_axaddr_0_addr),
                   .int_wr_req_desc_f_axaddr_1_addr(int_wr_req_desc_f_axaddr_1_addr),
                   .int_wr_req_desc_f_axaddr_2_addr(int_wr_req_desc_f_axaddr_2_addr),
                   .int_wr_req_desc_f_axaddr_3_addr(int_wr_req_desc_f_axaddr_3_addr),
                   .int_wr_req_desc_f_axid_0_axid(int_wr_req_desc_f_axid_0_axid),
                   .int_wr_req_desc_f_axid_1_axid(int_wr_req_desc_f_axid_1_axid),
                   .int_wr_req_desc_f_axid_2_axid(int_wr_req_desc_f_axid_2_axid),
                   .int_wr_req_desc_f_axid_3_axid(int_wr_req_desc_f_axid_3_axid),
                   .int_wr_req_desc_f_axuser_0_axuser(int_wr_req_desc_f_axuser_0_axuser),
                   .int_wr_req_desc_f_axuser_1_axuser(int_wr_req_desc_f_axuser_1_axuser),
                   .int_wr_req_desc_f_axuser_2_axuser(int_wr_req_desc_f_axuser_2_axuser),
                   .int_wr_req_desc_f_axuser_3_axuser(int_wr_req_desc_f_axuser_3_axuser),
                   .int_wr_req_desc_f_axuser_4_axuser(int_wr_req_desc_f_axuser_4_axuser),
                   .int_wr_req_desc_f_axuser_5_axuser(int_wr_req_desc_f_axuser_5_axuser),
                   .int_wr_req_desc_f_axuser_6_axuser(int_wr_req_desc_f_axuser_6_axuser),
                   .int_wr_req_desc_f_axuser_7_axuser(int_wr_req_desc_f_axuser_7_axuser),
                   .int_wr_req_desc_f_axuser_8_axuser(int_wr_req_desc_f_axuser_8_axuser),
                   .int_wr_req_desc_f_axuser_9_axuser(int_wr_req_desc_f_axuser_9_axuser),
                   .int_wr_req_desc_f_axuser_10_axuser(int_wr_req_desc_f_axuser_10_axuser),
                   .int_wr_req_desc_f_axuser_11_axuser(int_wr_req_desc_f_axuser_11_axuser),
                   .int_wr_req_desc_f_axuser_12_axuser(int_wr_req_desc_f_axuser_12_axuser),
                   .int_wr_req_desc_f_axuser_13_axuser(int_wr_req_desc_f_axuser_13_axuser),
                   .int_wr_req_desc_f_axuser_14_axuser(int_wr_req_desc_f_axuser_14_axuser),
                   .int_wr_req_desc_f_axuser_15_axuser(int_wr_req_desc_f_axuser_15_axuser),
                   .int_wr_req_desc_f_wuser_0_wuser(int_wr_req_desc_f_wuser_0_wuser),
                   .int_wr_req_desc_f_wuser_1_wuser(int_wr_req_desc_f_wuser_1_wuser),
                   .int_wr_req_desc_f_wuser_2_wuser(int_wr_req_desc_f_wuser_2_wuser),
                   .int_wr_req_desc_f_wuser_3_wuser(int_wr_req_desc_f_wuser_3_wuser),
                   .int_wr_req_desc_f_wuser_4_wuser(int_wr_req_desc_f_wuser_4_wuser),
                   .int_wr_req_desc_f_wuser_5_wuser(int_wr_req_desc_f_wuser_5_wuser),
                   .int_wr_req_desc_f_wuser_6_wuser(int_wr_req_desc_f_wuser_6_wuser),
                   .int_wr_req_desc_f_wuser_7_wuser(int_wr_req_desc_f_wuser_7_wuser),
                   .int_wr_req_desc_f_wuser_8_wuser(int_wr_req_desc_f_wuser_8_wuser),
                   .int_wr_req_desc_f_wuser_9_wuser(int_wr_req_desc_f_wuser_9_wuser),
                   .int_wr_req_desc_f_wuser_10_wuser(int_wr_req_desc_f_wuser_10_wuser),
                   .int_wr_req_desc_f_wuser_11_wuser(int_wr_req_desc_f_wuser_11_wuser),
                   .int_wr_req_desc_f_wuser_12_wuser(int_wr_req_desc_f_wuser_12_wuser),
                   .int_wr_req_desc_f_wuser_13_wuser(int_wr_req_desc_f_wuser_13_wuser),
                   .int_wr_req_desc_f_wuser_14_wuser(int_wr_req_desc_f_wuser_14_wuser),
                   .int_wr_req_desc_f_wuser_15_wuser(int_wr_req_desc_f_wuser_15_wuser),
                   .int_sn_resp_desc_f_resp_resp(int_sn_resp_desc_f_resp_resp),
                   // Inputs
                   .clk                    (clk),
                   .resetn                 (resetn),
                   .s_ace_usr_awid         (s_ace_usr_awid),
                   .s_ace_usr_awaddr       (s_ace_usr_awaddr),
                   .s_ace_usr_awlen        (s_ace_usr_awlen),
                   .s_ace_usr_awsize       (s_ace_usr_awsize),
                   .s_ace_usr_awburst      (s_ace_usr_awburst),
                   .s_ace_usr_awlock       (s_ace_usr_awlock),
                   .s_ace_usr_awcache      (s_ace_usr_awcache),
                   .s_ace_usr_awprot       (s_ace_usr_awprot),
                   .s_ace_usr_awqos        (s_ace_usr_awqos),
                   .s_ace_usr_awregion     (s_ace_usr_awregion),
                   .s_ace_usr_awuser       (s_ace_usr_awuser),
                   .s_ace_usr_awsnoop      (s_ace_usr_awsnoop),
                   .s_ace_usr_awdomain     (s_ace_usr_awdomain),
                   .s_ace_usr_awbar        (s_ace_usr_awbar),
                   .s_ace_usr_awunique     (s_ace_usr_awunique),
                   .s_ace_usr_awvalid      (s_ace_usr_awvalid),
                   .s_ace_usr_wdata        (s_ace_usr_wdata),
                   .s_ace_usr_wstrb        (s_ace_usr_wstrb),
                   .s_ace_usr_wlast        (s_ace_usr_wlast),
                   .s_ace_usr_wuser        (s_ace_usr_wuser),
                   .s_ace_usr_wvalid       (s_ace_usr_wvalid),
                   .s_ace_usr_bready       (s_ace_usr_bready),
                   .s_ace_usr_wack         (s_ace_usr_wack),
                   .s_ace_usr_arid         (s_ace_usr_arid),
                   .s_ace_usr_araddr       (s_ace_usr_araddr),
                   .s_ace_usr_arlen        (s_ace_usr_arlen),
                   .s_ace_usr_arsize       (s_ace_usr_arsize),
                   .s_ace_usr_arburst      (s_ace_usr_arburst),
                   .s_ace_usr_arlock       (s_ace_usr_arlock),
                   .s_ace_usr_arcache      (s_ace_usr_arcache),
                   .s_ace_usr_arprot       (s_ace_usr_arprot),
                   .s_ace_usr_arqos        (s_ace_usr_arqos),
                   .s_ace_usr_arregion     (s_ace_usr_arregion),
                   .s_ace_usr_aruser       (s_ace_usr_aruser),
                   .s_ace_usr_arsnoop      (s_ace_usr_arsnoop),
                   .s_ace_usr_ardomain     (s_ace_usr_ardomain),
                   .s_ace_usr_arbar        (s_ace_usr_arbar),
                   .s_ace_usr_arvalid      (s_ace_usr_arvalid),
                   .s_ace_usr_rready       (s_ace_usr_rready),
                   .s_ace_usr_rack         (s_ace_usr_rack),
                   .s_ace_usr_acready      (s_ace_usr_acready),
                   .s_ace_usr_crresp       (s_ace_usr_crresp),
                   .s_ace_usr_crvalid      (s_ace_usr_crvalid),
                   .s_ace_usr_cddata       (s_ace_usr_cddata),
                   .s_ace_usr_cdlast       (s_ace_usr_cdlast),
                   .s_ace_usr_cdvalid      (s_ace_usr_cdvalid),
                   .rb2uc_rd_data          (rb2uc_rd_data),
                   .rd_hm2uc_done          (rd_hm2uc_done),
                   .wr_hm2uc_done          (wr_hm2uc_done),
                   .rd_req_fifo_pop_desc_conn(rd_req_fifo_pop_desc_conn),
                   .wr_req_fifo_pop_desc_conn(wr_req_fifo_pop_desc_conn),
                   .sn_resp_fifo_pop_desc_conn(sn_resp_fifo_pop_desc_conn),
                   .sn_data_fifo_pop_desc_conn(sn_data_fifo_pop_desc_conn),
                   .int_bridge_identification_last_bridge(int_bridge_identification_last_bridge),
                   .int_version_major_ver  (int_version_major_ver),
                   .int_version_minor_ver  (int_version_minor_ver),
                   .int_bridge_type_type   (int_bridge_type_type),
                   .int_bridge_config_extend_wstrb(int_bridge_config_extend_wstrb),
                   .int_bridge_config_id_width(int_bridge_config_id_width),
                   .int_bridge_config_data_width(int_bridge_config_data_width),
                   .int_bridge_rd_user_config_ruser_width(int_bridge_rd_user_config_ruser_width),
                   .int_bridge_rd_user_config_aruser_width(int_bridge_rd_user_config_aruser_width),
                   .int_bridge_wr_user_config_buser_width(int_bridge_wr_user_config_buser_width),
                   .int_bridge_wr_user_config_wuser_width(int_bridge_wr_user_config_wuser_width),
                   .int_bridge_wr_user_config_awuser_width(int_bridge_wr_user_config_awuser_width),
                   .int_rd_max_desc_resp_max_desc(int_rd_max_desc_resp_max_desc),
                   .int_rd_max_desc_req_max_desc(int_rd_max_desc_req_max_desc),
                   .int_wr_max_desc_resp_max_desc(int_wr_max_desc_resp_max_desc),
                   .int_wr_max_desc_req_max_desc(int_wr_max_desc_req_max_desc),
                   .int_sn_max_desc_data_max_desc(int_sn_max_desc_data_max_desc),
                   .int_sn_max_desc_resp_max_desc(int_sn_max_desc_resp_max_desc),
                   .int_sn_max_desc_req_max_desc(int_sn_max_desc_req_max_desc),
                   .int_reset_dut_srst_3   (int_reset_dut_srst_3),
                   .int_reset_dut_srst_2   (int_reset_dut_srst_2),
                   .int_reset_dut_srst_1   (int_reset_dut_srst_1),
                   .int_reset_dut_srst_0   (int_reset_dut_srst_0),
                   .int_reset_srst         (int_reset_srst),
                   .int_mode_select_mode_0_1(int_mode_select_mode_0_1),
                   .int_intr_status_sn_data_fifo_nonempty(int_intr_status_sn_data_fifo_nonempty),
                   .int_intr_status_sn_resp_fifo_nonempty(int_intr_status_sn_resp_fifo_nonempty),
                   .int_intr_status_sn_req_comp(int_intr_status_sn_req_comp),
                   .int_intr_status_wr_resp_comp(int_intr_status_wr_resp_comp),
                   .int_intr_status_wr_req_fifo_nonempty(int_intr_status_wr_req_fifo_nonempty),
                   .int_intr_status_rd_resp_comp(int_intr_status_rd_resp_comp),
                   .int_intr_status_rd_req_fifo_nonempty(int_intr_status_rd_req_fifo_nonempty),
                   .int_intr_status_c2h    (int_intr_status_c2h),
                   .int_intr_status_error  (int_intr_status_error),
                   .int_intr_error_status_err_1(int_intr_error_status_err_1),
                   .int_intr_error_clear_clr_err_2(int_intr_error_clear_clr_err_2),
                   .int_intr_error_clear_clr_err_1(int_intr_error_clear_clr_err_1),
                   .int_intr_error_clear_clr_err_0(int_intr_error_clear_clr_err_0),
                   .int_intr_error_enable_en_err_2(int_intr_error_enable_en_err_2),
                   .int_intr_error_enable_en_err_1(int_intr_error_enable_en_err_1),
                   .int_intr_error_enable_en_err_0(int_intr_error_enable_en_err_0),
                   .int_rd_req_free_desc_desc(int_rd_req_free_desc_desc),
                   .int_rd_resp_fifo_push_desc_valid(int_rd_resp_fifo_push_desc_valid),
                   .int_rd_resp_fifo_push_desc_desc_index(int_rd_resp_fifo_push_desc_desc_index),
                   .int_rd_resp_intr_comp_clear_clr_comp(int_rd_resp_intr_comp_clear_clr_comp),
                   .int_rd_resp_intr_comp_enable_en_comp(int_rd_resp_intr_comp_enable_en_comp),
                   .int_wr_req_free_desc_desc(int_wr_req_free_desc_desc),
                   .int_wr_resp_fifo_push_desc_valid(int_wr_resp_fifo_push_desc_valid),
                   .int_wr_resp_fifo_push_desc_desc_index(int_wr_resp_fifo_push_desc_desc_index),
                   .int_wr_resp_intr_comp_clear_clr_comp(int_wr_resp_intr_comp_clear_clr_comp),
                   .int_wr_resp_intr_comp_enable_en_comp(int_wr_resp_intr_comp_enable_en_comp),
                   .int_sn_req_fifo_push_desc_valid(int_sn_req_fifo_push_desc_valid),
                   .int_sn_req_fifo_push_desc_desc_index(int_sn_req_fifo_push_desc_desc_index),
                   .int_sn_req_intr_comp_clear_clr_comp(int_sn_req_intr_comp_clear_clr_comp),
                   .int_sn_req_intr_comp_enable_en_comp(int_sn_req_intr_comp_enable_en_comp),
                   .int_sn_resp_free_desc_desc(int_sn_resp_free_desc_desc),
                   .int_sn_data_free_desc_desc(int_sn_data_free_desc_desc),
                   .int_intr_fifo_enable_en_sn_data_fifo_nonempty(int_intr_fifo_enable_en_sn_data_fifo_nonempty),
                   .int_intr_fifo_enable_en_sn_resp_fifo_nonempty(int_intr_fifo_enable_en_sn_resp_fifo_nonempty),
                   .int_intr_fifo_enable_en_wr_req_fifo_nonempty(int_intr_fifo_enable_en_wr_req_fifo_nonempty),
                   .int_intr_fifo_enable_en_rd_req_fifo_nonempty(int_intr_fifo_enable_en_rd_req_fifo_nonempty),
                   .int_rd_resp_desc_0_data_offset_addr(int_rd_resp_desc_0_data_offset_addr),
                   .int_rd_resp_desc_0_data_size_size(int_rd_resp_desc_0_data_size_size),
                   .int_rd_resp_desc_0_data_host_addr_0_addr(int_rd_resp_desc_0_data_host_addr_0_addr),
                   .int_rd_resp_desc_0_data_host_addr_1_addr(int_rd_resp_desc_0_data_host_addr_1_addr),
                   .int_rd_resp_desc_0_data_host_addr_2_addr(int_rd_resp_desc_0_data_host_addr_2_addr),
                   .int_rd_resp_desc_0_data_host_addr_3_addr(int_rd_resp_desc_0_data_host_addr_3_addr),
                   .int_rd_resp_desc_0_resp_resp(int_rd_resp_desc_0_resp_resp),
                   .int_rd_resp_desc_0_xid_0_xid(int_rd_resp_desc_0_xid_0_xid),
                   .int_rd_resp_desc_0_xid_1_xid(int_rd_resp_desc_0_xid_1_xid),
                   .int_rd_resp_desc_0_xid_2_xid(int_rd_resp_desc_0_xid_2_xid),
                   .int_rd_resp_desc_0_xid_3_xid(int_rd_resp_desc_0_xid_3_xid),
                   .int_rd_resp_desc_0_xuser_0_xuser(int_rd_resp_desc_0_xuser_0_xuser),
                   .int_rd_resp_desc_0_xuser_1_xuser(int_rd_resp_desc_0_xuser_1_xuser),
                   .int_rd_resp_desc_0_xuser_2_xuser(int_rd_resp_desc_0_xuser_2_xuser),
                   .int_rd_resp_desc_0_xuser_3_xuser(int_rd_resp_desc_0_xuser_3_xuser),
                   .int_rd_resp_desc_0_xuser_4_xuser(int_rd_resp_desc_0_xuser_4_xuser),
                   .int_rd_resp_desc_0_xuser_5_xuser(int_rd_resp_desc_0_xuser_5_xuser),
                   .int_rd_resp_desc_0_xuser_6_xuser(int_rd_resp_desc_0_xuser_6_xuser),
                   .int_rd_resp_desc_0_xuser_7_xuser(int_rd_resp_desc_0_xuser_7_xuser),
                   .int_rd_resp_desc_0_xuser_8_xuser(int_rd_resp_desc_0_xuser_8_xuser),
                   .int_rd_resp_desc_0_xuser_9_xuser(int_rd_resp_desc_0_xuser_9_xuser),
                   .int_rd_resp_desc_0_xuser_10_xuser(int_rd_resp_desc_0_xuser_10_xuser),
                   .int_rd_resp_desc_0_xuser_11_xuser(int_rd_resp_desc_0_xuser_11_xuser),
                   .int_rd_resp_desc_0_xuser_12_xuser(int_rd_resp_desc_0_xuser_12_xuser),
                   .int_rd_resp_desc_0_xuser_13_xuser(int_rd_resp_desc_0_xuser_13_xuser),
                   .int_rd_resp_desc_0_xuser_14_xuser(int_rd_resp_desc_0_xuser_14_xuser),
                   .int_rd_resp_desc_0_xuser_15_xuser(int_rd_resp_desc_0_xuser_15_xuser),
                   .int_wr_req_desc_0_data_host_addr_0_addr(int_wr_req_desc_0_data_host_addr_0_addr),
                   .int_wr_req_desc_0_data_host_addr_1_addr(int_wr_req_desc_0_data_host_addr_1_addr),
                   .int_wr_req_desc_0_data_host_addr_2_addr(int_wr_req_desc_0_data_host_addr_2_addr),
                   .int_wr_req_desc_0_data_host_addr_3_addr(int_wr_req_desc_0_data_host_addr_3_addr),
                   .int_wr_req_desc_0_wstrb_host_addr_0_addr(int_wr_req_desc_0_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_0_wstrb_host_addr_1_addr(int_wr_req_desc_0_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_0_wstrb_host_addr_2_addr(int_wr_req_desc_0_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_0_wstrb_host_addr_3_addr(int_wr_req_desc_0_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_0_resp_resp(int_wr_resp_desc_0_resp_resp),
                   .int_wr_resp_desc_0_xid_0_xid(int_wr_resp_desc_0_xid_0_xid),
                   .int_wr_resp_desc_0_xid_1_xid(int_wr_resp_desc_0_xid_1_xid),
                   .int_wr_resp_desc_0_xid_2_xid(int_wr_resp_desc_0_xid_2_xid),
                   .int_wr_resp_desc_0_xid_3_xid(int_wr_resp_desc_0_xid_3_xid),
                   .int_wr_resp_desc_0_xuser_0_xuser(int_wr_resp_desc_0_xuser_0_xuser),
                   .int_wr_resp_desc_0_xuser_1_xuser(int_wr_resp_desc_0_xuser_1_xuser),
                   .int_wr_resp_desc_0_xuser_2_xuser(int_wr_resp_desc_0_xuser_2_xuser),
                   .int_wr_resp_desc_0_xuser_3_xuser(int_wr_resp_desc_0_xuser_3_xuser),
                   .int_wr_resp_desc_0_xuser_4_xuser(int_wr_resp_desc_0_xuser_4_xuser),
                   .int_wr_resp_desc_0_xuser_5_xuser(int_wr_resp_desc_0_xuser_5_xuser),
                   .int_wr_resp_desc_0_xuser_6_xuser(int_wr_resp_desc_0_xuser_6_xuser),
                   .int_wr_resp_desc_0_xuser_7_xuser(int_wr_resp_desc_0_xuser_7_xuser),
                   .int_wr_resp_desc_0_xuser_8_xuser(int_wr_resp_desc_0_xuser_8_xuser),
                   .int_wr_resp_desc_0_xuser_9_xuser(int_wr_resp_desc_0_xuser_9_xuser),
                   .int_wr_resp_desc_0_xuser_10_xuser(int_wr_resp_desc_0_xuser_10_xuser),
                   .int_wr_resp_desc_0_xuser_11_xuser(int_wr_resp_desc_0_xuser_11_xuser),
                   .int_wr_resp_desc_0_xuser_12_xuser(int_wr_resp_desc_0_xuser_12_xuser),
                   .int_wr_resp_desc_0_xuser_13_xuser(int_wr_resp_desc_0_xuser_13_xuser),
                   .int_wr_resp_desc_0_xuser_14_xuser(int_wr_resp_desc_0_xuser_14_xuser),
                   .int_wr_resp_desc_0_xuser_15_xuser(int_wr_resp_desc_0_xuser_15_xuser),
                   .int_sn_req_desc_0_attr_acsnoop(int_sn_req_desc_0_attr_acsnoop),
                   .int_sn_req_desc_0_attr_acprot(int_sn_req_desc_0_attr_acprot),
                   .int_sn_req_desc_0_acaddr_0_addr(int_sn_req_desc_0_acaddr_0_addr),
                   .int_sn_req_desc_0_acaddr_1_addr(int_sn_req_desc_0_acaddr_1_addr),
                   .int_sn_req_desc_0_acaddr_2_addr(int_sn_req_desc_0_acaddr_2_addr),
                   .int_sn_req_desc_0_acaddr_3_addr(int_sn_req_desc_0_acaddr_3_addr),
                   .int_rd_resp_desc_1_data_offset_addr(int_rd_resp_desc_1_data_offset_addr),
                   .int_rd_resp_desc_1_data_size_size(int_rd_resp_desc_1_data_size_size),
                   .int_rd_resp_desc_1_data_host_addr_0_addr(int_rd_resp_desc_1_data_host_addr_0_addr),
                   .int_rd_resp_desc_1_data_host_addr_1_addr(int_rd_resp_desc_1_data_host_addr_1_addr),
                   .int_rd_resp_desc_1_data_host_addr_2_addr(int_rd_resp_desc_1_data_host_addr_2_addr),
                   .int_rd_resp_desc_1_data_host_addr_3_addr(int_rd_resp_desc_1_data_host_addr_3_addr),
                   .int_rd_resp_desc_1_resp_resp(int_rd_resp_desc_1_resp_resp),
                   .int_rd_resp_desc_1_xid_0_xid(int_rd_resp_desc_1_xid_0_xid),
                   .int_rd_resp_desc_1_xid_1_xid(int_rd_resp_desc_1_xid_1_xid),
                   .int_rd_resp_desc_1_xid_2_xid(int_rd_resp_desc_1_xid_2_xid),
                   .int_rd_resp_desc_1_xid_3_xid(int_rd_resp_desc_1_xid_3_xid),
                   .int_rd_resp_desc_1_xuser_0_xuser(int_rd_resp_desc_1_xuser_0_xuser),
                   .int_rd_resp_desc_1_xuser_1_xuser(int_rd_resp_desc_1_xuser_1_xuser),
                   .int_rd_resp_desc_1_xuser_2_xuser(int_rd_resp_desc_1_xuser_2_xuser),
                   .int_rd_resp_desc_1_xuser_3_xuser(int_rd_resp_desc_1_xuser_3_xuser),
                   .int_rd_resp_desc_1_xuser_4_xuser(int_rd_resp_desc_1_xuser_4_xuser),
                   .int_rd_resp_desc_1_xuser_5_xuser(int_rd_resp_desc_1_xuser_5_xuser),
                   .int_rd_resp_desc_1_xuser_6_xuser(int_rd_resp_desc_1_xuser_6_xuser),
                   .int_rd_resp_desc_1_xuser_7_xuser(int_rd_resp_desc_1_xuser_7_xuser),
                   .int_rd_resp_desc_1_xuser_8_xuser(int_rd_resp_desc_1_xuser_8_xuser),
                   .int_rd_resp_desc_1_xuser_9_xuser(int_rd_resp_desc_1_xuser_9_xuser),
                   .int_rd_resp_desc_1_xuser_10_xuser(int_rd_resp_desc_1_xuser_10_xuser),
                   .int_rd_resp_desc_1_xuser_11_xuser(int_rd_resp_desc_1_xuser_11_xuser),
                   .int_rd_resp_desc_1_xuser_12_xuser(int_rd_resp_desc_1_xuser_12_xuser),
                   .int_rd_resp_desc_1_xuser_13_xuser(int_rd_resp_desc_1_xuser_13_xuser),
                   .int_rd_resp_desc_1_xuser_14_xuser(int_rd_resp_desc_1_xuser_14_xuser),
                   .int_rd_resp_desc_1_xuser_15_xuser(int_rd_resp_desc_1_xuser_15_xuser),
                   .int_wr_req_desc_1_data_host_addr_0_addr(int_wr_req_desc_1_data_host_addr_0_addr),
                   .int_wr_req_desc_1_data_host_addr_1_addr(int_wr_req_desc_1_data_host_addr_1_addr),
                   .int_wr_req_desc_1_data_host_addr_2_addr(int_wr_req_desc_1_data_host_addr_2_addr),
                   .int_wr_req_desc_1_data_host_addr_3_addr(int_wr_req_desc_1_data_host_addr_3_addr),
                   .int_wr_req_desc_1_wstrb_host_addr_0_addr(int_wr_req_desc_1_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_1_wstrb_host_addr_1_addr(int_wr_req_desc_1_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_1_wstrb_host_addr_2_addr(int_wr_req_desc_1_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_1_wstrb_host_addr_3_addr(int_wr_req_desc_1_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_1_resp_resp(int_wr_resp_desc_1_resp_resp),
                   .int_wr_resp_desc_1_xid_0_xid(int_wr_resp_desc_1_xid_0_xid),
                   .int_wr_resp_desc_1_xid_1_xid(int_wr_resp_desc_1_xid_1_xid),
                   .int_wr_resp_desc_1_xid_2_xid(int_wr_resp_desc_1_xid_2_xid),
                   .int_wr_resp_desc_1_xid_3_xid(int_wr_resp_desc_1_xid_3_xid),
                   .int_wr_resp_desc_1_xuser_0_xuser(int_wr_resp_desc_1_xuser_0_xuser),
                   .int_wr_resp_desc_1_xuser_1_xuser(int_wr_resp_desc_1_xuser_1_xuser),
                   .int_wr_resp_desc_1_xuser_2_xuser(int_wr_resp_desc_1_xuser_2_xuser),
                   .int_wr_resp_desc_1_xuser_3_xuser(int_wr_resp_desc_1_xuser_3_xuser),
                   .int_wr_resp_desc_1_xuser_4_xuser(int_wr_resp_desc_1_xuser_4_xuser),
                   .int_wr_resp_desc_1_xuser_5_xuser(int_wr_resp_desc_1_xuser_5_xuser),
                   .int_wr_resp_desc_1_xuser_6_xuser(int_wr_resp_desc_1_xuser_6_xuser),
                   .int_wr_resp_desc_1_xuser_7_xuser(int_wr_resp_desc_1_xuser_7_xuser),
                   .int_wr_resp_desc_1_xuser_8_xuser(int_wr_resp_desc_1_xuser_8_xuser),
                   .int_wr_resp_desc_1_xuser_9_xuser(int_wr_resp_desc_1_xuser_9_xuser),
                   .int_wr_resp_desc_1_xuser_10_xuser(int_wr_resp_desc_1_xuser_10_xuser),
                   .int_wr_resp_desc_1_xuser_11_xuser(int_wr_resp_desc_1_xuser_11_xuser),
                   .int_wr_resp_desc_1_xuser_12_xuser(int_wr_resp_desc_1_xuser_12_xuser),
                   .int_wr_resp_desc_1_xuser_13_xuser(int_wr_resp_desc_1_xuser_13_xuser),
                   .int_wr_resp_desc_1_xuser_14_xuser(int_wr_resp_desc_1_xuser_14_xuser),
                   .int_wr_resp_desc_1_xuser_15_xuser(int_wr_resp_desc_1_xuser_15_xuser),
                   .int_sn_req_desc_1_attr_acsnoop(int_sn_req_desc_1_attr_acsnoop),
                   .int_sn_req_desc_1_attr_acprot(int_sn_req_desc_1_attr_acprot),
                   .int_sn_req_desc_1_acaddr_0_addr(int_sn_req_desc_1_acaddr_0_addr),
                   .int_sn_req_desc_1_acaddr_1_addr(int_sn_req_desc_1_acaddr_1_addr),
                   .int_sn_req_desc_1_acaddr_2_addr(int_sn_req_desc_1_acaddr_2_addr),
                   .int_sn_req_desc_1_acaddr_3_addr(int_sn_req_desc_1_acaddr_3_addr),
                   .int_rd_resp_desc_2_data_offset_addr(int_rd_resp_desc_2_data_offset_addr),
                   .int_rd_resp_desc_2_data_size_size(int_rd_resp_desc_2_data_size_size),
                   .int_rd_resp_desc_2_data_host_addr_0_addr(int_rd_resp_desc_2_data_host_addr_0_addr),
                   .int_rd_resp_desc_2_data_host_addr_1_addr(int_rd_resp_desc_2_data_host_addr_1_addr),
                   .int_rd_resp_desc_2_data_host_addr_2_addr(int_rd_resp_desc_2_data_host_addr_2_addr),
                   .int_rd_resp_desc_2_data_host_addr_3_addr(int_rd_resp_desc_2_data_host_addr_3_addr),
                   .int_rd_resp_desc_2_resp_resp(int_rd_resp_desc_2_resp_resp),
                   .int_rd_resp_desc_2_xid_0_xid(int_rd_resp_desc_2_xid_0_xid),
                   .int_rd_resp_desc_2_xid_1_xid(int_rd_resp_desc_2_xid_1_xid),
                   .int_rd_resp_desc_2_xid_2_xid(int_rd_resp_desc_2_xid_2_xid),
                   .int_rd_resp_desc_2_xid_3_xid(int_rd_resp_desc_2_xid_3_xid),
                   .int_rd_resp_desc_2_xuser_0_xuser(int_rd_resp_desc_2_xuser_0_xuser),
                   .int_rd_resp_desc_2_xuser_1_xuser(int_rd_resp_desc_2_xuser_1_xuser),
                   .int_rd_resp_desc_2_xuser_2_xuser(int_rd_resp_desc_2_xuser_2_xuser),
                   .int_rd_resp_desc_2_xuser_3_xuser(int_rd_resp_desc_2_xuser_3_xuser),
                   .int_rd_resp_desc_2_xuser_4_xuser(int_rd_resp_desc_2_xuser_4_xuser),
                   .int_rd_resp_desc_2_xuser_5_xuser(int_rd_resp_desc_2_xuser_5_xuser),
                   .int_rd_resp_desc_2_xuser_6_xuser(int_rd_resp_desc_2_xuser_6_xuser),
                   .int_rd_resp_desc_2_xuser_7_xuser(int_rd_resp_desc_2_xuser_7_xuser),
                   .int_rd_resp_desc_2_xuser_8_xuser(int_rd_resp_desc_2_xuser_8_xuser),
                   .int_rd_resp_desc_2_xuser_9_xuser(int_rd_resp_desc_2_xuser_9_xuser),
                   .int_rd_resp_desc_2_xuser_10_xuser(int_rd_resp_desc_2_xuser_10_xuser),
                   .int_rd_resp_desc_2_xuser_11_xuser(int_rd_resp_desc_2_xuser_11_xuser),
                   .int_rd_resp_desc_2_xuser_12_xuser(int_rd_resp_desc_2_xuser_12_xuser),
                   .int_rd_resp_desc_2_xuser_13_xuser(int_rd_resp_desc_2_xuser_13_xuser),
                   .int_rd_resp_desc_2_xuser_14_xuser(int_rd_resp_desc_2_xuser_14_xuser),
                   .int_rd_resp_desc_2_xuser_15_xuser(int_rd_resp_desc_2_xuser_15_xuser),
                   .int_wr_req_desc_2_data_host_addr_0_addr(int_wr_req_desc_2_data_host_addr_0_addr),
                   .int_wr_req_desc_2_data_host_addr_1_addr(int_wr_req_desc_2_data_host_addr_1_addr),
                   .int_wr_req_desc_2_data_host_addr_2_addr(int_wr_req_desc_2_data_host_addr_2_addr),
                   .int_wr_req_desc_2_data_host_addr_3_addr(int_wr_req_desc_2_data_host_addr_3_addr),
                   .int_wr_req_desc_2_wstrb_host_addr_0_addr(int_wr_req_desc_2_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_2_wstrb_host_addr_1_addr(int_wr_req_desc_2_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_2_wstrb_host_addr_2_addr(int_wr_req_desc_2_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_2_wstrb_host_addr_3_addr(int_wr_req_desc_2_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_2_resp_resp(int_wr_resp_desc_2_resp_resp),
                   .int_wr_resp_desc_2_xid_0_xid(int_wr_resp_desc_2_xid_0_xid),
                   .int_wr_resp_desc_2_xid_1_xid(int_wr_resp_desc_2_xid_1_xid),
                   .int_wr_resp_desc_2_xid_2_xid(int_wr_resp_desc_2_xid_2_xid),
                   .int_wr_resp_desc_2_xid_3_xid(int_wr_resp_desc_2_xid_3_xid),
                   .int_wr_resp_desc_2_xuser_0_xuser(int_wr_resp_desc_2_xuser_0_xuser),
                   .int_wr_resp_desc_2_xuser_1_xuser(int_wr_resp_desc_2_xuser_1_xuser),
                   .int_wr_resp_desc_2_xuser_2_xuser(int_wr_resp_desc_2_xuser_2_xuser),
                   .int_wr_resp_desc_2_xuser_3_xuser(int_wr_resp_desc_2_xuser_3_xuser),
                   .int_wr_resp_desc_2_xuser_4_xuser(int_wr_resp_desc_2_xuser_4_xuser),
                   .int_wr_resp_desc_2_xuser_5_xuser(int_wr_resp_desc_2_xuser_5_xuser),
                   .int_wr_resp_desc_2_xuser_6_xuser(int_wr_resp_desc_2_xuser_6_xuser),
                   .int_wr_resp_desc_2_xuser_7_xuser(int_wr_resp_desc_2_xuser_7_xuser),
                   .int_wr_resp_desc_2_xuser_8_xuser(int_wr_resp_desc_2_xuser_8_xuser),
                   .int_wr_resp_desc_2_xuser_9_xuser(int_wr_resp_desc_2_xuser_9_xuser),
                   .int_wr_resp_desc_2_xuser_10_xuser(int_wr_resp_desc_2_xuser_10_xuser),
                   .int_wr_resp_desc_2_xuser_11_xuser(int_wr_resp_desc_2_xuser_11_xuser),
                   .int_wr_resp_desc_2_xuser_12_xuser(int_wr_resp_desc_2_xuser_12_xuser),
                   .int_wr_resp_desc_2_xuser_13_xuser(int_wr_resp_desc_2_xuser_13_xuser),
                   .int_wr_resp_desc_2_xuser_14_xuser(int_wr_resp_desc_2_xuser_14_xuser),
                   .int_wr_resp_desc_2_xuser_15_xuser(int_wr_resp_desc_2_xuser_15_xuser),
                   .int_sn_req_desc_2_attr_acsnoop(int_sn_req_desc_2_attr_acsnoop),
                   .int_sn_req_desc_2_attr_acprot(int_sn_req_desc_2_attr_acprot),
                   .int_sn_req_desc_2_acaddr_0_addr(int_sn_req_desc_2_acaddr_0_addr),
                   .int_sn_req_desc_2_acaddr_1_addr(int_sn_req_desc_2_acaddr_1_addr),
                   .int_sn_req_desc_2_acaddr_2_addr(int_sn_req_desc_2_acaddr_2_addr),
                   .int_sn_req_desc_2_acaddr_3_addr(int_sn_req_desc_2_acaddr_3_addr),
                   .int_rd_resp_desc_3_data_offset_addr(int_rd_resp_desc_3_data_offset_addr),
                   .int_rd_resp_desc_3_data_size_size(int_rd_resp_desc_3_data_size_size),
                   .int_rd_resp_desc_3_data_host_addr_0_addr(int_rd_resp_desc_3_data_host_addr_0_addr),
                   .int_rd_resp_desc_3_data_host_addr_1_addr(int_rd_resp_desc_3_data_host_addr_1_addr),
                   .int_rd_resp_desc_3_data_host_addr_2_addr(int_rd_resp_desc_3_data_host_addr_2_addr),
                   .int_rd_resp_desc_3_data_host_addr_3_addr(int_rd_resp_desc_3_data_host_addr_3_addr),
                   .int_rd_resp_desc_3_resp_resp(int_rd_resp_desc_3_resp_resp),
                   .int_rd_resp_desc_3_xid_0_xid(int_rd_resp_desc_3_xid_0_xid),
                   .int_rd_resp_desc_3_xid_1_xid(int_rd_resp_desc_3_xid_1_xid),
                   .int_rd_resp_desc_3_xid_2_xid(int_rd_resp_desc_3_xid_2_xid),
                   .int_rd_resp_desc_3_xid_3_xid(int_rd_resp_desc_3_xid_3_xid),
                   .int_rd_resp_desc_3_xuser_0_xuser(int_rd_resp_desc_3_xuser_0_xuser),
                   .int_rd_resp_desc_3_xuser_1_xuser(int_rd_resp_desc_3_xuser_1_xuser),
                   .int_rd_resp_desc_3_xuser_2_xuser(int_rd_resp_desc_3_xuser_2_xuser),
                   .int_rd_resp_desc_3_xuser_3_xuser(int_rd_resp_desc_3_xuser_3_xuser),
                   .int_rd_resp_desc_3_xuser_4_xuser(int_rd_resp_desc_3_xuser_4_xuser),
                   .int_rd_resp_desc_3_xuser_5_xuser(int_rd_resp_desc_3_xuser_5_xuser),
                   .int_rd_resp_desc_3_xuser_6_xuser(int_rd_resp_desc_3_xuser_6_xuser),
                   .int_rd_resp_desc_3_xuser_7_xuser(int_rd_resp_desc_3_xuser_7_xuser),
                   .int_rd_resp_desc_3_xuser_8_xuser(int_rd_resp_desc_3_xuser_8_xuser),
                   .int_rd_resp_desc_3_xuser_9_xuser(int_rd_resp_desc_3_xuser_9_xuser),
                   .int_rd_resp_desc_3_xuser_10_xuser(int_rd_resp_desc_3_xuser_10_xuser),
                   .int_rd_resp_desc_3_xuser_11_xuser(int_rd_resp_desc_3_xuser_11_xuser),
                   .int_rd_resp_desc_3_xuser_12_xuser(int_rd_resp_desc_3_xuser_12_xuser),
                   .int_rd_resp_desc_3_xuser_13_xuser(int_rd_resp_desc_3_xuser_13_xuser),
                   .int_rd_resp_desc_3_xuser_14_xuser(int_rd_resp_desc_3_xuser_14_xuser),
                   .int_rd_resp_desc_3_xuser_15_xuser(int_rd_resp_desc_3_xuser_15_xuser),
                   .int_wr_req_desc_3_data_host_addr_0_addr(int_wr_req_desc_3_data_host_addr_0_addr),
                   .int_wr_req_desc_3_data_host_addr_1_addr(int_wr_req_desc_3_data_host_addr_1_addr),
                   .int_wr_req_desc_3_data_host_addr_2_addr(int_wr_req_desc_3_data_host_addr_2_addr),
                   .int_wr_req_desc_3_data_host_addr_3_addr(int_wr_req_desc_3_data_host_addr_3_addr),
                   .int_wr_req_desc_3_wstrb_host_addr_0_addr(int_wr_req_desc_3_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_3_wstrb_host_addr_1_addr(int_wr_req_desc_3_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_3_wstrb_host_addr_2_addr(int_wr_req_desc_3_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_3_wstrb_host_addr_3_addr(int_wr_req_desc_3_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_3_resp_resp(int_wr_resp_desc_3_resp_resp),
                   .int_wr_resp_desc_3_xid_0_xid(int_wr_resp_desc_3_xid_0_xid),
                   .int_wr_resp_desc_3_xid_1_xid(int_wr_resp_desc_3_xid_1_xid),
                   .int_wr_resp_desc_3_xid_2_xid(int_wr_resp_desc_3_xid_2_xid),
                   .int_wr_resp_desc_3_xid_3_xid(int_wr_resp_desc_3_xid_3_xid),
                   .int_wr_resp_desc_3_xuser_0_xuser(int_wr_resp_desc_3_xuser_0_xuser),
                   .int_wr_resp_desc_3_xuser_1_xuser(int_wr_resp_desc_3_xuser_1_xuser),
                   .int_wr_resp_desc_3_xuser_2_xuser(int_wr_resp_desc_3_xuser_2_xuser),
                   .int_wr_resp_desc_3_xuser_3_xuser(int_wr_resp_desc_3_xuser_3_xuser),
                   .int_wr_resp_desc_3_xuser_4_xuser(int_wr_resp_desc_3_xuser_4_xuser),
                   .int_wr_resp_desc_3_xuser_5_xuser(int_wr_resp_desc_3_xuser_5_xuser),
                   .int_wr_resp_desc_3_xuser_6_xuser(int_wr_resp_desc_3_xuser_6_xuser),
                   .int_wr_resp_desc_3_xuser_7_xuser(int_wr_resp_desc_3_xuser_7_xuser),
                   .int_wr_resp_desc_3_xuser_8_xuser(int_wr_resp_desc_3_xuser_8_xuser),
                   .int_wr_resp_desc_3_xuser_9_xuser(int_wr_resp_desc_3_xuser_9_xuser),
                   .int_wr_resp_desc_3_xuser_10_xuser(int_wr_resp_desc_3_xuser_10_xuser),
                   .int_wr_resp_desc_3_xuser_11_xuser(int_wr_resp_desc_3_xuser_11_xuser),
                   .int_wr_resp_desc_3_xuser_12_xuser(int_wr_resp_desc_3_xuser_12_xuser),
                   .int_wr_resp_desc_3_xuser_13_xuser(int_wr_resp_desc_3_xuser_13_xuser),
                   .int_wr_resp_desc_3_xuser_14_xuser(int_wr_resp_desc_3_xuser_14_xuser),
                   .int_wr_resp_desc_3_xuser_15_xuser(int_wr_resp_desc_3_xuser_15_xuser),
                   .int_sn_req_desc_3_attr_acsnoop(int_sn_req_desc_3_attr_acsnoop),
                   .int_sn_req_desc_3_attr_acprot(int_sn_req_desc_3_attr_acprot),
                   .int_sn_req_desc_3_acaddr_0_addr(int_sn_req_desc_3_acaddr_0_addr),
                   .int_sn_req_desc_3_acaddr_1_addr(int_sn_req_desc_3_acaddr_1_addr),
                   .int_sn_req_desc_3_acaddr_2_addr(int_sn_req_desc_3_acaddr_2_addr),
                   .int_sn_req_desc_3_acaddr_3_addr(int_sn_req_desc_3_acaddr_3_addr),
                   .int_rd_resp_desc_4_data_offset_addr(int_rd_resp_desc_4_data_offset_addr),
                   .int_rd_resp_desc_4_data_size_size(int_rd_resp_desc_4_data_size_size),
                   .int_rd_resp_desc_4_data_host_addr_0_addr(int_rd_resp_desc_4_data_host_addr_0_addr),
                   .int_rd_resp_desc_4_data_host_addr_1_addr(int_rd_resp_desc_4_data_host_addr_1_addr),
                   .int_rd_resp_desc_4_data_host_addr_2_addr(int_rd_resp_desc_4_data_host_addr_2_addr),
                   .int_rd_resp_desc_4_data_host_addr_3_addr(int_rd_resp_desc_4_data_host_addr_3_addr),
                   .int_rd_resp_desc_4_resp_resp(int_rd_resp_desc_4_resp_resp),
                   .int_rd_resp_desc_4_xid_0_xid(int_rd_resp_desc_4_xid_0_xid),
                   .int_rd_resp_desc_4_xid_1_xid(int_rd_resp_desc_4_xid_1_xid),
                   .int_rd_resp_desc_4_xid_2_xid(int_rd_resp_desc_4_xid_2_xid),
                   .int_rd_resp_desc_4_xid_3_xid(int_rd_resp_desc_4_xid_3_xid),
                   .int_rd_resp_desc_4_xuser_0_xuser(int_rd_resp_desc_4_xuser_0_xuser),
                   .int_rd_resp_desc_4_xuser_1_xuser(int_rd_resp_desc_4_xuser_1_xuser),
                   .int_rd_resp_desc_4_xuser_2_xuser(int_rd_resp_desc_4_xuser_2_xuser),
                   .int_rd_resp_desc_4_xuser_3_xuser(int_rd_resp_desc_4_xuser_3_xuser),
                   .int_rd_resp_desc_4_xuser_4_xuser(int_rd_resp_desc_4_xuser_4_xuser),
                   .int_rd_resp_desc_4_xuser_5_xuser(int_rd_resp_desc_4_xuser_5_xuser),
                   .int_rd_resp_desc_4_xuser_6_xuser(int_rd_resp_desc_4_xuser_6_xuser),
                   .int_rd_resp_desc_4_xuser_7_xuser(int_rd_resp_desc_4_xuser_7_xuser),
                   .int_rd_resp_desc_4_xuser_8_xuser(int_rd_resp_desc_4_xuser_8_xuser),
                   .int_rd_resp_desc_4_xuser_9_xuser(int_rd_resp_desc_4_xuser_9_xuser),
                   .int_rd_resp_desc_4_xuser_10_xuser(int_rd_resp_desc_4_xuser_10_xuser),
                   .int_rd_resp_desc_4_xuser_11_xuser(int_rd_resp_desc_4_xuser_11_xuser),
                   .int_rd_resp_desc_4_xuser_12_xuser(int_rd_resp_desc_4_xuser_12_xuser),
                   .int_rd_resp_desc_4_xuser_13_xuser(int_rd_resp_desc_4_xuser_13_xuser),
                   .int_rd_resp_desc_4_xuser_14_xuser(int_rd_resp_desc_4_xuser_14_xuser),
                   .int_rd_resp_desc_4_xuser_15_xuser(int_rd_resp_desc_4_xuser_15_xuser),
                   .int_wr_req_desc_4_data_host_addr_0_addr(int_wr_req_desc_4_data_host_addr_0_addr),
                   .int_wr_req_desc_4_data_host_addr_1_addr(int_wr_req_desc_4_data_host_addr_1_addr),
                   .int_wr_req_desc_4_data_host_addr_2_addr(int_wr_req_desc_4_data_host_addr_2_addr),
                   .int_wr_req_desc_4_data_host_addr_3_addr(int_wr_req_desc_4_data_host_addr_3_addr),
                   .int_wr_req_desc_4_wstrb_host_addr_0_addr(int_wr_req_desc_4_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_4_wstrb_host_addr_1_addr(int_wr_req_desc_4_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_4_wstrb_host_addr_2_addr(int_wr_req_desc_4_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_4_wstrb_host_addr_3_addr(int_wr_req_desc_4_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_4_resp_resp(int_wr_resp_desc_4_resp_resp),
                   .int_wr_resp_desc_4_xid_0_xid(int_wr_resp_desc_4_xid_0_xid),
                   .int_wr_resp_desc_4_xid_1_xid(int_wr_resp_desc_4_xid_1_xid),
                   .int_wr_resp_desc_4_xid_2_xid(int_wr_resp_desc_4_xid_2_xid),
                   .int_wr_resp_desc_4_xid_3_xid(int_wr_resp_desc_4_xid_3_xid),
                   .int_wr_resp_desc_4_xuser_0_xuser(int_wr_resp_desc_4_xuser_0_xuser),
                   .int_wr_resp_desc_4_xuser_1_xuser(int_wr_resp_desc_4_xuser_1_xuser),
                   .int_wr_resp_desc_4_xuser_2_xuser(int_wr_resp_desc_4_xuser_2_xuser),
                   .int_wr_resp_desc_4_xuser_3_xuser(int_wr_resp_desc_4_xuser_3_xuser),
                   .int_wr_resp_desc_4_xuser_4_xuser(int_wr_resp_desc_4_xuser_4_xuser),
                   .int_wr_resp_desc_4_xuser_5_xuser(int_wr_resp_desc_4_xuser_5_xuser),
                   .int_wr_resp_desc_4_xuser_6_xuser(int_wr_resp_desc_4_xuser_6_xuser),
                   .int_wr_resp_desc_4_xuser_7_xuser(int_wr_resp_desc_4_xuser_7_xuser),
                   .int_wr_resp_desc_4_xuser_8_xuser(int_wr_resp_desc_4_xuser_8_xuser),
                   .int_wr_resp_desc_4_xuser_9_xuser(int_wr_resp_desc_4_xuser_9_xuser),
                   .int_wr_resp_desc_4_xuser_10_xuser(int_wr_resp_desc_4_xuser_10_xuser),
                   .int_wr_resp_desc_4_xuser_11_xuser(int_wr_resp_desc_4_xuser_11_xuser),
                   .int_wr_resp_desc_4_xuser_12_xuser(int_wr_resp_desc_4_xuser_12_xuser),
                   .int_wr_resp_desc_4_xuser_13_xuser(int_wr_resp_desc_4_xuser_13_xuser),
                   .int_wr_resp_desc_4_xuser_14_xuser(int_wr_resp_desc_4_xuser_14_xuser),
                   .int_wr_resp_desc_4_xuser_15_xuser(int_wr_resp_desc_4_xuser_15_xuser),
                   .int_sn_req_desc_4_attr_acsnoop(int_sn_req_desc_4_attr_acsnoop),
                   .int_sn_req_desc_4_attr_acprot(int_sn_req_desc_4_attr_acprot),
                   .int_sn_req_desc_4_acaddr_0_addr(int_sn_req_desc_4_acaddr_0_addr),
                   .int_sn_req_desc_4_acaddr_1_addr(int_sn_req_desc_4_acaddr_1_addr),
                   .int_sn_req_desc_4_acaddr_2_addr(int_sn_req_desc_4_acaddr_2_addr),
                   .int_sn_req_desc_4_acaddr_3_addr(int_sn_req_desc_4_acaddr_3_addr),
                   .int_rd_resp_desc_5_data_offset_addr(int_rd_resp_desc_5_data_offset_addr),
                   .int_rd_resp_desc_5_data_size_size(int_rd_resp_desc_5_data_size_size),
                   .int_rd_resp_desc_5_data_host_addr_0_addr(int_rd_resp_desc_5_data_host_addr_0_addr),
                   .int_rd_resp_desc_5_data_host_addr_1_addr(int_rd_resp_desc_5_data_host_addr_1_addr),
                   .int_rd_resp_desc_5_data_host_addr_2_addr(int_rd_resp_desc_5_data_host_addr_2_addr),
                   .int_rd_resp_desc_5_data_host_addr_3_addr(int_rd_resp_desc_5_data_host_addr_3_addr),
                   .int_rd_resp_desc_5_resp_resp(int_rd_resp_desc_5_resp_resp),
                   .int_rd_resp_desc_5_xid_0_xid(int_rd_resp_desc_5_xid_0_xid),
                   .int_rd_resp_desc_5_xid_1_xid(int_rd_resp_desc_5_xid_1_xid),
                   .int_rd_resp_desc_5_xid_2_xid(int_rd_resp_desc_5_xid_2_xid),
                   .int_rd_resp_desc_5_xid_3_xid(int_rd_resp_desc_5_xid_3_xid),
                   .int_rd_resp_desc_5_xuser_0_xuser(int_rd_resp_desc_5_xuser_0_xuser),
                   .int_rd_resp_desc_5_xuser_1_xuser(int_rd_resp_desc_5_xuser_1_xuser),
                   .int_rd_resp_desc_5_xuser_2_xuser(int_rd_resp_desc_5_xuser_2_xuser),
                   .int_rd_resp_desc_5_xuser_3_xuser(int_rd_resp_desc_5_xuser_3_xuser),
                   .int_rd_resp_desc_5_xuser_4_xuser(int_rd_resp_desc_5_xuser_4_xuser),
                   .int_rd_resp_desc_5_xuser_5_xuser(int_rd_resp_desc_5_xuser_5_xuser),
                   .int_rd_resp_desc_5_xuser_6_xuser(int_rd_resp_desc_5_xuser_6_xuser),
                   .int_rd_resp_desc_5_xuser_7_xuser(int_rd_resp_desc_5_xuser_7_xuser),
                   .int_rd_resp_desc_5_xuser_8_xuser(int_rd_resp_desc_5_xuser_8_xuser),
                   .int_rd_resp_desc_5_xuser_9_xuser(int_rd_resp_desc_5_xuser_9_xuser),
                   .int_rd_resp_desc_5_xuser_10_xuser(int_rd_resp_desc_5_xuser_10_xuser),
                   .int_rd_resp_desc_5_xuser_11_xuser(int_rd_resp_desc_5_xuser_11_xuser),
                   .int_rd_resp_desc_5_xuser_12_xuser(int_rd_resp_desc_5_xuser_12_xuser),
                   .int_rd_resp_desc_5_xuser_13_xuser(int_rd_resp_desc_5_xuser_13_xuser),
                   .int_rd_resp_desc_5_xuser_14_xuser(int_rd_resp_desc_5_xuser_14_xuser),
                   .int_rd_resp_desc_5_xuser_15_xuser(int_rd_resp_desc_5_xuser_15_xuser),
                   .int_wr_req_desc_5_data_host_addr_0_addr(int_wr_req_desc_5_data_host_addr_0_addr),
                   .int_wr_req_desc_5_data_host_addr_1_addr(int_wr_req_desc_5_data_host_addr_1_addr),
                   .int_wr_req_desc_5_data_host_addr_2_addr(int_wr_req_desc_5_data_host_addr_2_addr),
                   .int_wr_req_desc_5_data_host_addr_3_addr(int_wr_req_desc_5_data_host_addr_3_addr),
                   .int_wr_req_desc_5_wstrb_host_addr_0_addr(int_wr_req_desc_5_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_5_wstrb_host_addr_1_addr(int_wr_req_desc_5_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_5_wstrb_host_addr_2_addr(int_wr_req_desc_5_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_5_wstrb_host_addr_3_addr(int_wr_req_desc_5_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_5_resp_resp(int_wr_resp_desc_5_resp_resp),
                   .int_wr_resp_desc_5_xid_0_xid(int_wr_resp_desc_5_xid_0_xid),
                   .int_wr_resp_desc_5_xid_1_xid(int_wr_resp_desc_5_xid_1_xid),
                   .int_wr_resp_desc_5_xid_2_xid(int_wr_resp_desc_5_xid_2_xid),
                   .int_wr_resp_desc_5_xid_3_xid(int_wr_resp_desc_5_xid_3_xid),
                   .int_wr_resp_desc_5_xuser_0_xuser(int_wr_resp_desc_5_xuser_0_xuser),
                   .int_wr_resp_desc_5_xuser_1_xuser(int_wr_resp_desc_5_xuser_1_xuser),
                   .int_wr_resp_desc_5_xuser_2_xuser(int_wr_resp_desc_5_xuser_2_xuser),
                   .int_wr_resp_desc_5_xuser_3_xuser(int_wr_resp_desc_5_xuser_3_xuser),
                   .int_wr_resp_desc_5_xuser_4_xuser(int_wr_resp_desc_5_xuser_4_xuser),
                   .int_wr_resp_desc_5_xuser_5_xuser(int_wr_resp_desc_5_xuser_5_xuser),
                   .int_wr_resp_desc_5_xuser_6_xuser(int_wr_resp_desc_5_xuser_6_xuser),
                   .int_wr_resp_desc_5_xuser_7_xuser(int_wr_resp_desc_5_xuser_7_xuser),
                   .int_wr_resp_desc_5_xuser_8_xuser(int_wr_resp_desc_5_xuser_8_xuser),
                   .int_wr_resp_desc_5_xuser_9_xuser(int_wr_resp_desc_5_xuser_9_xuser),
                   .int_wr_resp_desc_5_xuser_10_xuser(int_wr_resp_desc_5_xuser_10_xuser),
                   .int_wr_resp_desc_5_xuser_11_xuser(int_wr_resp_desc_5_xuser_11_xuser),
                   .int_wr_resp_desc_5_xuser_12_xuser(int_wr_resp_desc_5_xuser_12_xuser),
                   .int_wr_resp_desc_5_xuser_13_xuser(int_wr_resp_desc_5_xuser_13_xuser),
                   .int_wr_resp_desc_5_xuser_14_xuser(int_wr_resp_desc_5_xuser_14_xuser),
                   .int_wr_resp_desc_5_xuser_15_xuser(int_wr_resp_desc_5_xuser_15_xuser),
                   .int_sn_req_desc_5_attr_acsnoop(int_sn_req_desc_5_attr_acsnoop),
                   .int_sn_req_desc_5_attr_acprot(int_sn_req_desc_5_attr_acprot),
                   .int_sn_req_desc_5_acaddr_0_addr(int_sn_req_desc_5_acaddr_0_addr),
                   .int_sn_req_desc_5_acaddr_1_addr(int_sn_req_desc_5_acaddr_1_addr),
                   .int_sn_req_desc_5_acaddr_2_addr(int_sn_req_desc_5_acaddr_2_addr),
                   .int_sn_req_desc_5_acaddr_3_addr(int_sn_req_desc_5_acaddr_3_addr),
                   .int_rd_resp_desc_6_data_offset_addr(int_rd_resp_desc_6_data_offset_addr),
                   .int_rd_resp_desc_6_data_size_size(int_rd_resp_desc_6_data_size_size),
                   .int_rd_resp_desc_6_data_host_addr_0_addr(int_rd_resp_desc_6_data_host_addr_0_addr),
                   .int_rd_resp_desc_6_data_host_addr_1_addr(int_rd_resp_desc_6_data_host_addr_1_addr),
                   .int_rd_resp_desc_6_data_host_addr_2_addr(int_rd_resp_desc_6_data_host_addr_2_addr),
                   .int_rd_resp_desc_6_data_host_addr_3_addr(int_rd_resp_desc_6_data_host_addr_3_addr),
                   .int_rd_resp_desc_6_resp_resp(int_rd_resp_desc_6_resp_resp),
                   .int_rd_resp_desc_6_xid_0_xid(int_rd_resp_desc_6_xid_0_xid),
                   .int_rd_resp_desc_6_xid_1_xid(int_rd_resp_desc_6_xid_1_xid),
                   .int_rd_resp_desc_6_xid_2_xid(int_rd_resp_desc_6_xid_2_xid),
                   .int_rd_resp_desc_6_xid_3_xid(int_rd_resp_desc_6_xid_3_xid),
                   .int_rd_resp_desc_6_xuser_0_xuser(int_rd_resp_desc_6_xuser_0_xuser),
                   .int_rd_resp_desc_6_xuser_1_xuser(int_rd_resp_desc_6_xuser_1_xuser),
                   .int_rd_resp_desc_6_xuser_2_xuser(int_rd_resp_desc_6_xuser_2_xuser),
                   .int_rd_resp_desc_6_xuser_3_xuser(int_rd_resp_desc_6_xuser_3_xuser),
                   .int_rd_resp_desc_6_xuser_4_xuser(int_rd_resp_desc_6_xuser_4_xuser),
                   .int_rd_resp_desc_6_xuser_5_xuser(int_rd_resp_desc_6_xuser_5_xuser),
                   .int_rd_resp_desc_6_xuser_6_xuser(int_rd_resp_desc_6_xuser_6_xuser),
                   .int_rd_resp_desc_6_xuser_7_xuser(int_rd_resp_desc_6_xuser_7_xuser),
                   .int_rd_resp_desc_6_xuser_8_xuser(int_rd_resp_desc_6_xuser_8_xuser),
                   .int_rd_resp_desc_6_xuser_9_xuser(int_rd_resp_desc_6_xuser_9_xuser),
                   .int_rd_resp_desc_6_xuser_10_xuser(int_rd_resp_desc_6_xuser_10_xuser),
                   .int_rd_resp_desc_6_xuser_11_xuser(int_rd_resp_desc_6_xuser_11_xuser),
                   .int_rd_resp_desc_6_xuser_12_xuser(int_rd_resp_desc_6_xuser_12_xuser),
                   .int_rd_resp_desc_6_xuser_13_xuser(int_rd_resp_desc_6_xuser_13_xuser),
                   .int_rd_resp_desc_6_xuser_14_xuser(int_rd_resp_desc_6_xuser_14_xuser),
                   .int_rd_resp_desc_6_xuser_15_xuser(int_rd_resp_desc_6_xuser_15_xuser),
                   .int_wr_req_desc_6_data_host_addr_0_addr(int_wr_req_desc_6_data_host_addr_0_addr),
                   .int_wr_req_desc_6_data_host_addr_1_addr(int_wr_req_desc_6_data_host_addr_1_addr),
                   .int_wr_req_desc_6_data_host_addr_2_addr(int_wr_req_desc_6_data_host_addr_2_addr),
                   .int_wr_req_desc_6_data_host_addr_3_addr(int_wr_req_desc_6_data_host_addr_3_addr),
                   .int_wr_req_desc_6_wstrb_host_addr_0_addr(int_wr_req_desc_6_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_6_wstrb_host_addr_1_addr(int_wr_req_desc_6_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_6_wstrb_host_addr_2_addr(int_wr_req_desc_6_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_6_wstrb_host_addr_3_addr(int_wr_req_desc_6_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_6_resp_resp(int_wr_resp_desc_6_resp_resp),
                   .int_wr_resp_desc_6_xid_0_xid(int_wr_resp_desc_6_xid_0_xid),
                   .int_wr_resp_desc_6_xid_1_xid(int_wr_resp_desc_6_xid_1_xid),
                   .int_wr_resp_desc_6_xid_2_xid(int_wr_resp_desc_6_xid_2_xid),
                   .int_wr_resp_desc_6_xid_3_xid(int_wr_resp_desc_6_xid_3_xid),
                   .int_wr_resp_desc_6_xuser_0_xuser(int_wr_resp_desc_6_xuser_0_xuser),
                   .int_wr_resp_desc_6_xuser_1_xuser(int_wr_resp_desc_6_xuser_1_xuser),
                   .int_wr_resp_desc_6_xuser_2_xuser(int_wr_resp_desc_6_xuser_2_xuser),
                   .int_wr_resp_desc_6_xuser_3_xuser(int_wr_resp_desc_6_xuser_3_xuser),
                   .int_wr_resp_desc_6_xuser_4_xuser(int_wr_resp_desc_6_xuser_4_xuser),
                   .int_wr_resp_desc_6_xuser_5_xuser(int_wr_resp_desc_6_xuser_5_xuser),
                   .int_wr_resp_desc_6_xuser_6_xuser(int_wr_resp_desc_6_xuser_6_xuser),
                   .int_wr_resp_desc_6_xuser_7_xuser(int_wr_resp_desc_6_xuser_7_xuser),
                   .int_wr_resp_desc_6_xuser_8_xuser(int_wr_resp_desc_6_xuser_8_xuser),
                   .int_wr_resp_desc_6_xuser_9_xuser(int_wr_resp_desc_6_xuser_9_xuser),
                   .int_wr_resp_desc_6_xuser_10_xuser(int_wr_resp_desc_6_xuser_10_xuser),
                   .int_wr_resp_desc_6_xuser_11_xuser(int_wr_resp_desc_6_xuser_11_xuser),
                   .int_wr_resp_desc_6_xuser_12_xuser(int_wr_resp_desc_6_xuser_12_xuser),
                   .int_wr_resp_desc_6_xuser_13_xuser(int_wr_resp_desc_6_xuser_13_xuser),
                   .int_wr_resp_desc_6_xuser_14_xuser(int_wr_resp_desc_6_xuser_14_xuser),
                   .int_wr_resp_desc_6_xuser_15_xuser(int_wr_resp_desc_6_xuser_15_xuser),
                   .int_sn_req_desc_6_attr_acsnoop(int_sn_req_desc_6_attr_acsnoop),
                   .int_sn_req_desc_6_attr_acprot(int_sn_req_desc_6_attr_acprot),
                   .int_sn_req_desc_6_acaddr_0_addr(int_sn_req_desc_6_acaddr_0_addr),
                   .int_sn_req_desc_6_acaddr_1_addr(int_sn_req_desc_6_acaddr_1_addr),
                   .int_sn_req_desc_6_acaddr_2_addr(int_sn_req_desc_6_acaddr_2_addr),
                   .int_sn_req_desc_6_acaddr_3_addr(int_sn_req_desc_6_acaddr_3_addr),
                   .int_rd_resp_desc_7_data_offset_addr(int_rd_resp_desc_7_data_offset_addr),
                   .int_rd_resp_desc_7_data_size_size(int_rd_resp_desc_7_data_size_size),
                   .int_rd_resp_desc_7_data_host_addr_0_addr(int_rd_resp_desc_7_data_host_addr_0_addr),
                   .int_rd_resp_desc_7_data_host_addr_1_addr(int_rd_resp_desc_7_data_host_addr_1_addr),
                   .int_rd_resp_desc_7_data_host_addr_2_addr(int_rd_resp_desc_7_data_host_addr_2_addr),
                   .int_rd_resp_desc_7_data_host_addr_3_addr(int_rd_resp_desc_7_data_host_addr_3_addr),
                   .int_rd_resp_desc_7_resp_resp(int_rd_resp_desc_7_resp_resp),
                   .int_rd_resp_desc_7_xid_0_xid(int_rd_resp_desc_7_xid_0_xid),
                   .int_rd_resp_desc_7_xid_1_xid(int_rd_resp_desc_7_xid_1_xid),
                   .int_rd_resp_desc_7_xid_2_xid(int_rd_resp_desc_7_xid_2_xid),
                   .int_rd_resp_desc_7_xid_3_xid(int_rd_resp_desc_7_xid_3_xid),
                   .int_rd_resp_desc_7_xuser_0_xuser(int_rd_resp_desc_7_xuser_0_xuser),
                   .int_rd_resp_desc_7_xuser_1_xuser(int_rd_resp_desc_7_xuser_1_xuser),
                   .int_rd_resp_desc_7_xuser_2_xuser(int_rd_resp_desc_7_xuser_2_xuser),
                   .int_rd_resp_desc_7_xuser_3_xuser(int_rd_resp_desc_7_xuser_3_xuser),
                   .int_rd_resp_desc_7_xuser_4_xuser(int_rd_resp_desc_7_xuser_4_xuser),
                   .int_rd_resp_desc_7_xuser_5_xuser(int_rd_resp_desc_7_xuser_5_xuser),
                   .int_rd_resp_desc_7_xuser_6_xuser(int_rd_resp_desc_7_xuser_6_xuser),
                   .int_rd_resp_desc_7_xuser_7_xuser(int_rd_resp_desc_7_xuser_7_xuser),
                   .int_rd_resp_desc_7_xuser_8_xuser(int_rd_resp_desc_7_xuser_8_xuser),
                   .int_rd_resp_desc_7_xuser_9_xuser(int_rd_resp_desc_7_xuser_9_xuser),
                   .int_rd_resp_desc_7_xuser_10_xuser(int_rd_resp_desc_7_xuser_10_xuser),
                   .int_rd_resp_desc_7_xuser_11_xuser(int_rd_resp_desc_7_xuser_11_xuser),
                   .int_rd_resp_desc_7_xuser_12_xuser(int_rd_resp_desc_7_xuser_12_xuser),
                   .int_rd_resp_desc_7_xuser_13_xuser(int_rd_resp_desc_7_xuser_13_xuser),
                   .int_rd_resp_desc_7_xuser_14_xuser(int_rd_resp_desc_7_xuser_14_xuser),
                   .int_rd_resp_desc_7_xuser_15_xuser(int_rd_resp_desc_7_xuser_15_xuser),
                   .int_wr_req_desc_7_data_host_addr_0_addr(int_wr_req_desc_7_data_host_addr_0_addr),
                   .int_wr_req_desc_7_data_host_addr_1_addr(int_wr_req_desc_7_data_host_addr_1_addr),
                   .int_wr_req_desc_7_data_host_addr_2_addr(int_wr_req_desc_7_data_host_addr_2_addr),
                   .int_wr_req_desc_7_data_host_addr_3_addr(int_wr_req_desc_7_data_host_addr_3_addr),
                   .int_wr_req_desc_7_wstrb_host_addr_0_addr(int_wr_req_desc_7_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_7_wstrb_host_addr_1_addr(int_wr_req_desc_7_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_7_wstrb_host_addr_2_addr(int_wr_req_desc_7_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_7_wstrb_host_addr_3_addr(int_wr_req_desc_7_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_7_resp_resp(int_wr_resp_desc_7_resp_resp),
                   .int_wr_resp_desc_7_xid_0_xid(int_wr_resp_desc_7_xid_0_xid),
                   .int_wr_resp_desc_7_xid_1_xid(int_wr_resp_desc_7_xid_1_xid),
                   .int_wr_resp_desc_7_xid_2_xid(int_wr_resp_desc_7_xid_2_xid),
                   .int_wr_resp_desc_7_xid_3_xid(int_wr_resp_desc_7_xid_3_xid),
                   .int_wr_resp_desc_7_xuser_0_xuser(int_wr_resp_desc_7_xuser_0_xuser),
                   .int_wr_resp_desc_7_xuser_1_xuser(int_wr_resp_desc_7_xuser_1_xuser),
                   .int_wr_resp_desc_7_xuser_2_xuser(int_wr_resp_desc_7_xuser_2_xuser),
                   .int_wr_resp_desc_7_xuser_3_xuser(int_wr_resp_desc_7_xuser_3_xuser),
                   .int_wr_resp_desc_7_xuser_4_xuser(int_wr_resp_desc_7_xuser_4_xuser),
                   .int_wr_resp_desc_7_xuser_5_xuser(int_wr_resp_desc_7_xuser_5_xuser),
                   .int_wr_resp_desc_7_xuser_6_xuser(int_wr_resp_desc_7_xuser_6_xuser),
                   .int_wr_resp_desc_7_xuser_7_xuser(int_wr_resp_desc_7_xuser_7_xuser),
                   .int_wr_resp_desc_7_xuser_8_xuser(int_wr_resp_desc_7_xuser_8_xuser),
                   .int_wr_resp_desc_7_xuser_9_xuser(int_wr_resp_desc_7_xuser_9_xuser),
                   .int_wr_resp_desc_7_xuser_10_xuser(int_wr_resp_desc_7_xuser_10_xuser),
                   .int_wr_resp_desc_7_xuser_11_xuser(int_wr_resp_desc_7_xuser_11_xuser),
                   .int_wr_resp_desc_7_xuser_12_xuser(int_wr_resp_desc_7_xuser_12_xuser),
                   .int_wr_resp_desc_7_xuser_13_xuser(int_wr_resp_desc_7_xuser_13_xuser),
                   .int_wr_resp_desc_7_xuser_14_xuser(int_wr_resp_desc_7_xuser_14_xuser),
                   .int_wr_resp_desc_7_xuser_15_xuser(int_wr_resp_desc_7_xuser_15_xuser),
                   .int_sn_req_desc_7_attr_acsnoop(int_sn_req_desc_7_attr_acsnoop),
                   .int_sn_req_desc_7_attr_acprot(int_sn_req_desc_7_attr_acprot),
                   .int_sn_req_desc_7_acaddr_0_addr(int_sn_req_desc_7_acaddr_0_addr),
                   .int_sn_req_desc_7_acaddr_1_addr(int_sn_req_desc_7_acaddr_1_addr),
                   .int_sn_req_desc_7_acaddr_2_addr(int_sn_req_desc_7_acaddr_2_addr),
                   .int_sn_req_desc_7_acaddr_3_addr(int_sn_req_desc_7_acaddr_3_addr),
                   .int_rd_resp_desc_8_data_offset_addr(int_rd_resp_desc_8_data_offset_addr),
                   .int_rd_resp_desc_8_data_size_size(int_rd_resp_desc_8_data_size_size),
                   .int_rd_resp_desc_8_data_host_addr_0_addr(int_rd_resp_desc_8_data_host_addr_0_addr),
                   .int_rd_resp_desc_8_data_host_addr_1_addr(int_rd_resp_desc_8_data_host_addr_1_addr),
                   .int_rd_resp_desc_8_data_host_addr_2_addr(int_rd_resp_desc_8_data_host_addr_2_addr),
                   .int_rd_resp_desc_8_data_host_addr_3_addr(int_rd_resp_desc_8_data_host_addr_3_addr),
                   .int_rd_resp_desc_8_resp_resp(int_rd_resp_desc_8_resp_resp),
                   .int_rd_resp_desc_8_xid_0_xid(int_rd_resp_desc_8_xid_0_xid),
                   .int_rd_resp_desc_8_xid_1_xid(int_rd_resp_desc_8_xid_1_xid),
                   .int_rd_resp_desc_8_xid_2_xid(int_rd_resp_desc_8_xid_2_xid),
                   .int_rd_resp_desc_8_xid_3_xid(int_rd_resp_desc_8_xid_3_xid),
                   .int_rd_resp_desc_8_xuser_0_xuser(int_rd_resp_desc_8_xuser_0_xuser),
                   .int_rd_resp_desc_8_xuser_1_xuser(int_rd_resp_desc_8_xuser_1_xuser),
                   .int_rd_resp_desc_8_xuser_2_xuser(int_rd_resp_desc_8_xuser_2_xuser),
                   .int_rd_resp_desc_8_xuser_3_xuser(int_rd_resp_desc_8_xuser_3_xuser),
                   .int_rd_resp_desc_8_xuser_4_xuser(int_rd_resp_desc_8_xuser_4_xuser),
                   .int_rd_resp_desc_8_xuser_5_xuser(int_rd_resp_desc_8_xuser_5_xuser),
                   .int_rd_resp_desc_8_xuser_6_xuser(int_rd_resp_desc_8_xuser_6_xuser),
                   .int_rd_resp_desc_8_xuser_7_xuser(int_rd_resp_desc_8_xuser_7_xuser),
                   .int_rd_resp_desc_8_xuser_8_xuser(int_rd_resp_desc_8_xuser_8_xuser),
                   .int_rd_resp_desc_8_xuser_9_xuser(int_rd_resp_desc_8_xuser_9_xuser),
                   .int_rd_resp_desc_8_xuser_10_xuser(int_rd_resp_desc_8_xuser_10_xuser),
                   .int_rd_resp_desc_8_xuser_11_xuser(int_rd_resp_desc_8_xuser_11_xuser),
                   .int_rd_resp_desc_8_xuser_12_xuser(int_rd_resp_desc_8_xuser_12_xuser),
                   .int_rd_resp_desc_8_xuser_13_xuser(int_rd_resp_desc_8_xuser_13_xuser),
                   .int_rd_resp_desc_8_xuser_14_xuser(int_rd_resp_desc_8_xuser_14_xuser),
                   .int_rd_resp_desc_8_xuser_15_xuser(int_rd_resp_desc_8_xuser_15_xuser),
                   .int_wr_req_desc_8_data_host_addr_0_addr(int_wr_req_desc_8_data_host_addr_0_addr),
                   .int_wr_req_desc_8_data_host_addr_1_addr(int_wr_req_desc_8_data_host_addr_1_addr),
                   .int_wr_req_desc_8_data_host_addr_2_addr(int_wr_req_desc_8_data_host_addr_2_addr),
                   .int_wr_req_desc_8_data_host_addr_3_addr(int_wr_req_desc_8_data_host_addr_3_addr),
                   .int_wr_req_desc_8_wstrb_host_addr_0_addr(int_wr_req_desc_8_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_8_wstrb_host_addr_1_addr(int_wr_req_desc_8_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_8_wstrb_host_addr_2_addr(int_wr_req_desc_8_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_8_wstrb_host_addr_3_addr(int_wr_req_desc_8_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_8_resp_resp(int_wr_resp_desc_8_resp_resp),
                   .int_wr_resp_desc_8_xid_0_xid(int_wr_resp_desc_8_xid_0_xid),
                   .int_wr_resp_desc_8_xid_1_xid(int_wr_resp_desc_8_xid_1_xid),
                   .int_wr_resp_desc_8_xid_2_xid(int_wr_resp_desc_8_xid_2_xid),
                   .int_wr_resp_desc_8_xid_3_xid(int_wr_resp_desc_8_xid_3_xid),
                   .int_wr_resp_desc_8_xuser_0_xuser(int_wr_resp_desc_8_xuser_0_xuser),
                   .int_wr_resp_desc_8_xuser_1_xuser(int_wr_resp_desc_8_xuser_1_xuser),
                   .int_wr_resp_desc_8_xuser_2_xuser(int_wr_resp_desc_8_xuser_2_xuser),
                   .int_wr_resp_desc_8_xuser_3_xuser(int_wr_resp_desc_8_xuser_3_xuser),
                   .int_wr_resp_desc_8_xuser_4_xuser(int_wr_resp_desc_8_xuser_4_xuser),
                   .int_wr_resp_desc_8_xuser_5_xuser(int_wr_resp_desc_8_xuser_5_xuser),
                   .int_wr_resp_desc_8_xuser_6_xuser(int_wr_resp_desc_8_xuser_6_xuser),
                   .int_wr_resp_desc_8_xuser_7_xuser(int_wr_resp_desc_8_xuser_7_xuser),
                   .int_wr_resp_desc_8_xuser_8_xuser(int_wr_resp_desc_8_xuser_8_xuser),
                   .int_wr_resp_desc_8_xuser_9_xuser(int_wr_resp_desc_8_xuser_9_xuser),
                   .int_wr_resp_desc_8_xuser_10_xuser(int_wr_resp_desc_8_xuser_10_xuser),
                   .int_wr_resp_desc_8_xuser_11_xuser(int_wr_resp_desc_8_xuser_11_xuser),
                   .int_wr_resp_desc_8_xuser_12_xuser(int_wr_resp_desc_8_xuser_12_xuser),
                   .int_wr_resp_desc_8_xuser_13_xuser(int_wr_resp_desc_8_xuser_13_xuser),
                   .int_wr_resp_desc_8_xuser_14_xuser(int_wr_resp_desc_8_xuser_14_xuser),
                   .int_wr_resp_desc_8_xuser_15_xuser(int_wr_resp_desc_8_xuser_15_xuser),
                   .int_sn_req_desc_8_attr_acsnoop(int_sn_req_desc_8_attr_acsnoop),
                   .int_sn_req_desc_8_attr_acprot(int_sn_req_desc_8_attr_acprot),
                   .int_sn_req_desc_8_acaddr_0_addr(int_sn_req_desc_8_acaddr_0_addr),
                   .int_sn_req_desc_8_acaddr_1_addr(int_sn_req_desc_8_acaddr_1_addr),
                   .int_sn_req_desc_8_acaddr_2_addr(int_sn_req_desc_8_acaddr_2_addr),
                   .int_sn_req_desc_8_acaddr_3_addr(int_sn_req_desc_8_acaddr_3_addr),
                   .int_rd_resp_desc_9_data_offset_addr(int_rd_resp_desc_9_data_offset_addr),
                   .int_rd_resp_desc_9_data_size_size(int_rd_resp_desc_9_data_size_size),
                   .int_rd_resp_desc_9_data_host_addr_0_addr(int_rd_resp_desc_9_data_host_addr_0_addr),
                   .int_rd_resp_desc_9_data_host_addr_1_addr(int_rd_resp_desc_9_data_host_addr_1_addr),
                   .int_rd_resp_desc_9_data_host_addr_2_addr(int_rd_resp_desc_9_data_host_addr_2_addr),
                   .int_rd_resp_desc_9_data_host_addr_3_addr(int_rd_resp_desc_9_data_host_addr_3_addr),
                   .int_rd_resp_desc_9_resp_resp(int_rd_resp_desc_9_resp_resp),
                   .int_rd_resp_desc_9_xid_0_xid(int_rd_resp_desc_9_xid_0_xid),
                   .int_rd_resp_desc_9_xid_1_xid(int_rd_resp_desc_9_xid_1_xid),
                   .int_rd_resp_desc_9_xid_2_xid(int_rd_resp_desc_9_xid_2_xid),
                   .int_rd_resp_desc_9_xid_3_xid(int_rd_resp_desc_9_xid_3_xid),
                   .int_rd_resp_desc_9_xuser_0_xuser(int_rd_resp_desc_9_xuser_0_xuser),
                   .int_rd_resp_desc_9_xuser_1_xuser(int_rd_resp_desc_9_xuser_1_xuser),
                   .int_rd_resp_desc_9_xuser_2_xuser(int_rd_resp_desc_9_xuser_2_xuser),
                   .int_rd_resp_desc_9_xuser_3_xuser(int_rd_resp_desc_9_xuser_3_xuser),
                   .int_rd_resp_desc_9_xuser_4_xuser(int_rd_resp_desc_9_xuser_4_xuser),
                   .int_rd_resp_desc_9_xuser_5_xuser(int_rd_resp_desc_9_xuser_5_xuser),
                   .int_rd_resp_desc_9_xuser_6_xuser(int_rd_resp_desc_9_xuser_6_xuser),
                   .int_rd_resp_desc_9_xuser_7_xuser(int_rd_resp_desc_9_xuser_7_xuser),
                   .int_rd_resp_desc_9_xuser_8_xuser(int_rd_resp_desc_9_xuser_8_xuser),
                   .int_rd_resp_desc_9_xuser_9_xuser(int_rd_resp_desc_9_xuser_9_xuser),
                   .int_rd_resp_desc_9_xuser_10_xuser(int_rd_resp_desc_9_xuser_10_xuser),
                   .int_rd_resp_desc_9_xuser_11_xuser(int_rd_resp_desc_9_xuser_11_xuser),
                   .int_rd_resp_desc_9_xuser_12_xuser(int_rd_resp_desc_9_xuser_12_xuser),
                   .int_rd_resp_desc_9_xuser_13_xuser(int_rd_resp_desc_9_xuser_13_xuser),
                   .int_rd_resp_desc_9_xuser_14_xuser(int_rd_resp_desc_9_xuser_14_xuser),
                   .int_rd_resp_desc_9_xuser_15_xuser(int_rd_resp_desc_9_xuser_15_xuser),
                   .int_wr_req_desc_9_data_host_addr_0_addr(int_wr_req_desc_9_data_host_addr_0_addr),
                   .int_wr_req_desc_9_data_host_addr_1_addr(int_wr_req_desc_9_data_host_addr_1_addr),
                   .int_wr_req_desc_9_data_host_addr_2_addr(int_wr_req_desc_9_data_host_addr_2_addr),
                   .int_wr_req_desc_9_data_host_addr_3_addr(int_wr_req_desc_9_data_host_addr_3_addr),
                   .int_wr_req_desc_9_wstrb_host_addr_0_addr(int_wr_req_desc_9_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_9_wstrb_host_addr_1_addr(int_wr_req_desc_9_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_9_wstrb_host_addr_2_addr(int_wr_req_desc_9_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_9_wstrb_host_addr_3_addr(int_wr_req_desc_9_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_9_resp_resp(int_wr_resp_desc_9_resp_resp),
                   .int_wr_resp_desc_9_xid_0_xid(int_wr_resp_desc_9_xid_0_xid),
                   .int_wr_resp_desc_9_xid_1_xid(int_wr_resp_desc_9_xid_1_xid),
                   .int_wr_resp_desc_9_xid_2_xid(int_wr_resp_desc_9_xid_2_xid),
                   .int_wr_resp_desc_9_xid_3_xid(int_wr_resp_desc_9_xid_3_xid),
                   .int_wr_resp_desc_9_xuser_0_xuser(int_wr_resp_desc_9_xuser_0_xuser),
                   .int_wr_resp_desc_9_xuser_1_xuser(int_wr_resp_desc_9_xuser_1_xuser),
                   .int_wr_resp_desc_9_xuser_2_xuser(int_wr_resp_desc_9_xuser_2_xuser),
                   .int_wr_resp_desc_9_xuser_3_xuser(int_wr_resp_desc_9_xuser_3_xuser),
                   .int_wr_resp_desc_9_xuser_4_xuser(int_wr_resp_desc_9_xuser_4_xuser),
                   .int_wr_resp_desc_9_xuser_5_xuser(int_wr_resp_desc_9_xuser_5_xuser),
                   .int_wr_resp_desc_9_xuser_6_xuser(int_wr_resp_desc_9_xuser_6_xuser),
                   .int_wr_resp_desc_9_xuser_7_xuser(int_wr_resp_desc_9_xuser_7_xuser),
                   .int_wr_resp_desc_9_xuser_8_xuser(int_wr_resp_desc_9_xuser_8_xuser),
                   .int_wr_resp_desc_9_xuser_9_xuser(int_wr_resp_desc_9_xuser_9_xuser),
                   .int_wr_resp_desc_9_xuser_10_xuser(int_wr_resp_desc_9_xuser_10_xuser),
                   .int_wr_resp_desc_9_xuser_11_xuser(int_wr_resp_desc_9_xuser_11_xuser),
                   .int_wr_resp_desc_9_xuser_12_xuser(int_wr_resp_desc_9_xuser_12_xuser),
                   .int_wr_resp_desc_9_xuser_13_xuser(int_wr_resp_desc_9_xuser_13_xuser),
                   .int_wr_resp_desc_9_xuser_14_xuser(int_wr_resp_desc_9_xuser_14_xuser),
                   .int_wr_resp_desc_9_xuser_15_xuser(int_wr_resp_desc_9_xuser_15_xuser),
                   .int_sn_req_desc_9_attr_acsnoop(int_sn_req_desc_9_attr_acsnoop),
                   .int_sn_req_desc_9_attr_acprot(int_sn_req_desc_9_attr_acprot),
                   .int_sn_req_desc_9_acaddr_0_addr(int_sn_req_desc_9_acaddr_0_addr),
                   .int_sn_req_desc_9_acaddr_1_addr(int_sn_req_desc_9_acaddr_1_addr),
                   .int_sn_req_desc_9_acaddr_2_addr(int_sn_req_desc_9_acaddr_2_addr),
                   .int_sn_req_desc_9_acaddr_3_addr(int_sn_req_desc_9_acaddr_3_addr),
                   .int_rd_resp_desc_a_data_offset_addr(int_rd_resp_desc_a_data_offset_addr),
                   .int_rd_resp_desc_a_data_size_size(int_rd_resp_desc_a_data_size_size),
                   .int_rd_resp_desc_a_data_host_addr_0_addr(int_rd_resp_desc_a_data_host_addr_0_addr),
                   .int_rd_resp_desc_a_data_host_addr_1_addr(int_rd_resp_desc_a_data_host_addr_1_addr),
                   .int_rd_resp_desc_a_data_host_addr_2_addr(int_rd_resp_desc_a_data_host_addr_2_addr),
                   .int_rd_resp_desc_a_data_host_addr_3_addr(int_rd_resp_desc_a_data_host_addr_3_addr),
                   .int_rd_resp_desc_a_resp_resp(int_rd_resp_desc_a_resp_resp),
                   .int_rd_resp_desc_a_xid_0_xid(int_rd_resp_desc_a_xid_0_xid),
                   .int_rd_resp_desc_a_xid_1_xid(int_rd_resp_desc_a_xid_1_xid),
                   .int_rd_resp_desc_a_xid_2_xid(int_rd_resp_desc_a_xid_2_xid),
                   .int_rd_resp_desc_a_xid_3_xid(int_rd_resp_desc_a_xid_3_xid),
                   .int_rd_resp_desc_a_xuser_0_xuser(int_rd_resp_desc_a_xuser_0_xuser),
                   .int_rd_resp_desc_a_xuser_1_xuser(int_rd_resp_desc_a_xuser_1_xuser),
                   .int_rd_resp_desc_a_xuser_2_xuser(int_rd_resp_desc_a_xuser_2_xuser),
                   .int_rd_resp_desc_a_xuser_3_xuser(int_rd_resp_desc_a_xuser_3_xuser),
                   .int_rd_resp_desc_a_xuser_4_xuser(int_rd_resp_desc_a_xuser_4_xuser),
                   .int_rd_resp_desc_a_xuser_5_xuser(int_rd_resp_desc_a_xuser_5_xuser),
                   .int_rd_resp_desc_a_xuser_6_xuser(int_rd_resp_desc_a_xuser_6_xuser),
                   .int_rd_resp_desc_a_xuser_7_xuser(int_rd_resp_desc_a_xuser_7_xuser),
                   .int_rd_resp_desc_a_xuser_8_xuser(int_rd_resp_desc_a_xuser_8_xuser),
                   .int_rd_resp_desc_a_xuser_9_xuser(int_rd_resp_desc_a_xuser_9_xuser),
                   .int_rd_resp_desc_a_xuser_10_xuser(int_rd_resp_desc_a_xuser_10_xuser),
                   .int_rd_resp_desc_a_xuser_11_xuser(int_rd_resp_desc_a_xuser_11_xuser),
                   .int_rd_resp_desc_a_xuser_12_xuser(int_rd_resp_desc_a_xuser_12_xuser),
                   .int_rd_resp_desc_a_xuser_13_xuser(int_rd_resp_desc_a_xuser_13_xuser),
                   .int_rd_resp_desc_a_xuser_14_xuser(int_rd_resp_desc_a_xuser_14_xuser),
                   .int_rd_resp_desc_a_xuser_15_xuser(int_rd_resp_desc_a_xuser_15_xuser),
                   .int_wr_req_desc_a_data_host_addr_0_addr(int_wr_req_desc_a_data_host_addr_0_addr),
                   .int_wr_req_desc_a_data_host_addr_1_addr(int_wr_req_desc_a_data_host_addr_1_addr),
                   .int_wr_req_desc_a_data_host_addr_2_addr(int_wr_req_desc_a_data_host_addr_2_addr),
                   .int_wr_req_desc_a_data_host_addr_3_addr(int_wr_req_desc_a_data_host_addr_3_addr),
                   .int_wr_req_desc_a_wstrb_host_addr_0_addr(int_wr_req_desc_a_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_a_wstrb_host_addr_1_addr(int_wr_req_desc_a_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_a_wstrb_host_addr_2_addr(int_wr_req_desc_a_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_a_wstrb_host_addr_3_addr(int_wr_req_desc_a_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_a_resp_resp(int_wr_resp_desc_a_resp_resp),
                   .int_wr_resp_desc_a_xid_0_xid(int_wr_resp_desc_a_xid_0_xid),
                   .int_wr_resp_desc_a_xid_1_xid(int_wr_resp_desc_a_xid_1_xid),
                   .int_wr_resp_desc_a_xid_2_xid(int_wr_resp_desc_a_xid_2_xid),
                   .int_wr_resp_desc_a_xid_3_xid(int_wr_resp_desc_a_xid_3_xid),
                   .int_wr_resp_desc_a_xuser_0_xuser(int_wr_resp_desc_a_xuser_0_xuser),
                   .int_wr_resp_desc_a_xuser_1_xuser(int_wr_resp_desc_a_xuser_1_xuser),
                   .int_wr_resp_desc_a_xuser_2_xuser(int_wr_resp_desc_a_xuser_2_xuser),
                   .int_wr_resp_desc_a_xuser_3_xuser(int_wr_resp_desc_a_xuser_3_xuser),
                   .int_wr_resp_desc_a_xuser_4_xuser(int_wr_resp_desc_a_xuser_4_xuser),
                   .int_wr_resp_desc_a_xuser_5_xuser(int_wr_resp_desc_a_xuser_5_xuser),
                   .int_wr_resp_desc_a_xuser_6_xuser(int_wr_resp_desc_a_xuser_6_xuser),
                   .int_wr_resp_desc_a_xuser_7_xuser(int_wr_resp_desc_a_xuser_7_xuser),
                   .int_wr_resp_desc_a_xuser_8_xuser(int_wr_resp_desc_a_xuser_8_xuser),
                   .int_wr_resp_desc_a_xuser_9_xuser(int_wr_resp_desc_a_xuser_9_xuser),
                   .int_wr_resp_desc_a_xuser_10_xuser(int_wr_resp_desc_a_xuser_10_xuser),
                   .int_wr_resp_desc_a_xuser_11_xuser(int_wr_resp_desc_a_xuser_11_xuser),
                   .int_wr_resp_desc_a_xuser_12_xuser(int_wr_resp_desc_a_xuser_12_xuser),
                   .int_wr_resp_desc_a_xuser_13_xuser(int_wr_resp_desc_a_xuser_13_xuser),
                   .int_wr_resp_desc_a_xuser_14_xuser(int_wr_resp_desc_a_xuser_14_xuser),
                   .int_wr_resp_desc_a_xuser_15_xuser(int_wr_resp_desc_a_xuser_15_xuser),
                   .int_sn_req_desc_a_attr_acsnoop(int_sn_req_desc_a_attr_acsnoop),
                   .int_sn_req_desc_a_attr_acprot(int_sn_req_desc_a_attr_acprot),
                   .int_sn_req_desc_a_acaddr_0_addr(int_sn_req_desc_a_acaddr_0_addr),
                   .int_sn_req_desc_a_acaddr_1_addr(int_sn_req_desc_a_acaddr_1_addr),
                   .int_sn_req_desc_a_acaddr_2_addr(int_sn_req_desc_a_acaddr_2_addr),
                   .int_sn_req_desc_a_acaddr_3_addr(int_sn_req_desc_a_acaddr_3_addr),
                   .int_rd_resp_desc_b_data_offset_addr(int_rd_resp_desc_b_data_offset_addr),
                   .int_rd_resp_desc_b_data_size_size(int_rd_resp_desc_b_data_size_size),
                   .int_rd_resp_desc_b_data_host_addr_0_addr(int_rd_resp_desc_b_data_host_addr_0_addr),
                   .int_rd_resp_desc_b_data_host_addr_1_addr(int_rd_resp_desc_b_data_host_addr_1_addr),
                   .int_rd_resp_desc_b_data_host_addr_2_addr(int_rd_resp_desc_b_data_host_addr_2_addr),
                   .int_rd_resp_desc_b_data_host_addr_3_addr(int_rd_resp_desc_b_data_host_addr_3_addr),
                   .int_rd_resp_desc_b_resp_resp(int_rd_resp_desc_b_resp_resp),
                   .int_rd_resp_desc_b_xid_0_xid(int_rd_resp_desc_b_xid_0_xid),
                   .int_rd_resp_desc_b_xid_1_xid(int_rd_resp_desc_b_xid_1_xid),
                   .int_rd_resp_desc_b_xid_2_xid(int_rd_resp_desc_b_xid_2_xid),
                   .int_rd_resp_desc_b_xid_3_xid(int_rd_resp_desc_b_xid_3_xid),
                   .int_rd_resp_desc_b_xuser_0_xuser(int_rd_resp_desc_b_xuser_0_xuser),
                   .int_rd_resp_desc_b_xuser_1_xuser(int_rd_resp_desc_b_xuser_1_xuser),
                   .int_rd_resp_desc_b_xuser_2_xuser(int_rd_resp_desc_b_xuser_2_xuser),
                   .int_rd_resp_desc_b_xuser_3_xuser(int_rd_resp_desc_b_xuser_3_xuser),
                   .int_rd_resp_desc_b_xuser_4_xuser(int_rd_resp_desc_b_xuser_4_xuser),
                   .int_rd_resp_desc_b_xuser_5_xuser(int_rd_resp_desc_b_xuser_5_xuser),
                   .int_rd_resp_desc_b_xuser_6_xuser(int_rd_resp_desc_b_xuser_6_xuser),
                   .int_rd_resp_desc_b_xuser_7_xuser(int_rd_resp_desc_b_xuser_7_xuser),
                   .int_rd_resp_desc_b_xuser_8_xuser(int_rd_resp_desc_b_xuser_8_xuser),
                   .int_rd_resp_desc_b_xuser_9_xuser(int_rd_resp_desc_b_xuser_9_xuser),
                   .int_rd_resp_desc_b_xuser_10_xuser(int_rd_resp_desc_b_xuser_10_xuser),
                   .int_rd_resp_desc_b_xuser_11_xuser(int_rd_resp_desc_b_xuser_11_xuser),
                   .int_rd_resp_desc_b_xuser_12_xuser(int_rd_resp_desc_b_xuser_12_xuser),
                   .int_rd_resp_desc_b_xuser_13_xuser(int_rd_resp_desc_b_xuser_13_xuser),
                   .int_rd_resp_desc_b_xuser_14_xuser(int_rd_resp_desc_b_xuser_14_xuser),
                   .int_rd_resp_desc_b_xuser_15_xuser(int_rd_resp_desc_b_xuser_15_xuser),
                   .int_wr_req_desc_b_data_host_addr_0_addr(int_wr_req_desc_b_data_host_addr_0_addr),
                   .int_wr_req_desc_b_data_host_addr_1_addr(int_wr_req_desc_b_data_host_addr_1_addr),
                   .int_wr_req_desc_b_data_host_addr_2_addr(int_wr_req_desc_b_data_host_addr_2_addr),
                   .int_wr_req_desc_b_data_host_addr_3_addr(int_wr_req_desc_b_data_host_addr_3_addr),
                   .int_wr_req_desc_b_wstrb_host_addr_0_addr(int_wr_req_desc_b_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_b_wstrb_host_addr_1_addr(int_wr_req_desc_b_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_b_wstrb_host_addr_2_addr(int_wr_req_desc_b_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_b_wstrb_host_addr_3_addr(int_wr_req_desc_b_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_b_resp_resp(int_wr_resp_desc_b_resp_resp),
                   .int_wr_resp_desc_b_xid_0_xid(int_wr_resp_desc_b_xid_0_xid),
                   .int_wr_resp_desc_b_xid_1_xid(int_wr_resp_desc_b_xid_1_xid),
                   .int_wr_resp_desc_b_xid_2_xid(int_wr_resp_desc_b_xid_2_xid),
                   .int_wr_resp_desc_b_xid_3_xid(int_wr_resp_desc_b_xid_3_xid),
                   .int_wr_resp_desc_b_xuser_0_xuser(int_wr_resp_desc_b_xuser_0_xuser),
                   .int_wr_resp_desc_b_xuser_1_xuser(int_wr_resp_desc_b_xuser_1_xuser),
                   .int_wr_resp_desc_b_xuser_2_xuser(int_wr_resp_desc_b_xuser_2_xuser),
                   .int_wr_resp_desc_b_xuser_3_xuser(int_wr_resp_desc_b_xuser_3_xuser),
                   .int_wr_resp_desc_b_xuser_4_xuser(int_wr_resp_desc_b_xuser_4_xuser),
                   .int_wr_resp_desc_b_xuser_5_xuser(int_wr_resp_desc_b_xuser_5_xuser),
                   .int_wr_resp_desc_b_xuser_6_xuser(int_wr_resp_desc_b_xuser_6_xuser),
                   .int_wr_resp_desc_b_xuser_7_xuser(int_wr_resp_desc_b_xuser_7_xuser),
                   .int_wr_resp_desc_b_xuser_8_xuser(int_wr_resp_desc_b_xuser_8_xuser),
                   .int_wr_resp_desc_b_xuser_9_xuser(int_wr_resp_desc_b_xuser_9_xuser),
                   .int_wr_resp_desc_b_xuser_10_xuser(int_wr_resp_desc_b_xuser_10_xuser),
                   .int_wr_resp_desc_b_xuser_11_xuser(int_wr_resp_desc_b_xuser_11_xuser),
                   .int_wr_resp_desc_b_xuser_12_xuser(int_wr_resp_desc_b_xuser_12_xuser),
                   .int_wr_resp_desc_b_xuser_13_xuser(int_wr_resp_desc_b_xuser_13_xuser),
                   .int_wr_resp_desc_b_xuser_14_xuser(int_wr_resp_desc_b_xuser_14_xuser),
                   .int_wr_resp_desc_b_xuser_15_xuser(int_wr_resp_desc_b_xuser_15_xuser),
                   .int_sn_req_desc_b_attr_acsnoop(int_sn_req_desc_b_attr_acsnoop),
                   .int_sn_req_desc_b_attr_acprot(int_sn_req_desc_b_attr_acprot),
                   .int_sn_req_desc_b_acaddr_0_addr(int_sn_req_desc_b_acaddr_0_addr),
                   .int_sn_req_desc_b_acaddr_1_addr(int_sn_req_desc_b_acaddr_1_addr),
                   .int_sn_req_desc_b_acaddr_2_addr(int_sn_req_desc_b_acaddr_2_addr),
                   .int_sn_req_desc_b_acaddr_3_addr(int_sn_req_desc_b_acaddr_3_addr),
                   .int_rd_resp_desc_c_data_offset_addr(int_rd_resp_desc_c_data_offset_addr),
                   .int_rd_resp_desc_c_data_size_size(int_rd_resp_desc_c_data_size_size),
                   .int_rd_resp_desc_c_data_host_addr_0_addr(int_rd_resp_desc_c_data_host_addr_0_addr),
                   .int_rd_resp_desc_c_data_host_addr_1_addr(int_rd_resp_desc_c_data_host_addr_1_addr),
                   .int_rd_resp_desc_c_data_host_addr_2_addr(int_rd_resp_desc_c_data_host_addr_2_addr),
                   .int_rd_resp_desc_c_data_host_addr_3_addr(int_rd_resp_desc_c_data_host_addr_3_addr),
                   .int_rd_resp_desc_c_resp_resp(int_rd_resp_desc_c_resp_resp),
                   .int_rd_resp_desc_c_xid_0_xid(int_rd_resp_desc_c_xid_0_xid),
                   .int_rd_resp_desc_c_xid_1_xid(int_rd_resp_desc_c_xid_1_xid),
                   .int_rd_resp_desc_c_xid_2_xid(int_rd_resp_desc_c_xid_2_xid),
                   .int_rd_resp_desc_c_xid_3_xid(int_rd_resp_desc_c_xid_3_xid),
                   .int_rd_resp_desc_c_xuser_0_xuser(int_rd_resp_desc_c_xuser_0_xuser),
                   .int_rd_resp_desc_c_xuser_1_xuser(int_rd_resp_desc_c_xuser_1_xuser),
                   .int_rd_resp_desc_c_xuser_2_xuser(int_rd_resp_desc_c_xuser_2_xuser),
                   .int_rd_resp_desc_c_xuser_3_xuser(int_rd_resp_desc_c_xuser_3_xuser),
                   .int_rd_resp_desc_c_xuser_4_xuser(int_rd_resp_desc_c_xuser_4_xuser),
                   .int_rd_resp_desc_c_xuser_5_xuser(int_rd_resp_desc_c_xuser_5_xuser),
                   .int_rd_resp_desc_c_xuser_6_xuser(int_rd_resp_desc_c_xuser_6_xuser),
                   .int_rd_resp_desc_c_xuser_7_xuser(int_rd_resp_desc_c_xuser_7_xuser),
                   .int_rd_resp_desc_c_xuser_8_xuser(int_rd_resp_desc_c_xuser_8_xuser),
                   .int_rd_resp_desc_c_xuser_9_xuser(int_rd_resp_desc_c_xuser_9_xuser),
                   .int_rd_resp_desc_c_xuser_10_xuser(int_rd_resp_desc_c_xuser_10_xuser),
                   .int_rd_resp_desc_c_xuser_11_xuser(int_rd_resp_desc_c_xuser_11_xuser),
                   .int_rd_resp_desc_c_xuser_12_xuser(int_rd_resp_desc_c_xuser_12_xuser),
                   .int_rd_resp_desc_c_xuser_13_xuser(int_rd_resp_desc_c_xuser_13_xuser),
                   .int_rd_resp_desc_c_xuser_14_xuser(int_rd_resp_desc_c_xuser_14_xuser),
                   .int_rd_resp_desc_c_xuser_15_xuser(int_rd_resp_desc_c_xuser_15_xuser),
                   .int_wr_req_desc_c_data_host_addr_0_addr(int_wr_req_desc_c_data_host_addr_0_addr),
                   .int_wr_req_desc_c_data_host_addr_1_addr(int_wr_req_desc_c_data_host_addr_1_addr),
                   .int_wr_req_desc_c_data_host_addr_2_addr(int_wr_req_desc_c_data_host_addr_2_addr),
                   .int_wr_req_desc_c_data_host_addr_3_addr(int_wr_req_desc_c_data_host_addr_3_addr),
                   .int_wr_req_desc_c_wstrb_host_addr_0_addr(int_wr_req_desc_c_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_c_wstrb_host_addr_1_addr(int_wr_req_desc_c_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_c_wstrb_host_addr_2_addr(int_wr_req_desc_c_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_c_wstrb_host_addr_3_addr(int_wr_req_desc_c_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_c_resp_resp(int_wr_resp_desc_c_resp_resp),
                   .int_wr_resp_desc_c_xid_0_xid(int_wr_resp_desc_c_xid_0_xid),
                   .int_wr_resp_desc_c_xid_1_xid(int_wr_resp_desc_c_xid_1_xid),
                   .int_wr_resp_desc_c_xid_2_xid(int_wr_resp_desc_c_xid_2_xid),
                   .int_wr_resp_desc_c_xid_3_xid(int_wr_resp_desc_c_xid_3_xid),
                   .int_wr_resp_desc_c_xuser_0_xuser(int_wr_resp_desc_c_xuser_0_xuser),
                   .int_wr_resp_desc_c_xuser_1_xuser(int_wr_resp_desc_c_xuser_1_xuser),
                   .int_wr_resp_desc_c_xuser_2_xuser(int_wr_resp_desc_c_xuser_2_xuser),
                   .int_wr_resp_desc_c_xuser_3_xuser(int_wr_resp_desc_c_xuser_3_xuser),
                   .int_wr_resp_desc_c_xuser_4_xuser(int_wr_resp_desc_c_xuser_4_xuser),
                   .int_wr_resp_desc_c_xuser_5_xuser(int_wr_resp_desc_c_xuser_5_xuser),
                   .int_wr_resp_desc_c_xuser_6_xuser(int_wr_resp_desc_c_xuser_6_xuser),
                   .int_wr_resp_desc_c_xuser_7_xuser(int_wr_resp_desc_c_xuser_7_xuser),
                   .int_wr_resp_desc_c_xuser_8_xuser(int_wr_resp_desc_c_xuser_8_xuser),
                   .int_wr_resp_desc_c_xuser_9_xuser(int_wr_resp_desc_c_xuser_9_xuser),
                   .int_wr_resp_desc_c_xuser_10_xuser(int_wr_resp_desc_c_xuser_10_xuser),
                   .int_wr_resp_desc_c_xuser_11_xuser(int_wr_resp_desc_c_xuser_11_xuser),
                   .int_wr_resp_desc_c_xuser_12_xuser(int_wr_resp_desc_c_xuser_12_xuser),
                   .int_wr_resp_desc_c_xuser_13_xuser(int_wr_resp_desc_c_xuser_13_xuser),
                   .int_wr_resp_desc_c_xuser_14_xuser(int_wr_resp_desc_c_xuser_14_xuser),
                   .int_wr_resp_desc_c_xuser_15_xuser(int_wr_resp_desc_c_xuser_15_xuser),
                   .int_sn_req_desc_c_attr_acsnoop(int_sn_req_desc_c_attr_acsnoop),
                   .int_sn_req_desc_c_attr_acprot(int_sn_req_desc_c_attr_acprot),
                   .int_sn_req_desc_c_acaddr_0_addr(int_sn_req_desc_c_acaddr_0_addr),
                   .int_sn_req_desc_c_acaddr_1_addr(int_sn_req_desc_c_acaddr_1_addr),
                   .int_sn_req_desc_c_acaddr_2_addr(int_sn_req_desc_c_acaddr_2_addr),
                   .int_sn_req_desc_c_acaddr_3_addr(int_sn_req_desc_c_acaddr_3_addr),
                   .int_rd_resp_desc_d_data_offset_addr(int_rd_resp_desc_d_data_offset_addr),
                   .int_rd_resp_desc_d_data_size_size(int_rd_resp_desc_d_data_size_size),
                   .int_rd_resp_desc_d_data_host_addr_0_addr(int_rd_resp_desc_d_data_host_addr_0_addr),
                   .int_rd_resp_desc_d_data_host_addr_1_addr(int_rd_resp_desc_d_data_host_addr_1_addr),
                   .int_rd_resp_desc_d_data_host_addr_2_addr(int_rd_resp_desc_d_data_host_addr_2_addr),
                   .int_rd_resp_desc_d_data_host_addr_3_addr(int_rd_resp_desc_d_data_host_addr_3_addr),
                   .int_rd_resp_desc_d_resp_resp(int_rd_resp_desc_d_resp_resp),
                   .int_rd_resp_desc_d_xid_0_xid(int_rd_resp_desc_d_xid_0_xid),
                   .int_rd_resp_desc_d_xid_1_xid(int_rd_resp_desc_d_xid_1_xid),
                   .int_rd_resp_desc_d_xid_2_xid(int_rd_resp_desc_d_xid_2_xid),
                   .int_rd_resp_desc_d_xid_3_xid(int_rd_resp_desc_d_xid_3_xid),
                   .int_rd_resp_desc_d_xuser_0_xuser(int_rd_resp_desc_d_xuser_0_xuser),
                   .int_rd_resp_desc_d_xuser_1_xuser(int_rd_resp_desc_d_xuser_1_xuser),
                   .int_rd_resp_desc_d_xuser_2_xuser(int_rd_resp_desc_d_xuser_2_xuser),
                   .int_rd_resp_desc_d_xuser_3_xuser(int_rd_resp_desc_d_xuser_3_xuser),
                   .int_rd_resp_desc_d_xuser_4_xuser(int_rd_resp_desc_d_xuser_4_xuser),
                   .int_rd_resp_desc_d_xuser_5_xuser(int_rd_resp_desc_d_xuser_5_xuser),
                   .int_rd_resp_desc_d_xuser_6_xuser(int_rd_resp_desc_d_xuser_6_xuser),
                   .int_rd_resp_desc_d_xuser_7_xuser(int_rd_resp_desc_d_xuser_7_xuser),
                   .int_rd_resp_desc_d_xuser_8_xuser(int_rd_resp_desc_d_xuser_8_xuser),
                   .int_rd_resp_desc_d_xuser_9_xuser(int_rd_resp_desc_d_xuser_9_xuser),
                   .int_rd_resp_desc_d_xuser_10_xuser(int_rd_resp_desc_d_xuser_10_xuser),
                   .int_rd_resp_desc_d_xuser_11_xuser(int_rd_resp_desc_d_xuser_11_xuser),
                   .int_rd_resp_desc_d_xuser_12_xuser(int_rd_resp_desc_d_xuser_12_xuser),
                   .int_rd_resp_desc_d_xuser_13_xuser(int_rd_resp_desc_d_xuser_13_xuser),
                   .int_rd_resp_desc_d_xuser_14_xuser(int_rd_resp_desc_d_xuser_14_xuser),
                   .int_rd_resp_desc_d_xuser_15_xuser(int_rd_resp_desc_d_xuser_15_xuser),
                   .int_wr_req_desc_d_data_host_addr_0_addr(int_wr_req_desc_d_data_host_addr_0_addr),
                   .int_wr_req_desc_d_data_host_addr_1_addr(int_wr_req_desc_d_data_host_addr_1_addr),
                   .int_wr_req_desc_d_data_host_addr_2_addr(int_wr_req_desc_d_data_host_addr_2_addr),
                   .int_wr_req_desc_d_data_host_addr_3_addr(int_wr_req_desc_d_data_host_addr_3_addr),
                   .int_wr_req_desc_d_wstrb_host_addr_0_addr(int_wr_req_desc_d_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_d_wstrb_host_addr_1_addr(int_wr_req_desc_d_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_d_wstrb_host_addr_2_addr(int_wr_req_desc_d_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_d_wstrb_host_addr_3_addr(int_wr_req_desc_d_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_d_resp_resp(int_wr_resp_desc_d_resp_resp),
                   .int_wr_resp_desc_d_xid_0_xid(int_wr_resp_desc_d_xid_0_xid),
                   .int_wr_resp_desc_d_xid_1_xid(int_wr_resp_desc_d_xid_1_xid),
                   .int_wr_resp_desc_d_xid_2_xid(int_wr_resp_desc_d_xid_2_xid),
                   .int_wr_resp_desc_d_xid_3_xid(int_wr_resp_desc_d_xid_3_xid),
                   .int_wr_resp_desc_d_xuser_0_xuser(int_wr_resp_desc_d_xuser_0_xuser),
                   .int_wr_resp_desc_d_xuser_1_xuser(int_wr_resp_desc_d_xuser_1_xuser),
                   .int_wr_resp_desc_d_xuser_2_xuser(int_wr_resp_desc_d_xuser_2_xuser),
                   .int_wr_resp_desc_d_xuser_3_xuser(int_wr_resp_desc_d_xuser_3_xuser),
                   .int_wr_resp_desc_d_xuser_4_xuser(int_wr_resp_desc_d_xuser_4_xuser),
                   .int_wr_resp_desc_d_xuser_5_xuser(int_wr_resp_desc_d_xuser_5_xuser),
                   .int_wr_resp_desc_d_xuser_6_xuser(int_wr_resp_desc_d_xuser_6_xuser),
                   .int_wr_resp_desc_d_xuser_7_xuser(int_wr_resp_desc_d_xuser_7_xuser),
                   .int_wr_resp_desc_d_xuser_8_xuser(int_wr_resp_desc_d_xuser_8_xuser),
                   .int_wr_resp_desc_d_xuser_9_xuser(int_wr_resp_desc_d_xuser_9_xuser),
                   .int_wr_resp_desc_d_xuser_10_xuser(int_wr_resp_desc_d_xuser_10_xuser),
                   .int_wr_resp_desc_d_xuser_11_xuser(int_wr_resp_desc_d_xuser_11_xuser),
                   .int_wr_resp_desc_d_xuser_12_xuser(int_wr_resp_desc_d_xuser_12_xuser),
                   .int_wr_resp_desc_d_xuser_13_xuser(int_wr_resp_desc_d_xuser_13_xuser),
                   .int_wr_resp_desc_d_xuser_14_xuser(int_wr_resp_desc_d_xuser_14_xuser),
                   .int_wr_resp_desc_d_xuser_15_xuser(int_wr_resp_desc_d_xuser_15_xuser),
                   .int_sn_req_desc_d_attr_acsnoop(int_sn_req_desc_d_attr_acsnoop),
                   .int_sn_req_desc_d_attr_acprot(int_sn_req_desc_d_attr_acprot),
                   .int_sn_req_desc_d_acaddr_0_addr(int_sn_req_desc_d_acaddr_0_addr),
                   .int_sn_req_desc_d_acaddr_1_addr(int_sn_req_desc_d_acaddr_1_addr),
                   .int_sn_req_desc_d_acaddr_2_addr(int_sn_req_desc_d_acaddr_2_addr),
                   .int_sn_req_desc_d_acaddr_3_addr(int_sn_req_desc_d_acaddr_3_addr),
                   .int_rd_resp_desc_e_data_offset_addr(int_rd_resp_desc_e_data_offset_addr),
                   .int_rd_resp_desc_e_data_size_size(int_rd_resp_desc_e_data_size_size),
                   .int_rd_resp_desc_e_data_host_addr_0_addr(int_rd_resp_desc_e_data_host_addr_0_addr),
                   .int_rd_resp_desc_e_data_host_addr_1_addr(int_rd_resp_desc_e_data_host_addr_1_addr),
                   .int_rd_resp_desc_e_data_host_addr_2_addr(int_rd_resp_desc_e_data_host_addr_2_addr),
                   .int_rd_resp_desc_e_data_host_addr_3_addr(int_rd_resp_desc_e_data_host_addr_3_addr),
                   .int_rd_resp_desc_e_resp_resp(int_rd_resp_desc_e_resp_resp),
                   .int_rd_resp_desc_e_xid_0_xid(int_rd_resp_desc_e_xid_0_xid),
                   .int_rd_resp_desc_e_xid_1_xid(int_rd_resp_desc_e_xid_1_xid),
                   .int_rd_resp_desc_e_xid_2_xid(int_rd_resp_desc_e_xid_2_xid),
                   .int_rd_resp_desc_e_xid_3_xid(int_rd_resp_desc_e_xid_3_xid),
                   .int_rd_resp_desc_e_xuser_0_xuser(int_rd_resp_desc_e_xuser_0_xuser),
                   .int_rd_resp_desc_e_xuser_1_xuser(int_rd_resp_desc_e_xuser_1_xuser),
                   .int_rd_resp_desc_e_xuser_2_xuser(int_rd_resp_desc_e_xuser_2_xuser),
                   .int_rd_resp_desc_e_xuser_3_xuser(int_rd_resp_desc_e_xuser_3_xuser),
                   .int_rd_resp_desc_e_xuser_4_xuser(int_rd_resp_desc_e_xuser_4_xuser),
                   .int_rd_resp_desc_e_xuser_5_xuser(int_rd_resp_desc_e_xuser_5_xuser),
                   .int_rd_resp_desc_e_xuser_6_xuser(int_rd_resp_desc_e_xuser_6_xuser),
                   .int_rd_resp_desc_e_xuser_7_xuser(int_rd_resp_desc_e_xuser_7_xuser),
                   .int_rd_resp_desc_e_xuser_8_xuser(int_rd_resp_desc_e_xuser_8_xuser),
                   .int_rd_resp_desc_e_xuser_9_xuser(int_rd_resp_desc_e_xuser_9_xuser),
                   .int_rd_resp_desc_e_xuser_10_xuser(int_rd_resp_desc_e_xuser_10_xuser),
                   .int_rd_resp_desc_e_xuser_11_xuser(int_rd_resp_desc_e_xuser_11_xuser),
                   .int_rd_resp_desc_e_xuser_12_xuser(int_rd_resp_desc_e_xuser_12_xuser),
                   .int_rd_resp_desc_e_xuser_13_xuser(int_rd_resp_desc_e_xuser_13_xuser),
                   .int_rd_resp_desc_e_xuser_14_xuser(int_rd_resp_desc_e_xuser_14_xuser),
                   .int_rd_resp_desc_e_xuser_15_xuser(int_rd_resp_desc_e_xuser_15_xuser),
                   .int_wr_req_desc_e_data_host_addr_0_addr(int_wr_req_desc_e_data_host_addr_0_addr),
                   .int_wr_req_desc_e_data_host_addr_1_addr(int_wr_req_desc_e_data_host_addr_1_addr),
                   .int_wr_req_desc_e_data_host_addr_2_addr(int_wr_req_desc_e_data_host_addr_2_addr),
                   .int_wr_req_desc_e_data_host_addr_3_addr(int_wr_req_desc_e_data_host_addr_3_addr),
                   .int_wr_req_desc_e_wstrb_host_addr_0_addr(int_wr_req_desc_e_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_e_wstrb_host_addr_1_addr(int_wr_req_desc_e_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_e_wstrb_host_addr_2_addr(int_wr_req_desc_e_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_e_wstrb_host_addr_3_addr(int_wr_req_desc_e_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_e_resp_resp(int_wr_resp_desc_e_resp_resp),
                   .int_wr_resp_desc_e_xid_0_xid(int_wr_resp_desc_e_xid_0_xid),
                   .int_wr_resp_desc_e_xid_1_xid(int_wr_resp_desc_e_xid_1_xid),
                   .int_wr_resp_desc_e_xid_2_xid(int_wr_resp_desc_e_xid_2_xid),
                   .int_wr_resp_desc_e_xid_3_xid(int_wr_resp_desc_e_xid_3_xid),
                   .int_wr_resp_desc_e_xuser_0_xuser(int_wr_resp_desc_e_xuser_0_xuser),
                   .int_wr_resp_desc_e_xuser_1_xuser(int_wr_resp_desc_e_xuser_1_xuser),
                   .int_wr_resp_desc_e_xuser_2_xuser(int_wr_resp_desc_e_xuser_2_xuser),
                   .int_wr_resp_desc_e_xuser_3_xuser(int_wr_resp_desc_e_xuser_3_xuser),
                   .int_wr_resp_desc_e_xuser_4_xuser(int_wr_resp_desc_e_xuser_4_xuser),
                   .int_wr_resp_desc_e_xuser_5_xuser(int_wr_resp_desc_e_xuser_5_xuser),
                   .int_wr_resp_desc_e_xuser_6_xuser(int_wr_resp_desc_e_xuser_6_xuser),
                   .int_wr_resp_desc_e_xuser_7_xuser(int_wr_resp_desc_e_xuser_7_xuser),
                   .int_wr_resp_desc_e_xuser_8_xuser(int_wr_resp_desc_e_xuser_8_xuser),
                   .int_wr_resp_desc_e_xuser_9_xuser(int_wr_resp_desc_e_xuser_9_xuser),
                   .int_wr_resp_desc_e_xuser_10_xuser(int_wr_resp_desc_e_xuser_10_xuser),
                   .int_wr_resp_desc_e_xuser_11_xuser(int_wr_resp_desc_e_xuser_11_xuser),
                   .int_wr_resp_desc_e_xuser_12_xuser(int_wr_resp_desc_e_xuser_12_xuser),
                   .int_wr_resp_desc_e_xuser_13_xuser(int_wr_resp_desc_e_xuser_13_xuser),
                   .int_wr_resp_desc_e_xuser_14_xuser(int_wr_resp_desc_e_xuser_14_xuser),
                   .int_wr_resp_desc_e_xuser_15_xuser(int_wr_resp_desc_e_xuser_15_xuser),
                   .int_sn_req_desc_e_attr_acsnoop(int_sn_req_desc_e_attr_acsnoop),
                   .int_sn_req_desc_e_attr_acprot(int_sn_req_desc_e_attr_acprot),
                   .int_sn_req_desc_e_acaddr_0_addr(int_sn_req_desc_e_acaddr_0_addr),
                   .int_sn_req_desc_e_acaddr_1_addr(int_sn_req_desc_e_acaddr_1_addr),
                   .int_sn_req_desc_e_acaddr_2_addr(int_sn_req_desc_e_acaddr_2_addr),
                   .int_sn_req_desc_e_acaddr_3_addr(int_sn_req_desc_e_acaddr_3_addr),
                   .int_rd_resp_desc_f_data_offset_addr(int_rd_resp_desc_f_data_offset_addr),
                   .int_rd_resp_desc_f_data_size_size(int_rd_resp_desc_f_data_size_size),
                   .int_rd_resp_desc_f_data_host_addr_0_addr(int_rd_resp_desc_f_data_host_addr_0_addr),
                   .int_rd_resp_desc_f_data_host_addr_1_addr(int_rd_resp_desc_f_data_host_addr_1_addr),
                   .int_rd_resp_desc_f_data_host_addr_2_addr(int_rd_resp_desc_f_data_host_addr_2_addr),
                   .int_rd_resp_desc_f_data_host_addr_3_addr(int_rd_resp_desc_f_data_host_addr_3_addr),
                   .int_rd_resp_desc_f_resp_resp(int_rd_resp_desc_f_resp_resp),
                   .int_rd_resp_desc_f_xid_0_xid(int_rd_resp_desc_f_xid_0_xid),
                   .int_rd_resp_desc_f_xid_1_xid(int_rd_resp_desc_f_xid_1_xid),
                   .int_rd_resp_desc_f_xid_2_xid(int_rd_resp_desc_f_xid_2_xid),
                   .int_rd_resp_desc_f_xid_3_xid(int_rd_resp_desc_f_xid_3_xid),
                   .int_rd_resp_desc_f_xuser_0_xuser(int_rd_resp_desc_f_xuser_0_xuser),
                   .int_rd_resp_desc_f_xuser_1_xuser(int_rd_resp_desc_f_xuser_1_xuser),
                   .int_rd_resp_desc_f_xuser_2_xuser(int_rd_resp_desc_f_xuser_2_xuser),
                   .int_rd_resp_desc_f_xuser_3_xuser(int_rd_resp_desc_f_xuser_3_xuser),
                   .int_rd_resp_desc_f_xuser_4_xuser(int_rd_resp_desc_f_xuser_4_xuser),
                   .int_rd_resp_desc_f_xuser_5_xuser(int_rd_resp_desc_f_xuser_5_xuser),
                   .int_rd_resp_desc_f_xuser_6_xuser(int_rd_resp_desc_f_xuser_6_xuser),
                   .int_rd_resp_desc_f_xuser_7_xuser(int_rd_resp_desc_f_xuser_7_xuser),
                   .int_rd_resp_desc_f_xuser_8_xuser(int_rd_resp_desc_f_xuser_8_xuser),
                   .int_rd_resp_desc_f_xuser_9_xuser(int_rd_resp_desc_f_xuser_9_xuser),
                   .int_rd_resp_desc_f_xuser_10_xuser(int_rd_resp_desc_f_xuser_10_xuser),
                   .int_rd_resp_desc_f_xuser_11_xuser(int_rd_resp_desc_f_xuser_11_xuser),
                   .int_rd_resp_desc_f_xuser_12_xuser(int_rd_resp_desc_f_xuser_12_xuser),
                   .int_rd_resp_desc_f_xuser_13_xuser(int_rd_resp_desc_f_xuser_13_xuser),
                   .int_rd_resp_desc_f_xuser_14_xuser(int_rd_resp_desc_f_xuser_14_xuser),
                   .int_rd_resp_desc_f_xuser_15_xuser(int_rd_resp_desc_f_xuser_15_xuser),
                   .int_wr_req_desc_f_data_host_addr_0_addr(int_wr_req_desc_f_data_host_addr_0_addr),
                   .int_wr_req_desc_f_data_host_addr_1_addr(int_wr_req_desc_f_data_host_addr_1_addr),
                   .int_wr_req_desc_f_data_host_addr_2_addr(int_wr_req_desc_f_data_host_addr_2_addr),
                   .int_wr_req_desc_f_data_host_addr_3_addr(int_wr_req_desc_f_data_host_addr_3_addr),
                   .int_wr_req_desc_f_wstrb_host_addr_0_addr(int_wr_req_desc_f_wstrb_host_addr_0_addr),
                   .int_wr_req_desc_f_wstrb_host_addr_1_addr(int_wr_req_desc_f_wstrb_host_addr_1_addr),
                   .int_wr_req_desc_f_wstrb_host_addr_2_addr(int_wr_req_desc_f_wstrb_host_addr_2_addr),
                   .int_wr_req_desc_f_wstrb_host_addr_3_addr(int_wr_req_desc_f_wstrb_host_addr_3_addr),
                   .int_wr_resp_desc_f_resp_resp(int_wr_resp_desc_f_resp_resp),
                   .int_wr_resp_desc_f_xid_0_xid(int_wr_resp_desc_f_xid_0_xid),
                   .int_wr_resp_desc_f_xid_1_xid(int_wr_resp_desc_f_xid_1_xid),
                   .int_wr_resp_desc_f_xid_2_xid(int_wr_resp_desc_f_xid_2_xid),
                   .int_wr_resp_desc_f_xid_3_xid(int_wr_resp_desc_f_xid_3_xid),
                   .int_wr_resp_desc_f_xuser_0_xuser(int_wr_resp_desc_f_xuser_0_xuser),
                   .int_wr_resp_desc_f_xuser_1_xuser(int_wr_resp_desc_f_xuser_1_xuser),
                   .int_wr_resp_desc_f_xuser_2_xuser(int_wr_resp_desc_f_xuser_2_xuser),
                   .int_wr_resp_desc_f_xuser_3_xuser(int_wr_resp_desc_f_xuser_3_xuser),
                   .int_wr_resp_desc_f_xuser_4_xuser(int_wr_resp_desc_f_xuser_4_xuser),
                   .int_wr_resp_desc_f_xuser_5_xuser(int_wr_resp_desc_f_xuser_5_xuser),
                   .int_wr_resp_desc_f_xuser_6_xuser(int_wr_resp_desc_f_xuser_6_xuser),
                   .int_wr_resp_desc_f_xuser_7_xuser(int_wr_resp_desc_f_xuser_7_xuser),
                   .int_wr_resp_desc_f_xuser_8_xuser(int_wr_resp_desc_f_xuser_8_xuser),
                   .int_wr_resp_desc_f_xuser_9_xuser(int_wr_resp_desc_f_xuser_9_xuser),
                   .int_wr_resp_desc_f_xuser_10_xuser(int_wr_resp_desc_f_xuser_10_xuser),
                   .int_wr_resp_desc_f_xuser_11_xuser(int_wr_resp_desc_f_xuser_11_xuser),
                   .int_wr_resp_desc_f_xuser_12_xuser(int_wr_resp_desc_f_xuser_12_xuser),
                   .int_wr_resp_desc_f_xuser_13_xuser(int_wr_resp_desc_f_xuser_13_xuser),
                   .int_wr_resp_desc_f_xuser_14_xuser(int_wr_resp_desc_f_xuser_14_xuser),
                   .int_wr_resp_desc_f_xuser_15_xuser(int_wr_resp_desc_f_xuser_15_xuser),
                   .int_sn_req_desc_f_attr_acsnoop(int_sn_req_desc_f_attr_acsnoop),
                   .int_sn_req_desc_f_attr_acprot(int_sn_req_desc_f_attr_acprot),
                   .int_sn_req_desc_f_acaddr_0_addr(int_sn_req_desc_f_acaddr_0_addr),
                   .int_sn_req_desc_f_acaddr_1_addr(int_sn_req_desc_f_acaddr_1_addr),
                   .int_sn_req_desc_f_acaddr_2_addr(int_sn_req_desc_f_acaddr_2_addr),
                   .int_sn_req_desc_f_acaddr_3_addr(int_sn_req_desc_f_acaddr_3_addr),
                   .rd_req_fifo_out(rd_req_fifo_out),
                   .rd_req_fifo_out_valid(rd_req_fifo_out_valid),
                   .wr_req_fifo_out(wr_req_fifo_out),
                   .wr_req_fifo_out_valid(wr_req_fifo_out_valid),
                   .sn_resp_fifo_out(sn_resp_fifo_out),
                   .sn_resp_fifo_out_valid(sn_resp_fifo_out_valid),
                   .sn_data_fifo_out(sn_data_fifo_out),
                   .sn_data_fifo_out_valid(sn_data_fifo_out_valid)
      
      
      
      
                   );


   //        `include "int_desc_port_inst.vh"
   
   

endmodule

