/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *   This Module Implements Register Module for Slave Bridge for 128KB memory requirement.
 *
 *
 */


`include "ace_defines_common.vh"
`include "ace_defines_slv_regspace.vh"
module ace_regs_slv #(

                       parameter ACE_PROTOCOL                   = "FULLACE" 
                       
                       ,parameter S_AXI_ADDR_WIDTH               = 64 
                       ,parameter S_AXI_DATA_WIDTH               = 32 
                       
                       ,parameter S_ACE_USR_ADDR_WIDTH           = 64 
                       ,parameter S_ACE_USR_XX_DATA_WIDTH        = 128       
                       ,parameter S_ACE_USR_SN_DATA_WIDTH        = 128       
                       ,parameter S_ACE_USR_ID_WIDTH             = 16 
                       ,parameter S_ACE_USR_AWUSER_WIDTH         = 32 
                       ,parameter S_ACE_USR_WUSER_WIDTH          = 32 
                       ,parameter S_ACE_USR_BUSER_WIDTH          = 32 
                       ,parameter S_ACE_USR_ARUSER_WIDTH         = 32 
                       ,parameter S_ACE_USR_RUSER_WIDTH          = 32 
                       
                       ,parameter CACHE_LINE_SIZE                = 64 
                       ,parameter XX_MAX_DESC                    = 16         
                       ,parameter SN_MAX_DESC                    = 16         
                       ,parameter XX_RAM_SIZE                    = 16384     
                       ,parameter SN_RAM_SIZE                    = 1024       
                       ,parameter USR_RST_NUM                    = 4     

                       ,parameter LAST_BRIDGE                    = 0
                       ,parameter EXTEND_WSTRB                   = 1 
                       
                       


                       )
   (
    input clk
    ,input resetn // Top level AXI reset. Typically derived from Reset issued by Pcie Host. Drives AXI FSM and 'reset_reg' of this module.
    ,input rst_n // combination of 'resetn' and Bridge SRST. Drives all Regs and RAMs in this module. 
    
    // S_AXI - AXI4-Lite
    ,input wire [S_AXI_ADDR_WIDTH-1:0] s_axi_awaddr
    ,input wire [2:0] s_axi_awprot
    ,input wire s_axi_awvalid
    ,output wire s_axi_awready
    ,input wire [S_AXI_DATA_WIDTH-1:0] s_axi_wdata
    ,input wire [(S_AXI_DATA_WIDTH/8)-1:0] s_axi_wstrb
    ,input wire s_axi_wvalid
    ,output wire s_axi_wready
    ,output wire [1:0] s_axi_bresp
    ,output wire s_axi_bvalid
    ,input wire s_axi_bready
    ,input wire [S_AXI_ADDR_WIDTH-1:0] s_axi_araddr
    ,input wire [2:0] s_axi_arprot
    ,input wire s_axi_arvalid
    ,output wire s_axi_arready
    ,output wire [S_AXI_DATA_WIDTH-1:0] s_axi_rdata
    ,output wire [1:0] s_axi_rresp
    ,output wire s_axi_rvalid
    ,input wire s_axi_rready
    
    //RDATA_RAM
    ,input [(`CLOG2((XX_RAM_SIZE*8)/S_ACE_USR_XX_DATA_WIDTH))-1:0] uc2rb_rd_addr 
    ,output [S_ACE_USR_XX_DATA_WIDTH-1:0] rb2uc_rd_data 
    
    //WDATA_RAM and WSTRB_RAM                               
    ,input uc2rb_wr_we 
    ,input [(S_ACE_USR_XX_DATA_WIDTH/8)-1:0] uc2rb_wr_bwe 
    ,input [(`CLOG2((XX_RAM_SIZE*8)/S_ACE_USR_XX_DATA_WIDTH))-1:0] uc2rb_wr_addr 
    ,input [S_ACE_USR_XX_DATA_WIDTH-1:0] uc2rb_wr_data 
    ,input [(S_ACE_USR_XX_DATA_WIDTH/8)-1:0] uc2rb_wr_wstrb 
    
    //CDDATA_RAM                               
    ,input uc2rb_sn_we 
    ,input [(S_ACE_USR_SN_DATA_WIDTH/8)-1:0] uc2rb_sn_bwe 
    ,input [(`CLOG2((SN_RAM_SIZE*8)/S_ACE_USR_SN_DATA_WIDTH))-1:0] uc2rb_sn_addr 
    ,input [S_ACE_USR_SN_DATA_WIDTH-1:0] uc2rb_sn_data 
    
    // Mode 1 Signals
    // Read port of WR DataRam
    ,input [(`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8)))-1:0] hm2rb_rd_addr 
    ,output reg [S_ACE_USR_XX_DATA_WIDTH-1:0] rb2hm_rd_data 
    ,output reg [(S_ACE_USR_XX_DATA_WIDTH/8 -1):0] rb2hm_rd_wstrb
    // Write port of RD DataRam
    ,input hm2rb_wr_we 
    ,input [(S_ACE_USR_XX_DATA_WIDTH/8 -1):0] hm2rb_wr_bwe 
    ,input [(`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8)))-1:0] hm2rb_wr_addr 
    ,input [S_ACE_USR_XX_DATA_WIDTH-1:0] hm2rb_wr_data
    
    //pop request to FIFO
    ,output reg rd_req_fifo_pop_desc_conn 
    ,output reg wr_req_fifo_pop_desc_conn 
    ,output reg sn_resp_fifo_pop_desc_conn
    ,output reg sn_data_fifo_pop_desc_conn
    
    //output from FIFO
    ,input [(`CLOG2(XX_MAX_DESC))-1:0] rd_req_fifo_out
    ,input rd_req_fifo_out_valid //it is one clock cycle pulse
    ,input [(`CLOG2(XX_MAX_DESC))-1:0] wr_req_fifo_out
    ,input wr_req_fifo_out_valid //it is one clock cycle pulse
    ,input [(`CLOG2(SN_MAX_DESC))-1:0] sn_resp_fifo_out
    ,input sn_resp_fifo_out_valid //it is one clock cycle pulse
    ,input [(`CLOG2(SN_MAX_DESC))-1:0] sn_data_fifo_out
    ,input sn_data_fifo_out_valid //it is one clock cycle pulse
    
    
    
    // Registers
    ,output reg [31:0] bridge_identification_reg
    ,output reg [31:0] last_bridge_reg
    ,output reg [31:0] version_reg
    ,output reg [31:0] bridge_type_reg
    ,output reg [31:0] mode_select_reg
    ,output reg [31:0] reset_reg
    ,output reg [31:0] h2c_intr_0_reg
    ,output reg [31:0] h2c_intr_1_reg
    ,output reg [31:0] h2c_intr_2_reg
    ,output reg [31:0] h2c_intr_3_reg
    ,output reg [31:0] c2h_intr_status_0_reg
    ,output reg [31:0] intr_c2h_toggle_status_0_reg
    ,output reg [31:0] intr_c2h_toggle_clear_0_reg
    ,output reg [31:0] intr_c2h_toggle_enable_0_reg
    ,output reg [31:0] c2h_intr_status_1_reg
    ,output reg [31:0] intr_c2h_toggle_status_1_reg
    ,output reg [31:0] intr_c2h_toggle_clear_1_reg
    ,output reg [31:0] intr_c2h_toggle_enable_1_reg
    ,output reg [31:0] c2h_gpio_0_reg
    ,output reg [31:0] c2h_gpio_1_reg
    ,output reg [31:0] c2h_gpio_2_reg
    ,output reg [31:0] c2h_gpio_3_reg
    ,output reg [31:0] c2h_gpio_4_reg
    ,output reg [31:0] c2h_gpio_5_reg
    ,output reg [31:0] c2h_gpio_6_reg
    ,output reg [31:0] c2h_gpio_7_reg
    ,output reg [31:0] c2h_gpio_8_reg
    ,output reg [31:0] c2h_gpio_9_reg
    ,output reg [31:0] c2h_gpio_10_reg
    ,output reg [31:0] c2h_gpio_11_reg
    ,output reg [31:0] c2h_gpio_12_reg
    ,output reg [31:0] c2h_gpio_13_reg
    ,output reg [31:0] c2h_gpio_14_reg
    ,output reg [31:0] c2h_gpio_15_reg
    ,output reg [31:0] h2c_gpio_0_reg
    ,output reg [31:0] h2c_gpio_1_reg
    ,output reg [31:0] h2c_gpio_2_reg
    ,output reg [31:0] h2c_gpio_3_reg
    ,output reg [31:0] h2c_gpio_4_reg
    ,output reg [31:0] h2c_gpio_5_reg
    ,output reg [31:0] h2c_gpio_6_reg
    ,output reg [31:0] h2c_gpio_7_reg
    ,output reg [31:0] h2c_gpio_8_reg
    ,output reg [31:0] h2c_gpio_9_reg
    ,output reg [31:0] h2c_gpio_10_reg
    ,output reg [31:0] h2c_gpio_11_reg
    ,output reg [31:0] h2c_gpio_12_reg
    ,output reg [31:0] h2c_gpio_13_reg
    ,output reg [31:0] h2c_gpio_14_reg
    ,output reg [31:0] h2c_gpio_15_reg
    ,output reg [31:0] bridge_config_reg
    ,output reg [31:0] intr_status_reg
    ,output reg [31:0] intr_error_status_reg
    ,output reg [31:0] intr_error_clear_reg
    ,output reg [31:0] intr_error_enable_reg
    ,output reg [31:0] bridge_rd_user_config_reg
    ,output reg [31:0] bridge_wr_user_config_reg
    ,output reg [31:0] rd_max_desc_reg
    ,output reg [31:0] wr_max_desc_reg
    ,output reg [31:0] sn_max_desc_reg
    ,output reg [31:0] rd_req_free_desc_reg
    ,output reg [31:0] rd_req_fifo_pop_desc_reg
    ,output reg [31:0] rd_req_fifo_fill_level_reg
    ,output reg [31:0] rd_resp_fifo_push_desc_reg
    ,output reg [31:0] rd_resp_fifo_free_level_reg
    ,output reg [31:0] rd_resp_intr_comp_status_reg
    ,output reg [31:0] rd_resp_intr_comp_clear_reg
    ,output reg [31:0] rd_resp_intr_comp_enable_reg
    ,output reg [31:0] wr_req_free_desc_reg
    ,output reg [31:0] wr_req_fifo_pop_desc_reg
    ,output reg [31:0] wr_req_fifo_fill_level_reg
    ,output reg [31:0] wr_resp_fifo_push_desc_reg
    ,output reg [31:0] wr_resp_fifo_free_level_reg
    ,output reg [31:0] wr_resp_intr_comp_status_reg
    ,output reg [31:0] wr_resp_intr_comp_clear_reg
    ,output reg [31:0] wr_resp_intr_comp_enable_reg
    ,output reg [31:0] sn_req_fifo_push_desc_reg
    ,output reg [31:0] sn_req_fifo_free_level_reg
    ,output reg [31:0] sn_req_intr_comp_status_reg
    ,output reg [31:0] sn_req_intr_comp_clear_reg
    ,output reg [31:0] sn_req_intr_comp_enable_reg
    ,output reg [31:0] sn_resp_free_desc_reg
    ,output reg [31:0] sn_resp_fifo_pop_desc_reg
    ,output reg [31:0] sn_resp_fifo_fill_level_reg
    ,output reg [31:0] sn_data_free_desc_reg
    ,output reg [31:0] sn_data_fifo_pop_desc_reg
    ,output reg [31:0] sn_data_fifo_fill_level_reg
    ,output reg [31:0] intr_fifo_enable_reg
    ,output reg [31:0] rd_req_desc_0_txn_type_reg
    ,output reg [31:0] rd_req_desc_0_size_reg
    ,output reg [31:0] rd_req_desc_0_axsize_reg
    ,output reg [31:0] rd_req_desc_0_attr_reg
    ,output reg [31:0] rd_req_desc_0_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_0_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_0_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_0_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_0_axid_0_reg
    ,output reg [31:0] rd_req_desc_0_axid_1_reg
    ,output reg [31:0] rd_req_desc_0_axid_2_reg
    ,output reg [31:0] rd_req_desc_0_axid_3_reg
    ,output reg [31:0] rd_req_desc_0_axuser_0_reg
    ,output reg [31:0] rd_req_desc_0_axuser_1_reg
    ,output reg [31:0] rd_req_desc_0_axuser_2_reg
    ,output reg [31:0] rd_req_desc_0_axuser_3_reg
    ,output reg [31:0] rd_req_desc_0_axuser_4_reg
    ,output reg [31:0] rd_req_desc_0_axuser_5_reg
    ,output reg [31:0] rd_req_desc_0_axuser_6_reg
    ,output reg [31:0] rd_req_desc_0_axuser_7_reg
    ,output reg [31:0] rd_req_desc_0_axuser_8_reg
    ,output reg [31:0] rd_req_desc_0_axuser_9_reg
    ,output reg [31:0] rd_req_desc_0_axuser_10_reg
    ,output reg [31:0] rd_req_desc_0_axuser_11_reg
    ,output reg [31:0] rd_req_desc_0_axuser_12_reg
    ,output reg [31:0] rd_req_desc_0_axuser_13_reg
    ,output reg [31:0] rd_req_desc_0_axuser_14_reg
    ,output reg [31:0] rd_req_desc_0_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_0_data_offset_reg
    ,output reg [31:0] rd_resp_desc_0_data_size_reg
    ,output reg [31:0] rd_resp_desc_0_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_0_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_0_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_0_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_0_resp_reg
    ,output reg [31:0] rd_resp_desc_0_xid_0_reg
    ,output reg [31:0] rd_resp_desc_0_xid_1_reg
    ,output reg [31:0] rd_resp_desc_0_xid_2_reg
    ,output reg [31:0] rd_resp_desc_0_xid_3_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_0_xuser_15_reg
    ,output reg [31:0] wr_req_desc_0_txn_type_reg
    ,output reg [31:0] wr_req_desc_0_size_reg
    ,output reg [31:0] wr_req_desc_0_data_offset_reg
    ,output reg [31:0] wr_req_desc_0_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_0_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_0_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_0_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_0_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_0_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_0_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_0_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_0_axsize_reg
    ,output reg [31:0] wr_req_desc_0_attr_reg
    ,output reg [31:0] wr_req_desc_0_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_0_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_0_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_0_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_0_axid_0_reg
    ,output reg [31:0] wr_req_desc_0_axid_1_reg
    ,output reg [31:0] wr_req_desc_0_axid_2_reg
    ,output reg [31:0] wr_req_desc_0_axid_3_reg
    ,output reg [31:0] wr_req_desc_0_axuser_0_reg
    ,output reg [31:0] wr_req_desc_0_axuser_1_reg
    ,output reg [31:0] wr_req_desc_0_axuser_2_reg
    ,output reg [31:0] wr_req_desc_0_axuser_3_reg
    ,output reg [31:0] wr_req_desc_0_axuser_4_reg
    ,output reg [31:0] wr_req_desc_0_axuser_5_reg
    ,output reg [31:0] wr_req_desc_0_axuser_6_reg
    ,output reg [31:0] wr_req_desc_0_axuser_7_reg
    ,output reg [31:0] wr_req_desc_0_axuser_8_reg
    ,output reg [31:0] wr_req_desc_0_axuser_9_reg
    ,output reg [31:0] wr_req_desc_0_axuser_10_reg
    ,output reg [31:0] wr_req_desc_0_axuser_11_reg
    ,output reg [31:0] wr_req_desc_0_axuser_12_reg
    ,output reg [31:0] wr_req_desc_0_axuser_13_reg
    ,output reg [31:0] wr_req_desc_0_axuser_14_reg
    ,output reg [31:0] wr_req_desc_0_axuser_15_reg
    ,output reg [31:0] wr_req_desc_0_wuser_0_reg
    ,output reg [31:0] wr_req_desc_0_wuser_1_reg
    ,output reg [31:0] wr_req_desc_0_wuser_2_reg
    ,output reg [31:0] wr_req_desc_0_wuser_3_reg
    ,output reg [31:0] wr_req_desc_0_wuser_4_reg
    ,output reg [31:0] wr_req_desc_0_wuser_5_reg
    ,output reg [31:0] wr_req_desc_0_wuser_6_reg
    ,output reg [31:0] wr_req_desc_0_wuser_7_reg
    ,output reg [31:0] wr_req_desc_0_wuser_8_reg
    ,output reg [31:0] wr_req_desc_0_wuser_9_reg
    ,output reg [31:0] wr_req_desc_0_wuser_10_reg
    ,output reg [31:0] wr_req_desc_0_wuser_11_reg
    ,output reg [31:0] wr_req_desc_0_wuser_12_reg
    ,output reg [31:0] wr_req_desc_0_wuser_13_reg
    ,output reg [31:0] wr_req_desc_0_wuser_14_reg
    ,output reg [31:0] wr_req_desc_0_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_0_resp_reg
    ,output reg [31:0] wr_resp_desc_0_xid_0_reg
    ,output reg [31:0] wr_resp_desc_0_xid_1_reg
    ,output reg [31:0] wr_resp_desc_0_xid_2_reg
    ,output reg [31:0] wr_resp_desc_0_xid_3_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_0_xuser_15_reg
    ,output reg [31:0] sn_req_desc_0_attr_reg
    ,output reg [31:0] sn_req_desc_0_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_0_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_0_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_0_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_0_resp_reg
    ,output reg [31:0] rd_req_desc_1_txn_type_reg
    ,output reg [31:0] rd_req_desc_1_size_reg
    ,output reg [31:0] rd_req_desc_1_axsize_reg
    ,output reg [31:0] rd_req_desc_1_attr_reg
    ,output reg [31:0] rd_req_desc_1_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_1_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_1_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_1_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_1_axid_0_reg
    ,output reg [31:0] rd_req_desc_1_axid_1_reg
    ,output reg [31:0] rd_req_desc_1_axid_2_reg
    ,output reg [31:0] rd_req_desc_1_axid_3_reg
    ,output reg [31:0] rd_req_desc_1_axuser_0_reg
    ,output reg [31:0] rd_req_desc_1_axuser_1_reg
    ,output reg [31:0] rd_req_desc_1_axuser_2_reg
    ,output reg [31:0] rd_req_desc_1_axuser_3_reg
    ,output reg [31:0] rd_req_desc_1_axuser_4_reg
    ,output reg [31:0] rd_req_desc_1_axuser_5_reg
    ,output reg [31:0] rd_req_desc_1_axuser_6_reg
    ,output reg [31:0] rd_req_desc_1_axuser_7_reg
    ,output reg [31:0] rd_req_desc_1_axuser_8_reg
    ,output reg [31:0] rd_req_desc_1_axuser_9_reg
    ,output reg [31:0] rd_req_desc_1_axuser_10_reg
    ,output reg [31:0] rd_req_desc_1_axuser_11_reg
    ,output reg [31:0] rd_req_desc_1_axuser_12_reg
    ,output reg [31:0] rd_req_desc_1_axuser_13_reg
    ,output reg [31:0] rd_req_desc_1_axuser_14_reg
    ,output reg [31:0] rd_req_desc_1_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_1_data_offset_reg
    ,output reg [31:0] rd_resp_desc_1_data_size_reg
    ,output reg [31:0] rd_resp_desc_1_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_1_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_1_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_1_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_1_resp_reg
    ,output reg [31:0] rd_resp_desc_1_xid_0_reg
    ,output reg [31:0] rd_resp_desc_1_xid_1_reg
    ,output reg [31:0] rd_resp_desc_1_xid_2_reg
    ,output reg [31:0] rd_resp_desc_1_xid_3_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_1_xuser_15_reg
    ,output reg [31:0] wr_req_desc_1_txn_type_reg
    ,output reg [31:0] wr_req_desc_1_size_reg
    ,output reg [31:0] wr_req_desc_1_data_offset_reg
    ,output reg [31:0] wr_req_desc_1_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_1_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_1_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_1_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_1_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_1_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_1_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_1_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_1_axsize_reg
    ,output reg [31:0] wr_req_desc_1_attr_reg
    ,output reg [31:0] wr_req_desc_1_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_1_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_1_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_1_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_1_axid_0_reg
    ,output reg [31:0] wr_req_desc_1_axid_1_reg
    ,output reg [31:0] wr_req_desc_1_axid_2_reg
    ,output reg [31:0] wr_req_desc_1_axid_3_reg
    ,output reg [31:0] wr_req_desc_1_axuser_0_reg
    ,output reg [31:0] wr_req_desc_1_axuser_1_reg
    ,output reg [31:0] wr_req_desc_1_axuser_2_reg
    ,output reg [31:0] wr_req_desc_1_axuser_3_reg
    ,output reg [31:0] wr_req_desc_1_axuser_4_reg
    ,output reg [31:0] wr_req_desc_1_axuser_5_reg
    ,output reg [31:0] wr_req_desc_1_axuser_6_reg
    ,output reg [31:0] wr_req_desc_1_axuser_7_reg
    ,output reg [31:0] wr_req_desc_1_axuser_8_reg
    ,output reg [31:0] wr_req_desc_1_axuser_9_reg
    ,output reg [31:0] wr_req_desc_1_axuser_10_reg
    ,output reg [31:0] wr_req_desc_1_axuser_11_reg
    ,output reg [31:0] wr_req_desc_1_axuser_12_reg
    ,output reg [31:0] wr_req_desc_1_axuser_13_reg
    ,output reg [31:0] wr_req_desc_1_axuser_14_reg
    ,output reg [31:0] wr_req_desc_1_axuser_15_reg
    ,output reg [31:0] wr_req_desc_1_wuser_0_reg
    ,output reg [31:0] wr_req_desc_1_wuser_1_reg
    ,output reg [31:0] wr_req_desc_1_wuser_2_reg
    ,output reg [31:0] wr_req_desc_1_wuser_3_reg
    ,output reg [31:0] wr_req_desc_1_wuser_4_reg
    ,output reg [31:0] wr_req_desc_1_wuser_5_reg
    ,output reg [31:0] wr_req_desc_1_wuser_6_reg
    ,output reg [31:0] wr_req_desc_1_wuser_7_reg
    ,output reg [31:0] wr_req_desc_1_wuser_8_reg
    ,output reg [31:0] wr_req_desc_1_wuser_9_reg
    ,output reg [31:0] wr_req_desc_1_wuser_10_reg
    ,output reg [31:0] wr_req_desc_1_wuser_11_reg
    ,output reg [31:0] wr_req_desc_1_wuser_12_reg
    ,output reg [31:0] wr_req_desc_1_wuser_13_reg
    ,output reg [31:0] wr_req_desc_1_wuser_14_reg
    ,output reg [31:0] wr_req_desc_1_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_1_resp_reg
    ,output reg [31:0] wr_resp_desc_1_xid_0_reg
    ,output reg [31:0] wr_resp_desc_1_xid_1_reg
    ,output reg [31:0] wr_resp_desc_1_xid_2_reg
    ,output reg [31:0] wr_resp_desc_1_xid_3_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_1_xuser_15_reg
    ,output reg [31:0] sn_req_desc_1_attr_reg
    ,output reg [31:0] sn_req_desc_1_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_1_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_1_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_1_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_1_resp_reg
    ,output reg [31:0] rd_req_desc_2_txn_type_reg
    ,output reg [31:0] rd_req_desc_2_size_reg
    ,output reg [31:0] rd_req_desc_2_axsize_reg
    ,output reg [31:0] rd_req_desc_2_attr_reg
    ,output reg [31:0] rd_req_desc_2_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_2_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_2_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_2_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_2_axid_0_reg
    ,output reg [31:0] rd_req_desc_2_axid_1_reg
    ,output reg [31:0] rd_req_desc_2_axid_2_reg
    ,output reg [31:0] rd_req_desc_2_axid_3_reg
    ,output reg [31:0] rd_req_desc_2_axuser_0_reg
    ,output reg [31:0] rd_req_desc_2_axuser_1_reg
    ,output reg [31:0] rd_req_desc_2_axuser_2_reg
    ,output reg [31:0] rd_req_desc_2_axuser_3_reg
    ,output reg [31:0] rd_req_desc_2_axuser_4_reg
    ,output reg [31:0] rd_req_desc_2_axuser_5_reg
    ,output reg [31:0] rd_req_desc_2_axuser_6_reg
    ,output reg [31:0] rd_req_desc_2_axuser_7_reg
    ,output reg [31:0] rd_req_desc_2_axuser_8_reg
    ,output reg [31:0] rd_req_desc_2_axuser_9_reg
    ,output reg [31:0] rd_req_desc_2_axuser_10_reg
    ,output reg [31:0] rd_req_desc_2_axuser_11_reg
    ,output reg [31:0] rd_req_desc_2_axuser_12_reg
    ,output reg [31:0] rd_req_desc_2_axuser_13_reg
    ,output reg [31:0] rd_req_desc_2_axuser_14_reg
    ,output reg [31:0] rd_req_desc_2_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_2_data_offset_reg
    ,output reg [31:0] rd_resp_desc_2_data_size_reg
    ,output reg [31:0] rd_resp_desc_2_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_2_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_2_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_2_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_2_resp_reg
    ,output reg [31:0] rd_resp_desc_2_xid_0_reg
    ,output reg [31:0] rd_resp_desc_2_xid_1_reg
    ,output reg [31:0] rd_resp_desc_2_xid_2_reg
    ,output reg [31:0] rd_resp_desc_2_xid_3_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_2_xuser_15_reg
    ,output reg [31:0] wr_req_desc_2_txn_type_reg
    ,output reg [31:0] wr_req_desc_2_size_reg
    ,output reg [31:0] wr_req_desc_2_data_offset_reg
    ,output reg [31:0] wr_req_desc_2_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_2_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_2_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_2_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_2_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_2_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_2_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_2_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_2_axsize_reg
    ,output reg [31:0] wr_req_desc_2_attr_reg
    ,output reg [31:0] wr_req_desc_2_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_2_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_2_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_2_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_2_axid_0_reg
    ,output reg [31:0] wr_req_desc_2_axid_1_reg
    ,output reg [31:0] wr_req_desc_2_axid_2_reg
    ,output reg [31:0] wr_req_desc_2_axid_3_reg
    ,output reg [31:0] wr_req_desc_2_axuser_0_reg
    ,output reg [31:0] wr_req_desc_2_axuser_1_reg
    ,output reg [31:0] wr_req_desc_2_axuser_2_reg
    ,output reg [31:0] wr_req_desc_2_axuser_3_reg
    ,output reg [31:0] wr_req_desc_2_axuser_4_reg
    ,output reg [31:0] wr_req_desc_2_axuser_5_reg
    ,output reg [31:0] wr_req_desc_2_axuser_6_reg
    ,output reg [31:0] wr_req_desc_2_axuser_7_reg
    ,output reg [31:0] wr_req_desc_2_axuser_8_reg
    ,output reg [31:0] wr_req_desc_2_axuser_9_reg
    ,output reg [31:0] wr_req_desc_2_axuser_10_reg
    ,output reg [31:0] wr_req_desc_2_axuser_11_reg
    ,output reg [31:0] wr_req_desc_2_axuser_12_reg
    ,output reg [31:0] wr_req_desc_2_axuser_13_reg
    ,output reg [31:0] wr_req_desc_2_axuser_14_reg
    ,output reg [31:0] wr_req_desc_2_axuser_15_reg
    ,output reg [31:0] wr_req_desc_2_wuser_0_reg
    ,output reg [31:0] wr_req_desc_2_wuser_1_reg
    ,output reg [31:0] wr_req_desc_2_wuser_2_reg
    ,output reg [31:0] wr_req_desc_2_wuser_3_reg
    ,output reg [31:0] wr_req_desc_2_wuser_4_reg
    ,output reg [31:0] wr_req_desc_2_wuser_5_reg
    ,output reg [31:0] wr_req_desc_2_wuser_6_reg
    ,output reg [31:0] wr_req_desc_2_wuser_7_reg
    ,output reg [31:0] wr_req_desc_2_wuser_8_reg
    ,output reg [31:0] wr_req_desc_2_wuser_9_reg
    ,output reg [31:0] wr_req_desc_2_wuser_10_reg
    ,output reg [31:0] wr_req_desc_2_wuser_11_reg
    ,output reg [31:0] wr_req_desc_2_wuser_12_reg
    ,output reg [31:0] wr_req_desc_2_wuser_13_reg
    ,output reg [31:0] wr_req_desc_2_wuser_14_reg
    ,output reg [31:0] wr_req_desc_2_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_2_resp_reg
    ,output reg [31:0] wr_resp_desc_2_xid_0_reg
    ,output reg [31:0] wr_resp_desc_2_xid_1_reg
    ,output reg [31:0] wr_resp_desc_2_xid_2_reg
    ,output reg [31:0] wr_resp_desc_2_xid_3_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_2_xuser_15_reg
    ,output reg [31:0] sn_req_desc_2_attr_reg
    ,output reg [31:0] sn_req_desc_2_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_2_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_2_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_2_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_2_resp_reg
    ,output reg [31:0] rd_req_desc_3_txn_type_reg
    ,output reg [31:0] rd_req_desc_3_size_reg
    ,output reg [31:0] rd_req_desc_3_axsize_reg
    ,output reg [31:0] rd_req_desc_3_attr_reg
    ,output reg [31:0] rd_req_desc_3_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_3_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_3_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_3_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_3_axid_0_reg
    ,output reg [31:0] rd_req_desc_3_axid_1_reg
    ,output reg [31:0] rd_req_desc_3_axid_2_reg
    ,output reg [31:0] rd_req_desc_3_axid_3_reg
    ,output reg [31:0] rd_req_desc_3_axuser_0_reg
    ,output reg [31:0] rd_req_desc_3_axuser_1_reg
    ,output reg [31:0] rd_req_desc_3_axuser_2_reg
    ,output reg [31:0] rd_req_desc_3_axuser_3_reg
    ,output reg [31:0] rd_req_desc_3_axuser_4_reg
    ,output reg [31:0] rd_req_desc_3_axuser_5_reg
    ,output reg [31:0] rd_req_desc_3_axuser_6_reg
    ,output reg [31:0] rd_req_desc_3_axuser_7_reg
    ,output reg [31:0] rd_req_desc_3_axuser_8_reg
    ,output reg [31:0] rd_req_desc_3_axuser_9_reg
    ,output reg [31:0] rd_req_desc_3_axuser_10_reg
    ,output reg [31:0] rd_req_desc_3_axuser_11_reg
    ,output reg [31:0] rd_req_desc_3_axuser_12_reg
    ,output reg [31:0] rd_req_desc_3_axuser_13_reg
    ,output reg [31:0] rd_req_desc_3_axuser_14_reg
    ,output reg [31:0] rd_req_desc_3_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_3_data_offset_reg
    ,output reg [31:0] rd_resp_desc_3_data_size_reg
    ,output reg [31:0] rd_resp_desc_3_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_3_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_3_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_3_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_3_resp_reg
    ,output reg [31:0] rd_resp_desc_3_xid_0_reg
    ,output reg [31:0] rd_resp_desc_3_xid_1_reg
    ,output reg [31:0] rd_resp_desc_3_xid_2_reg
    ,output reg [31:0] rd_resp_desc_3_xid_3_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_3_xuser_15_reg
    ,output reg [31:0] wr_req_desc_3_txn_type_reg
    ,output reg [31:0] wr_req_desc_3_size_reg
    ,output reg [31:0] wr_req_desc_3_data_offset_reg
    ,output reg [31:0] wr_req_desc_3_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_3_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_3_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_3_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_3_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_3_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_3_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_3_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_3_axsize_reg
    ,output reg [31:0] wr_req_desc_3_attr_reg
    ,output reg [31:0] wr_req_desc_3_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_3_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_3_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_3_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_3_axid_0_reg
    ,output reg [31:0] wr_req_desc_3_axid_1_reg
    ,output reg [31:0] wr_req_desc_3_axid_2_reg
    ,output reg [31:0] wr_req_desc_3_axid_3_reg
    ,output reg [31:0] wr_req_desc_3_axuser_0_reg
    ,output reg [31:0] wr_req_desc_3_axuser_1_reg
    ,output reg [31:0] wr_req_desc_3_axuser_2_reg
    ,output reg [31:0] wr_req_desc_3_axuser_3_reg
    ,output reg [31:0] wr_req_desc_3_axuser_4_reg
    ,output reg [31:0] wr_req_desc_3_axuser_5_reg
    ,output reg [31:0] wr_req_desc_3_axuser_6_reg
    ,output reg [31:0] wr_req_desc_3_axuser_7_reg
    ,output reg [31:0] wr_req_desc_3_axuser_8_reg
    ,output reg [31:0] wr_req_desc_3_axuser_9_reg
    ,output reg [31:0] wr_req_desc_3_axuser_10_reg
    ,output reg [31:0] wr_req_desc_3_axuser_11_reg
    ,output reg [31:0] wr_req_desc_3_axuser_12_reg
    ,output reg [31:0] wr_req_desc_3_axuser_13_reg
    ,output reg [31:0] wr_req_desc_3_axuser_14_reg
    ,output reg [31:0] wr_req_desc_3_axuser_15_reg
    ,output reg [31:0] wr_req_desc_3_wuser_0_reg
    ,output reg [31:0] wr_req_desc_3_wuser_1_reg
    ,output reg [31:0] wr_req_desc_3_wuser_2_reg
    ,output reg [31:0] wr_req_desc_3_wuser_3_reg
    ,output reg [31:0] wr_req_desc_3_wuser_4_reg
    ,output reg [31:0] wr_req_desc_3_wuser_5_reg
    ,output reg [31:0] wr_req_desc_3_wuser_6_reg
    ,output reg [31:0] wr_req_desc_3_wuser_7_reg
    ,output reg [31:0] wr_req_desc_3_wuser_8_reg
    ,output reg [31:0] wr_req_desc_3_wuser_9_reg
    ,output reg [31:0] wr_req_desc_3_wuser_10_reg
    ,output reg [31:0] wr_req_desc_3_wuser_11_reg
    ,output reg [31:0] wr_req_desc_3_wuser_12_reg
    ,output reg [31:0] wr_req_desc_3_wuser_13_reg
    ,output reg [31:0] wr_req_desc_3_wuser_14_reg
    ,output reg [31:0] wr_req_desc_3_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_3_resp_reg
    ,output reg [31:0] wr_resp_desc_3_xid_0_reg
    ,output reg [31:0] wr_resp_desc_3_xid_1_reg
    ,output reg [31:0] wr_resp_desc_3_xid_2_reg
    ,output reg [31:0] wr_resp_desc_3_xid_3_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_3_xuser_15_reg
    ,output reg [31:0] sn_req_desc_3_attr_reg
    ,output reg [31:0] sn_req_desc_3_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_3_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_3_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_3_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_3_resp_reg
    ,output reg [31:0] rd_req_desc_4_txn_type_reg
    ,output reg [31:0] rd_req_desc_4_size_reg
    ,output reg [31:0] rd_req_desc_4_axsize_reg
    ,output reg [31:0] rd_req_desc_4_attr_reg
    ,output reg [31:0] rd_req_desc_4_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_4_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_4_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_4_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_4_axid_0_reg
    ,output reg [31:0] rd_req_desc_4_axid_1_reg
    ,output reg [31:0] rd_req_desc_4_axid_2_reg
    ,output reg [31:0] rd_req_desc_4_axid_3_reg
    ,output reg [31:0] rd_req_desc_4_axuser_0_reg
    ,output reg [31:0] rd_req_desc_4_axuser_1_reg
    ,output reg [31:0] rd_req_desc_4_axuser_2_reg
    ,output reg [31:0] rd_req_desc_4_axuser_3_reg
    ,output reg [31:0] rd_req_desc_4_axuser_4_reg
    ,output reg [31:0] rd_req_desc_4_axuser_5_reg
    ,output reg [31:0] rd_req_desc_4_axuser_6_reg
    ,output reg [31:0] rd_req_desc_4_axuser_7_reg
    ,output reg [31:0] rd_req_desc_4_axuser_8_reg
    ,output reg [31:0] rd_req_desc_4_axuser_9_reg
    ,output reg [31:0] rd_req_desc_4_axuser_10_reg
    ,output reg [31:0] rd_req_desc_4_axuser_11_reg
    ,output reg [31:0] rd_req_desc_4_axuser_12_reg
    ,output reg [31:0] rd_req_desc_4_axuser_13_reg
    ,output reg [31:0] rd_req_desc_4_axuser_14_reg
    ,output reg [31:0] rd_req_desc_4_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_4_data_offset_reg
    ,output reg [31:0] rd_resp_desc_4_data_size_reg
    ,output reg [31:0] rd_resp_desc_4_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_4_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_4_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_4_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_4_resp_reg
    ,output reg [31:0] rd_resp_desc_4_xid_0_reg
    ,output reg [31:0] rd_resp_desc_4_xid_1_reg
    ,output reg [31:0] rd_resp_desc_4_xid_2_reg
    ,output reg [31:0] rd_resp_desc_4_xid_3_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_4_xuser_15_reg
    ,output reg [31:0] wr_req_desc_4_txn_type_reg
    ,output reg [31:0] wr_req_desc_4_size_reg
    ,output reg [31:0] wr_req_desc_4_data_offset_reg
    ,output reg [31:0] wr_req_desc_4_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_4_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_4_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_4_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_4_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_4_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_4_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_4_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_4_axsize_reg
    ,output reg [31:0] wr_req_desc_4_attr_reg
    ,output reg [31:0] wr_req_desc_4_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_4_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_4_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_4_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_4_axid_0_reg
    ,output reg [31:0] wr_req_desc_4_axid_1_reg
    ,output reg [31:0] wr_req_desc_4_axid_2_reg
    ,output reg [31:0] wr_req_desc_4_axid_3_reg
    ,output reg [31:0] wr_req_desc_4_axuser_0_reg
    ,output reg [31:0] wr_req_desc_4_axuser_1_reg
    ,output reg [31:0] wr_req_desc_4_axuser_2_reg
    ,output reg [31:0] wr_req_desc_4_axuser_3_reg
    ,output reg [31:0] wr_req_desc_4_axuser_4_reg
    ,output reg [31:0] wr_req_desc_4_axuser_5_reg
    ,output reg [31:0] wr_req_desc_4_axuser_6_reg
    ,output reg [31:0] wr_req_desc_4_axuser_7_reg
    ,output reg [31:0] wr_req_desc_4_axuser_8_reg
    ,output reg [31:0] wr_req_desc_4_axuser_9_reg
    ,output reg [31:0] wr_req_desc_4_axuser_10_reg
    ,output reg [31:0] wr_req_desc_4_axuser_11_reg
    ,output reg [31:0] wr_req_desc_4_axuser_12_reg
    ,output reg [31:0] wr_req_desc_4_axuser_13_reg
    ,output reg [31:0] wr_req_desc_4_axuser_14_reg
    ,output reg [31:0] wr_req_desc_4_axuser_15_reg
    ,output reg [31:0] wr_req_desc_4_wuser_0_reg
    ,output reg [31:0] wr_req_desc_4_wuser_1_reg
    ,output reg [31:0] wr_req_desc_4_wuser_2_reg
    ,output reg [31:0] wr_req_desc_4_wuser_3_reg
    ,output reg [31:0] wr_req_desc_4_wuser_4_reg
    ,output reg [31:0] wr_req_desc_4_wuser_5_reg
    ,output reg [31:0] wr_req_desc_4_wuser_6_reg
    ,output reg [31:0] wr_req_desc_4_wuser_7_reg
    ,output reg [31:0] wr_req_desc_4_wuser_8_reg
    ,output reg [31:0] wr_req_desc_4_wuser_9_reg
    ,output reg [31:0] wr_req_desc_4_wuser_10_reg
    ,output reg [31:0] wr_req_desc_4_wuser_11_reg
    ,output reg [31:0] wr_req_desc_4_wuser_12_reg
    ,output reg [31:0] wr_req_desc_4_wuser_13_reg
    ,output reg [31:0] wr_req_desc_4_wuser_14_reg
    ,output reg [31:0] wr_req_desc_4_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_4_resp_reg
    ,output reg [31:0] wr_resp_desc_4_xid_0_reg
    ,output reg [31:0] wr_resp_desc_4_xid_1_reg
    ,output reg [31:0] wr_resp_desc_4_xid_2_reg
    ,output reg [31:0] wr_resp_desc_4_xid_3_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_4_xuser_15_reg
    ,output reg [31:0] sn_req_desc_4_attr_reg
    ,output reg [31:0] sn_req_desc_4_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_4_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_4_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_4_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_4_resp_reg
    ,output reg [31:0] rd_req_desc_5_txn_type_reg
    ,output reg [31:0] rd_req_desc_5_size_reg
    ,output reg [31:0] rd_req_desc_5_axsize_reg
    ,output reg [31:0] rd_req_desc_5_attr_reg
    ,output reg [31:0] rd_req_desc_5_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_5_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_5_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_5_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_5_axid_0_reg
    ,output reg [31:0] rd_req_desc_5_axid_1_reg
    ,output reg [31:0] rd_req_desc_5_axid_2_reg
    ,output reg [31:0] rd_req_desc_5_axid_3_reg
    ,output reg [31:0] rd_req_desc_5_axuser_0_reg
    ,output reg [31:0] rd_req_desc_5_axuser_1_reg
    ,output reg [31:0] rd_req_desc_5_axuser_2_reg
    ,output reg [31:0] rd_req_desc_5_axuser_3_reg
    ,output reg [31:0] rd_req_desc_5_axuser_4_reg
    ,output reg [31:0] rd_req_desc_5_axuser_5_reg
    ,output reg [31:0] rd_req_desc_5_axuser_6_reg
    ,output reg [31:0] rd_req_desc_5_axuser_7_reg
    ,output reg [31:0] rd_req_desc_5_axuser_8_reg
    ,output reg [31:0] rd_req_desc_5_axuser_9_reg
    ,output reg [31:0] rd_req_desc_5_axuser_10_reg
    ,output reg [31:0] rd_req_desc_5_axuser_11_reg
    ,output reg [31:0] rd_req_desc_5_axuser_12_reg
    ,output reg [31:0] rd_req_desc_5_axuser_13_reg
    ,output reg [31:0] rd_req_desc_5_axuser_14_reg
    ,output reg [31:0] rd_req_desc_5_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_5_data_offset_reg
    ,output reg [31:0] rd_resp_desc_5_data_size_reg
    ,output reg [31:0] rd_resp_desc_5_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_5_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_5_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_5_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_5_resp_reg
    ,output reg [31:0] rd_resp_desc_5_xid_0_reg
    ,output reg [31:0] rd_resp_desc_5_xid_1_reg
    ,output reg [31:0] rd_resp_desc_5_xid_2_reg
    ,output reg [31:0] rd_resp_desc_5_xid_3_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_5_xuser_15_reg
    ,output reg [31:0] wr_req_desc_5_txn_type_reg
    ,output reg [31:0] wr_req_desc_5_size_reg
    ,output reg [31:0] wr_req_desc_5_data_offset_reg
    ,output reg [31:0] wr_req_desc_5_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_5_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_5_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_5_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_5_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_5_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_5_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_5_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_5_axsize_reg
    ,output reg [31:0] wr_req_desc_5_attr_reg
    ,output reg [31:0] wr_req_desc_5_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_5_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_5_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_5_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_5_axid_0_reg
    ,output reg [31:0] wr_req_desc_5_axid_1_reg
    ,output reg [31:0] wr_req_desc_5_axid_2_reg
    ,output reg [31:0] wr_req_desc_5_axid_3_reg
    ,output reg [31:0] wr_req_desc_5_axuser_0_reg
    ,output reg [31:0] wr_req_desc_5_axuser_1_reg
    ,output reg [31:0] wr_req_desc_5_axuser_2_reg
    ,output reg [31:0] wr_req_desc_5_axuser_3_reg
    ,output reg [31:0] wr_req_desc_5_axuser_4_reg
    ,output reg [31:0] wr_req_desc_5_axuser_5_reg
    ,output reg [31:0] wr_req_desc_5_axuser_6_reg
    ,output reg [31:0] wr_req_desc_5_axuser_7_reg
    ,output reg [31:0] wr_req_desc_5_axuser_8_reg
    ,output reg [31:0] wr_req_desc_5_axuser_9_reg
    ,output reg [31:0] wr_req_desc_5_axuser_10_reg
    ,output reg [31:0] wr_req_desc_5_axuser_11_reg
    ,output reg [31:0] wr_req_desc_5_axuser_12_reg
    ,output reg [31:0] wr_req_desc_5_axuser_13_reg
    ,output reg [31:0] wr_req_desc_5_axuser_14_reg
    ,output reg [31:0] wr_req_desc_5_axuser_15_reg
    ,output reg [31:0] wr_req_desc_5_wuser_0_reg
    ,output reg [31:0] wr_req_desc_5_wuser_1_reg
    ,output reg [31:0] wr_req_desc_5_wuser_2_reg
    ,output reg [31:0] wr_req_desc_5_wuser_3_reg
    ,output reg [31:0] wr_req_desc_5_wuser_4_reg
    ,output reg [31:0] wr_req_desc_5_wuser_5_reg
    ,output reg [31:0] wr_req_desc_5_wuser_6_reg
    ,output reg [31:0] wr_req_desc_5_wuser_7_reg
    ,output reg [31:0] wr_req_desc_5_wuser_8_reg
    ,output reg [31:0] wr_req_desc_5_wuser_9_reg
    ,output reg [31:0] wr_req_desc_5_wuser_10_reg
    ,output reg [31:0] wr_req_desc_5_wuser_11_reg
    ,output reg [31:0] wr_req_desc_5_wuser_12_reg
    ,output reg [31:0] wr_req_desc_5_wuser_13_reg
    ,output reg [31:0] wr_req_desc_5_wuser_14_reg
    ,output reg [31:0] wr_req_desc_5_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_5_resp_reg
    ,output reg [31:0] wr_resp_desc_5_xid_0_reg
    ,output reg [31:0] wr_resp_desc_5_xid_1_reg
    ,output reg [31:0] wr_resp_desc_5_xid_2_reg
    ,output reg [31:0] wr_resp_desc_5_xid_3_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_5_xuser_15_reg
    ,output reg [31:0] sn_req_desc_5_attr_reg
    ,output reg [31:0] sn_req_desc_5_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_5_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_5_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_5_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_5_resp_reg
    ,output reg [31:0] rd_req_desc_6_txn_type_reg
    ,output reg [31:0] rd_req_desc_6_size_reg
    ,output reg [31:0] rd_req_desc_6_axsize_reg
    ,output reg [31:0] rd_req_desc_6_attr_reg
    ,output reg [31:0] rd_req_desc_6_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_6_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_6_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_6_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_6_axid_0_reg
    ,output reg [31:0] rd_req_desc_6_axid_1_reg
    ,output reg [31:0] rd_req_desc_6_axid_2_reg
    ,output reg [31:0] rd_req_desc_6_axid_3_reg
    ,output reg [31:0] rd_req_desc_6_axuser_0_reg
    ,output reg [31:0] rd_req_desc_6_axuser_1_reg
    ,output reg [31:0] rd_req_desc_6_axuser_2_reg
    ,output reg [31:0] rd_req_desc_6_axuser_3_reg
    ,output reg [31:0] rd_req_desc_6_axuser_4_reg
    ,output reg [31:0] rd_req_desc_6_axuser_5_reg
    ,output reg [31:0] rd_req_desc_6_axuser_6_reg
    ,output reg [31:0] rd_req_desc_6_axuser_7_reg
    ,output reg [31:0] rd_req_desc_6_axuser_8_reg
    ,output reg [31:0] rd_req_desc_6_axuser_9_reg
    ,output reg [31:0] rd_req_desc_6_axuser_10_reg
    ,output reg [31:0] rd_req_desc_6_axuser_11_reg
    ,output reg [31:0] rd_req_desc_6_axuser_12_reg
    ,output reg [31:0] rd_req_desc_6_axuser_13_reg
    ,output reg [31:0] rd_req_desc_6_axuser_14_reg
    ,output reg [31:0] rd_req_desc_6_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_6_data_offset_reg
    ,output reg [31:0] rd_resp_desc_6_data_size_reg
    ,output reg [31:0] rd_resp_desc_6_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_6_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_6_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_6_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_6_resp_reg
    ,output reg [31:0] rd_resp_desc_6_xid_0_reg
    ,output reg [31:0] rd_resp_desc_6_xid_1_reg
    ,output reg [31:0] rd_resp_desc_6_xid_2_reg
    ,output reg [31:0] rd_resp_desc_6_xid_3_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_6_xuser_15_reg
    ,output reg [31:0] wr_req_desc_6_txn_type_reg
    ,output reg [31:0] wr_req_desc_6_size_reg
    ,output reg [31:0] wr_req_desc_6_data_offset_reg
    ,output reg [31:0] wr_req_desc_6_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_6_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_6_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_6_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_6_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_6_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_6_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_6_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_6_axsize_reg
    ,output reg [31:0] wr_req_desc_6_attr_reg
    ,output reg [31:0] wr_req_desc_6_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_6_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_6_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_6_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_6_axid_0_reg
    ,output reg [31:0] wr_req_desc_6_axid_1_reg
    ,output reg [31:0] wr_req_desc_6_axid_2_reg
    ,output reg [31:0] wr_req_desc_6_axid_3_reg
    ,output reg [31:0] wr_req_desc_6_axuser_0_reg
    ,output reg [31:0] wr_req_desc_6_axuser_1_reg
    ,output reg [31:0] wr_req_desc_6_axuser_2_reg
    ,output reg [31:0] wr_req_desc_6_axuser_3_reg
    ,output reg [31:0] wr_req_desc_6_axuser_4_reg
    ,output reg [31:0] wr_req_desc_6_axuser_5_reg
    ,output reg [31:0] wr_req_desc_6_axuser_6_reg
    ,output reg [31:0] wr_req_desc_6_axuser_7_reg
    ,output reg [31:0] wr_req_desc_6_axuser_8_reg
    ,output reg [31:0] wr_req_desc_6_axuser_9_reg
    ,output reg [31:0] wr_req_desc_6_axuser_10_reg
    ,output reg [31:0] wr_req_desc_6_axuser_11_reg
    ,output reg [31:0] wr_req_desc_6_axuser_12_reg
    ,output reg [31:0] wr_req_desc_6_axuser_13_reg
    ,output reg [31:0] wr_req_desc_6_axuser_14_reg
    ,output reg [31:0] wr_req_desc_6_axuser_15_reg
    ,output reg [31:0] wr_req_desc_6_wuser_0_reg
    ,output reg [31:0] wr_req_desc_6_wuser_1_reg
    ,output reg [31:0] wr_req_desc_6_wuser_2_reg
    ,output reg [31:0] wr_req_desc_6_wuser_3_reg
    ,output reg [31:0] wr_req_desc_6_wuser_4_reg
    ,output reg [31:0] wr_req_desc_6_wuser_5_reg
    ,output reg [31:0] wr_req_desc_6_wuser_6_reg
    ,output reg [31:0] wr_req_desc_6_wuser_7_reg
    ,output reg [31:0] wr_req_desc_6_wuser_8_reg
    ,output reg [31:0] wr_req_desc_6_wuser_9_reg
    ,output reg [31:0] wr_req_desc_6_wuser_10_reg
    ,output reg [31:0] wr_req_desc_6_wuser_11_reg
    ,output reg [31:0] wr_req_desc_6_wuser_12_reg
    ,output reg [31:0] wr_req_desc_6_wuser_13_reg
    ,output reg [31:0] wr_req_desc_6_wuser_14_reg
    ,output reg [31:0] wr_req_desc_6_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_6_resp_reg
    ,output reg [31:0] wr_resp_desc_6_xid_0_reg
    ,output reg [31:0] wr_resp_desc_6_xid_1_reg
    ,output reg [31:0] wr_resp_desc_6_xid_2_reg
    ,output reg [31:0] wr_resp_desc_6_xid_3_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_6_xuser_15_reg
    ,output reg [31:0] sn_req_desc_6_attr_reg
    ,output reg [31:0] sn_req_desc_6_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_6_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_6_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_6_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_6_resp_reg
    ,output reg [31:0] rd_req_desc_7_txn_type_reg
    ,output reg [31:0] rd_req_desc_7_size_reg
    ,output reg [31:0] rd_req_desc_7_axsize_reg
    ,output reg [31:0] rd_req_desc_7_attr_reg
    ,output reg [31:0] rd_req_desc_7_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_7_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_7_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_7_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_7_axid_0_reg
    ,output reg [31:0] rd_req_desc_7_axid_1_reg
    ,output reg [31:0] rd_req_desc_7_axid_2_reg
    ,output reg [31:0] rd_req_desc_7_axid_3_reg
    ,output reg [31:0] rd_req_desc_7_axuser_0_reg
    ,output reg [31:0] rd_req_desc_7_axuser_1_reg
    ,output reg [31:0] rd_req_desc_7_axuser_2_reg
    ,output reg [31:0] rd_req_desc_7_axuser_3_reg
    ,output reg [31:0] rd_req_desc_7_axuser_4_reg
    ,output reg [31:0] rd_req_desc_7_axuser_5_reg
    ,output reg [31:0] rd_req_desc_7_axuser_6_reg
    ,output reg [31:0] rd_req_desc_7_axuser_7_reg
    ,output reg [31:0] rd_req_desc_7_axuser_8_reg
    ,output reg [31:0] rd_req_desc_7_axuser_9_reg
    ,output reg [31:0] rd_req_desc_7_axuser_10_reg
    ,output reg [31:0] rd_req_desc_7_axuser_11_reg
    ,output reg [31:0] rd_req_desc_7_axuser_12_reg
    ,output reg [31:0] rd_req_desc_7_axuser_13_reg
    ,output reg [31:0] rd_req_desc_7_axuser_14_reg
    ,output reg [31:0] rd_req_desc_7_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_7_data_offset_reg
    ,output reg [31:0] rd_resp_desc_7_data_size_reg
    ,output reg [31:0] rd_resp_desc_7_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_7_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_7_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_7_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_7_resp_reg
    ,output reg [31:0] rd_resp_desc_7_xid_0_reg
    ,output reg [31:0] rd_resp_desc_7_xid_1_reg
    ,output reg [31:0] rd_resp_desc_7_xid_2_reg
    ,output reg [31:0] rd_resp_desc_7_xid_3_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_7_xuser_15_reg
    ,output reg [31:0] wr_req_desc_7_txn_type_reg
    ,output reg [31:0] wr_req_desc_7_size_reg
    ,output reg [31:0] wr_req_desc_7_data_offset_reg
    ,output reg [31:0] wr_req_desc_7_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_7_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_7_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_7_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_7_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_7_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_7_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_7_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_7_axsize_reg
    ,output reg [31:0] wr_req_desc_7_attr_reg
    ,output reg [31:0] wr_req_desc_7_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_7_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_7_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_7_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_7_axid_0_reg
    ,output reg [31:0] wr_req_desc_7_axid_1_reg
    ,output reg [31:0] wr_req_desc_7_axid_2_reg
    ,output reg [31:0] wr_req_desc_7_axid_3_reg
    ,output reg [31:0] wr_req_desc_7_axuser_0_reg
    ,output reg [31:0] wr_req_desc_7_axuser_1_reg
    ,output reg [31:0] wr_req_desc_7_axuser_2_reg
    ,output reg [31:0] wr_req_desc_7_axuser_3_reg
    ,output reg [31:0] wr_req_desc_7_axuser_4_reg
    ,output reg [31:0] wr_req_desc_7_axuser_5_reg
    ,output reg [31:0] wr_req_desc_7_axuser_6_reg
    ,output reg [31:0] wr_req_desc_7_axuser_7_reg
    ,output reg [31:0] wr_req_desc_7_axuser_8_reg
    ,output reg [31:0] wr_req_desc_7_axuser_9_reg
    ,output reg [31:0] wr_req_desc_7_axuser_10_reg
    ,output reg [31:0] wr_req_desc_7_axuser_11_reg
    ,output reg [31:0] wr_req_desc_7_axuser_12_reg
    ,output reg [31:0] wr_req_desc_7_axuser_13_reg
    ,output reg [31:0] wr_req_desc_7_axuser_14_reg
    ,output reg [31:0] wr_req_desc_7_axuser_15_reg
    ,output reg [31:0] wr_req_desc_7_wuser_0_reg
    ,output reg [31:0] wr_req_desc_7_wuser_1_reg
    ,output reg [31:0] wr_req_desc_7_wuser_2_reg
    ,output reg [31:0] wr_req_desc_7_wuser_3_reg
    ,output reg [31:0] wr_req_desc_7_wuser_4_reg
    ,output reg [31:0] wr_req_desc_7_wuser_5_reg
    ,output reg [31:0] wr_req_desc_7_wuser_6_reg
    ,output reg [31:0] wr_req_desc_7_wuser_7_reg
    ,output reg [31:0] wr_req_desc_7_wuser_8_reg
    ,output reg [31:0] wr_req_desc_7_wuser_9_reg
    ,output reg [31:0] wr_req_desc_7_wuser_10_reg
    ,output reg [31:0] wr_req_desc_7_wuser_11_reg
    ,output reg [31:0] wr_req_desc_7_wuser_12_reg
    ,output reg [31:0] wr_req_desc_7_wuser_13_reg
    ,output reg [31:0] wr_req_desc_7_wuser_14_reg
    ,output reg [31:0] wr_req_desc_7_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_7_resp_reg
    ,output reg [31:0] wr_resp_desc_7_xid_0_reg
    ,output reg [31:0] wr_resp_desc_7_xid_1_reg
    ,output reg [31:0] wr_resp_desc_7_xid_2_reg
    ,output reg [31:0] wr_resp_desc_7_xid_3_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_7_xuser_15_reg
    ,output reg [31:0] sn_req_desc_7_attr_reg
    ,output reg [31:0] sn_req_desc_7_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_7_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_7_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_7_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_7_resp_reg
    ,output reg [31:0] rd_req_desc_8_txn_type_reg
    ,output reg [31:0] rd_req_desc_8_size_reg
    ,output reg [31:0] rd_req_desc_8_axsize_reg
    ,output reg [31:0] rd_req_desc_8_attr_reg
    ,output reg [31:0] rd_req_desc_8_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_8_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_8_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_8_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_8_axid_0_reg
    ,output reg [31:0] rd_req_desc_8_axid_1_reg
    ,output reg [31:0] rd_req_desc_8_axid_2_reg
    ,output reg [31:0] rd_req_desc_8_axid_3_reg
    ,output reg [31:0] rd_req_desc_8_axuser_0_reg
    ,output reg [31:0] rd_req_desc_8_axuser_1_reg
    ,output reg [31:0] rd_req_desc_8_axuser_2_reg
    ,output reg [31:0] rd_req_desc_8_axuser_3_reg
    ,output reg [31:0] rd_req_desc_8_axuser_4_reg
    ,output reg [31:0] rd_req_desc_8_axuser_5_reg
    ,output reg [31:0] rd_req_desc_8_axuser_6_reg
    ,output reg [31:0] rd_req_desc_8_axuser_7_reg
    ,output reg [31:0] rd_req_desc_8_axuser_8_reg
    ,output reg [31:0] rd_req_desc_8_axuser_9_reg
    ,output reg [31:0] rd_req_desc_8_axuser_10_reg
    ,output reg [31:0] rd_req_desc_8_axuser_11_reg
    ,output reg [31:0] rd_req_desc_8_axuser_12_reg
    ,output reg [31:0] rd_req_desc_8_axuser_13_reg
    ,output reg [31:0] rd_req_desc_8_axuser_14_reg
    ,output reg [31:0] rd_req_desc_8_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_8_data_offset_reg
    ,output reg [31:0] rd_resp_desc_8_data_size_reg
    ,output reg [31:0] rd_resp_desc_8_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_8_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_8_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_8_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_8_resp_reg
    ,output reg [31:0] rd_resp_desc_8_xid_0_reg
    ,output reg [31:0] rd_resp_desc_8_xid_1_reg
    ,output reg [31:0] rd_resp_desc_8_xid_2_reg
    ,output reg [31:0] rd_resp_desc_8_xid_3_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_8_xuser_15_reg
    ,output reg [31:0] wr_req_desc_8_txn_type_reg
    ,output reg [31:0] wr_req_desc_8_size_reg
    ,output reg [31:0] wr_req_desc_8_data_offset_reg
    ,output reg [31:0] wr_req_desc_8_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_8_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_8_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_8_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_8_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_8_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_8_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_8_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_8_axsize_reg
    ,output reg [31:0] wr_req_desc_8_attr_reg
    ,output reg [31:0] wr_req_desc_8_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_8_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_8_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_8_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_8_axid_0_reg
    ,output reg [31:0] wr_req_desc_8_axid_1_reg
    ,output reg [31:0] wr_req_desc_8_axid_2_reg
    ,output reg [31:0] wr_req_desc_8_axid_3_reg
    ,output reg [31:0] wr_req_desc_8_axuser_0_reg
    ,output reg [31:0] wr_req_desc_8_axuser_1_reg
    ,output reg [31:0] wr_req_desc_8_axuser_2_reg
    ,output reg [31:0] wr_req_desc_8_axuser_3_reg
    ,output reg [31:0] wr_req_desc_8_axuser_4_reg
    ,output reg [31:0] wr_req_desc_8_axuser_5_reg
    ,output reg [31:0] wr_req_desc_8_axuser_6_reg
    ,output reg [31:0] wr_req_desc_8_axuser_7_reg
    ,output reg [31:0] wr_req_desc_8_axuser_8_reg
    ,output reg [31:0] wr_req_desc_8_axuser_9_reg
    ,output reg [31:0] wr_req_desc_8_axuser_10_reg
    ,output reg [31:0] wr_req_desc_8_axuser_11_reg
    ,output reg [31:0] wr_req_desc_8_axuser_12_reg
    ,output reg [31:0] wr_req_desc_8_axuser_13_reg
    ,output reg [31:0] wr_req_desc_8_axuser_14_reg
    ,output reg [31:0] wr_req_desc_8_axuser_15_reg
    ,output reg [31:0] wr_req_desc_8_wuser_0_reg
    ,output reg [31:0] wr_req_desc_8_wuser_1_reg
    ,output reg [31:0] wr_req_desc_8_wuser_2_reg
    ,output reg [31:0] wr_req_desc_8_wuser_3_reg
    ,output reg [31:0] wr_req_desc_8_wuser_4_reg
    ,output reg [31:0] wr_req_desc_8_wuser_5_reg
    ,output reg [31:0] wr_req_desc_8_wuser_6_reg
    ,output reg [31:0] wr_req_desc_8_wuser_7_reg
    ,output reg [31:0] wr_req_desc_8_wuser_8_reg
    ,output reg [31:0] wr_req_desc_8_wuser_9_reg
    ,output reg [31:0] wr_req_desc_8_wuser_10_reg
    ,output reg [31:0] wr_req_desc_8_wuser_11_reg
    ,output reg [31:0] wr_req_desc_8_wuser_12_reg
    ,output reg [31:0] wr_req_desc_8_wuser_13_reg
    ,output reg [31:0] wr_req_desc_8_wuser_14_reg
    ,output reg [31:0] wr_req_desc_8_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_8_resp_reg
    ,output reg [31:0] wr_resp_desc_8_xid_0_reg
    ,output reg [31:0] wr_resp_desc_8_xid_1_reg
    ,output reg [31:0] wr_resp_desc_8_xid_2_reg
    ,output reg [31:0] wr_resp_desc_8_xid_3_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_8_xuser_15_reg
    ,output reg [31:0] sn_req_desc_8_attr_reg
    ,output reg [31:0] sn_req_desc_8_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_8_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_8_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_8_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_8_resp_reg
    ,output reg [31:0] rd_req_desc_9_txn_type_reg
    ,output reg [31:0] rd_req_desc_9_size_reg
    ,output reg [31:0] rd_req_desc_9_axsize_reg
    ,output reg [31:0] rd_req_desc_9_attr_reg
    ,output reg [31:0] rd_req_desc_9_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_9_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_9_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_9_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_9_axid_0_reg
    ,output reg [31:0] rd_req_desc_9_axid_1_reg
    ,output reg [31:0] rd_req_desc_9_axid_2_reg
    ,output reg [31:0] rd_req_desc_9_axid_3_reg
    ,output reg [31:0] rd_req_desc_9_axuser_0_reg
    ,output reg [31:0] rd_req_desc_9_axuser_1_reg
    ,output reg [31:0] rd_req_desc_9_axuser_2_reg
    ,output reg [31:0] rd_req_desc_9_axuser_3_reg
    ,output reg [31:0] rd_req_desc_9_axuser_4_reg
    ,output reg [31:0] rd_req_desc_9_axuser_5_reg
    ,output reg [31:0] rd_req_desc_9_axuser_6_reg
    ,output reg [31:0] rd_req_desc_9_axuser_7_reg
    ,output reg [31:0] rd_req_desc_9_axuser_8_reg
    ,output reg [31:0] rd_req_desc_9_axuser_9_reg
    ,output reg [31:0] rd_req_desc_9_axuser_10_reg
    ,output reg [31:0] rd_req_desc_9_axuser_11_reg
    ,output reg [31:0] rd_req_desc_9_axuser_12_reg
    ,output reg [31:0] rd_req_desc_9_axuser_13_reg
    ,output reg [31:0] rd_req_desc_9_axuser_14_reg
    ,output reg [31:0] rd_req_desc_9_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_9_data_offset_reg
    ,output reg [31:0] rd_resp_desc_9_data_size_reg
    ,output reg [31:0] rd_resp_desc_9_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_9_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_9_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_9_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_9_resp_reg
    ,output reg [31:0] rd_resp_desc_9_xid_0_reg
    ,output reg [31:0] rd_resp_desc_9_xid_1_reg
    ,output reg [31:0] rd_resp_desc_9_xid_2_reg
    ,output reg [31:0] rd_resp_desc_9_xid_3_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_9_xuser_15_reg
    ,output reg [31:0] wr_req_desc_9_txn_type_reg
    ,output reg [31:0] wr_req_desc_9_size_reg
    ,output reg [31:0] wr_req_desc_9_data_offset_reg
    ,output reg [31:0] wr_req_desc_9_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_9_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_9_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_9_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_9_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_9_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_9_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_9_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_9_axsize_reg
    ,output reg [31:0] wr_req_desc_9_attr_reg
    ,output reg [31:0] wr_req_desc_9_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_9_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_9_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_9_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_9_axid_0_reg
    ,output reg [31:0] wr_req_desc_9_axid_1_reg
    ,output reg [31:0] wr_req_desc_9_axid_2_reg
    ,output reg [31:0] wr_req_desc_9_axid_3_reg
    ,output reg [31:0] wr_req_desc_9_axuser_0_reg
    ,output reg [31:0] wr_req_desc_9_axuser_1_reg
    ,output reg [31:0] wr_req_desc_9_axuser_2_reg
    ,output reg [31:0] wr_req_desc_9_axuser_3_reg
    ,output reg [31:0] wr_req_desc_9_axuser_4_reg
    ,output reg [31:0] wr_req_desc_9_axuser_5_reg
    ,output reg [31:0] wr_req_desc_9_axuser_6_reg
    ,output reg [31:0] wr_req_desc_9_axuser_7_reg
    ,output reg [31:0] wr_req_desc_9_axuser_8_reg
    ,output reg [31:0] wr_req_desc_9_axuser_9_reg
    ,output reg [31:0] wr_req_desc_9_axuser_10_reg
    ,output reg [31:0] wr_req_desc_9_axuser_11_reg
    ,output reg [31:0] wr_req_desc_9_axuser_12_reg
    ,output reg [31:0] wr_req_desc_9_axuser_13_reg
    ,output reg [31:0] wr_req_desc_9_axuser_14_reg
    ,output reg [31:0] wr_req_desc_9_axuser_15_reg
    ,output reg [31:0] wr_req_desc_9_wuser_0_reg
    ,output reg [31:0] wr_req_desc_9_wuser_1_reg
    ,output reg [31:0] wr_req_desc_9_wuser_2_reg
    ,output reg [31:0] wr_req_desc_9_wuser_3_reg
    ,output reg [31:0] wr_req_desc_9_wuser_4_reg
    ,output reg [31:0] wr_req_desc_9_wuser_5_reg
    ,output reg [31:0] wr_req_desc_9_wuser_6_reg
    ,output reg [31:0] wr_req_desc_9_wuser_7_reg
    ,output reg [31:0] wr_req_desc_9_wuser_8_reg
    ,output reg [31:0] wr_req_desc_9_wuser_9_reg
    ,output reg [31:0] wr_req_desc_9_wuser_10_reg
    ,output reg [31:0] wr_req_desc_9_wuser_11_reg
    ,output reg [31:0] wr_req_desc_9_wuser_12_reg
    ,output reg [31:0] wr_req_desc_9_wuser_13_reg
    ,output reg [31:0] wr_req_desc_9_wuser_14_reg
    ,output reg [31:0] wr_req_desc_9_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_9_resp_reg
    ,output reg [31:0] wr_resp_desc_9_xid_0_reg
    ,output reg [31:0] wr_resp_desc_9_xid_1_reg
    ,output reg [31:0] wr_resp_desc_9_xid_2_reg
    ,output reg [31:0] wr_resp_desc_9_xid_3_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_9_xuser_15_reg
    ,output reg [31:0] sn_req_desc_9_attr_reg
    ,output reg [31:0] sn_req_desc_9_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_9_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_9_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_9_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_9_resp_reg
    ,output reg [31:0] rd_req_desc_a_txn_type_reg
    ,output reg [31:0] rd_req_desc_a_size_reg
    ,output reg [31:0] rd_req_desc_a_axsize_reg
    ,output reg [31:0] rd_req_desc_a_attr_reg
    ,output reg [31:0] rd_req_desc_a_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_a_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_a_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_a_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_a_axid_0_reg
    ,output reg [31:0] rd_req_desc_a_axid_1_reg
    ,output reg [31:0] rd_req_desc_a_axid_2_reg
    ,output reg [31:0] rd_req_desc_a_axid_3_reg
    ,output reg [31:0] rd_req_desc_a_axuser_0_reg
    ,output reg [31:0] rd_req_desc_a_axuser_1_reg
    ,output reg [31:0] rd_req_desc_a_axuser_2_reg
    ,output reg [31:0] rd_req_desc_a_axuser_3_reg
    ,output reg [31:0] rd_req_desc_a_axuser_4_reg
    ,output reg [31:0] rd_req_desc_a_axuser_5_reg
    ,output reg [31:0] rd_req_desc_a_axuser_6_reg
    ,output reg [31:0] rd_req_desc_a_axuser_7_reg
    ,output reg [31:0] rd_req_desc_a_axuser_8_reg
    ,output reg [31:0] rd_req_desc_a_axuser_9_reg
    ,output reg [31:0] rd_req_desc_a_axuser_10_reg
    ,output reg [31:0] rd_req_desc_a_axuser_11_reg
    ,output reg [31:0] rd_req_desc_a_axuser_12_reg
    ,output reg [31:0] rd_req_desc_a_axuser_13_reg
    ,output reg [31:0] rd_req_desc_a_axuser_14_reg
    ,output reg [31:0] rd_req_desc_a_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_a_data_offset_reg
    ,output reg [31:0] rd_resp_desc_a_data_size_reg
    ,output reg [31:0] rd_resp_desc_a_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_a_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_a_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_a_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_a_resp_reg
    ,output reg [31:0] rd_resp_desc_a_xid_0_reg
    ,output reg [31:0] rd_resp_desc_a_xid_1_reg
    ,output reg [31:0] rd_resp_desc_a_xid_2_reg
    ,output reg [31:0] rd_resp_desc_a_xid_3_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_a_xuser_15_reg
    ,output reg [31:0] wr_req_desc_a_txn_type_reg
    ,output reg [31:0] wr_req_desc_a_size_reg
    ,output reg [31:0] wr_req_desc_a_data_offset_reg
    ,output reg [31:0] wr_req_desc_a_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_a_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_a_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_a_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_a_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_a_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_a_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_a_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_a_axsize_reg
    ,output reg [31:0] wr_req_desc_a_attr_reg
    ,output reg [31:0] wr_req_desc_a_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_a_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_a_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_a_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_a_axid_0_reg
    ,output reg [31:0] wr_req_desc_a_axid_1_reg
    ,output reg [31:0] wr_req_desc_a_axid_2_reg
    ,output reg [31:0] wr_req_desc_a_axid_3_reg
    ,output reg [31:0] wr_req_desc_a_axuser_0_reg
    ,output reg [31:0] wr_req_desc_a_axuser_1_reg
    ,output reg [31:0] wr_req_desc_a_axuser_2_reg
    ,output reg [31:0] wr_req_desc_a_axuser_3_reg
    ,output reg [31:0] wr_req_desc_a_axuser_4_reg
    ,output reg [31:0] wr_req_desc_a_axuser_5_reg
    ,output reg [31:0] wr_req_desc_a_axuser_6_reg
    ,output reg [31:0] wr_req_desc_a_axuser_7_reg
    ,output reg [31:0] wr_req_desc_a_axuser_8_reg
    ,output reg [31:0] wr_req_desc_a_axuser_9_reg
    ,output reg [31:0] wr_req_desc_a_axuser_10_reg
    ,output reg [31:0] wr_req_desc_a_axuser_11_reg
    ,output reg [31:0] wr_req_desc_a_axuser_12_reg
    ,output reg [31:0] wr_req_desc_a_axuser_13_reg
    ,output reg [31:0] wr_req_desc_a_axuser_14_reg
    ,output reg [31:0] wr_req_desc_a_axuser_15_reg
    ,output reg [31:0] wr_req_desc_a_wuser_0_reg
    ,output reg [31:0] wr_req_desc_a_wuser_1_reg
    ,output reg [31:0] wr_req_desc_a_wuser_2_reg
    ,output reg [31:0] wr_req_desc_a_wuser_3_reg
    ,output reg [31:0] wr_req_desc_a_wuser_4_reg
    ,output reg [31:0] wr_req_desc_a_wuser_5_reg
    ,output reg [31:0] wr_req_desc_a_wuser_6_reg
    ,output reg [31:0] wr_req_desc_a_wuser_7_reg
    ,output reg [31:0] wr_req_desc_a_wuser_8_reg
    ,output reg [31:0] wr_req_desc_a_wuser_9_reg
    ,output reg [31:0] wr_req_desc_a_wuser_10_reg
    ,output reg [31:0] wr_req_desc_a_wuser_11_reg
    ,output reg [31:0] wr_req_desc_a_wuser_12_reg
    ,output reg [31:0] wr_req_desc_a_wuser_13_reg
    ,output reg [31:0] wr_req_desc_a_wuser_14_reg
    ,output reg [31:0] wr_req_desc_a_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_a_resp_reg
    ,output reg [31:0] wr_resp_desc_a_xid_0_reg
    ,output reg [31:0] wr_resp_desc_a_xid_1_reg
    ,output reg [31:0] wr_resp_desc_a_xid_2_reg
    ,output reg [31:0] wr_resp_desc_a_xid_3_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_a_xuser_15_reg
    ,output reg [31:0] sn_req_desc_a_attr_reg
    ,output reg [31:0] sn_req_desc_a_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_a_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_a_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_a_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_a_resp_reg
    ,output reg [31:0] rd_req_desc_b_txn_type_reg
    ,output reg [31:0] rd_req_desc_b_size_reg
    ,output reg [31:0] rd_req_desc_b_axsize_reg
    ,output reg [31:0] rd_req_desc_b_attr_reg
    ,output reg [31:0] rd_req_desc_b_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_b_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_b_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_b_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_b_axid_0_reg
    ,output reg [31:0] rd_req_desc_b_axid_1_reg
    ,output reg [31:0] rd_req_desc_b_axid_2_reg
    ,output reg [31:0] rd_req_desc_b_axid_3_reg
    ,output reg [31:0] rd_req_desc_b_axuser_0_reg
    ,output reg [31:0] rd_req_desc_b_axuser_1_reg
    ,output reg [31:0] rd_req_desc_b_axuser_2_reg
    ,output reg [31:0] rd_req_desc_b_axuser_3_reg
    ,output reg [31:0] rd_req_desc_b_axuser_4_reg
    ,output reg [31:0] rd_req_desc_b_axuser_5_reg
    ,output reg [31:0] rd_req_desc_b_axuser_6_reg
    ,output reg [31:0] rd_req_desc_b_axuser_7_reg
    ,output reg [31:0] rd_req_desc_b_axuser_8_reg
    ,output reg [31:0] rd_req_desc_b_axuser_9_reg
    ,output reg [31:0] rd_req_desc_b_axuser_10_reg
    ,output reg [31:0] rd_req_desc_b_axuser_11_reg
    ,output reg [31:0] rd_req_desc_b_axuser_12_reg
    ,output reg [31:0] rd_req_desc_b_axuser_13_reg
    ,output reg [31:0] rd_req_desc_b_axuser_14_reg
    ,output reg [31:0] rd_req_desc_b_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_b_data_offset_reg
    ,output reg [31:0] rd_resp_desc_b_data_size_reg
    ,output reg [31:0] rd_resp_desc_b_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_b_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_b_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_b_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_b_resp_reg
    ,output reg [31:0] rd_resp_desc_b_xid_0_reg
    ,output reg [31:0] rd_resp_desc_b_xid_1_reg
    ,output reg [31:0] rd_resp_desc_b_xid_2_reg
    ,output reg [31:0] rd_resp_desc_b_xid_3_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_b_xuser_15_reg
    ,output reg [31:0] wr_req_desc_b_txn_type_reg
    ,output reg [31:0] wr_req_desc_b_size_reg
    ,output reg [31:0] wr_req_desc_b_data_offset_reg
    ,output reg [31:0] wr_req_desc_b_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_b_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_b_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_b_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_b_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_b_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_b_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_b_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_b_axsize_reg
    ,output reg [31:0] wr_req_desc_b_attr_reg
    ,output reg [31:0] wr_req_desc_b_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_b_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_b_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_b_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_b_axid_0_reg
    ,output reg [31:0] wr_req_desc_b_axid_1_reg
    ,output reg [31:0] wr_req_desc_b_axid_2_reg
    ,output reg [31:0] wr_req_desc_b_axid_3_reg
    ,output reg [31:0] wr_req_desc_b_axuser_0_reg
    ,output reg [31:0] wr_req_desc_b_axuser_1_reg
    ,output reg [31:0] wr_req_desc_b_axuser_2_reg
    ,output reg [31:0] wr_req_desc_b_axuser_3_reg
    ,output reg [31:0] wr_req_desc_b_axuser_4_reg
    ,output reg [31:0] wr_req_desc_b_axuser_5_reg
    ,output reg [31:0] wr_req_desc_b_axuser_6_reg
    ,output reg [31:0] wr_req_desc_b_axuser_7_reg
    ,output reg [31:0] wr_req_desc_b_axuser_8_reg
    ,output reg [31:0] wr_req_desc_b_axuser_9_reg
    ,output reg [31:0] wr_req_desc_b_axuser_10_reg
    ,output reg [31:0] wr_req_desc_b_axuser_11_reg
    ,output reg [31:0] wr_req_desc_b_axuser_12_reg
    ,output reg [31:0] wr_req_desc_b_axuser_13_reg
    ,output reg [31:0] wr_req_desc_b_axuser_14_reg
    ,output reg [31:0] wr_req_desc_b_axuser_15_reg
    ,output reg [31:0] wr_req_desc_b_wuser_0_reg
    ,output reg [31:0] wr_req_desc_b_wuser_1_reg
    ,output reg [31:0] wr_req_desc_b_wuser_2_reg
    ,output reg [31:0] wr_req_desc_b_wuser_3_reg
    ,output reg [31:0] wr_req_desc_b_wuser_4_reg
    ,output reg [31:0] wr_req_desc_b_wuser_5_reg
    ,output reg [31:0] wr_req_desc_b_wuser_6_reg
    ,output reg [31:0] wr_req_desc_b_wuser_7_reg
    ,output reg [31:0] wr_req_desc_b_wuser_8_reg
    ,output reg [31:0] wr_req_desc_b_wuser_9_reg
    ,output reg [31:0] wr_req_desc_b_wuser_10_reg
    ,output reg [31:0] wr_req_desc_b_wuser_11_reg
    ,output reg [31:0] wr_req_desc_b_wuser_12_reg
    ,output reg [31:0] wr_req_desc_b_wuser_13_reg
    ,output reg [31:0] wr_req_desc_b_wuser_14_reg
    ,output reg [31:0] wr_req_desc_b_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_b_resp_reg
    ,output reg [31:0] wr_resp_desc_b_xid_0_reg
    ,output reg [31:0] wr_resp_desc_b_xid_1_reg
    ,output reg [31:0] wr_resp_desc_b_xid_2_reg
    ,output reg [31:0] wr_resp_desc_b_xid_3_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_b_xuser_15_reg
    ,output reg [31:0] sn_req_desc_b_attr_reg
    ,output reg [31:0] sn_req_desc_b_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_b_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_b_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_b_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_b_resp_reg
    ,output reg [31:0] rd_req_desc_c_txn_type_reg
    ,output reg [31:0] rd_req_desc_c_size_reg
    ,output reg [31:0] rd_req_desc_c_axsize_reg
    ,output reg [31:0] rd_req_desc_c_attr_reg
    ,output reg [31:0] rd_req_desc_c_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_c_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_c_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_c_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_c_axid_0_reg
    ,output reg [31:0] rd_req_desc_c_axid_1_reg
    ,output reg [31:0] rd_req_desc_c_axid_2_reg
    ,output reg [31:0] rd_req_desc_c_axid_3_reg
    ,output reg [31:0] rd_req_desc_c_axuser_0_reg
    ,output reg [31:0] rd_req_desc_c_axuser_1_reg
    ,output reg [31:0] rd_req_desc_c_axuser_2_reg
    ,output reg [31:0] rd_req_desc_c_axuser_3_reg
    ,output reg [31:0] rd_req_desc_c_axuser_4_reg
    ,output reg [31:0] rd_req_desc_c_axuser_5_reg
    ,output reg [31:0] rd_req_desc_c_axuser_6_reg
    ,output reg [31:0] rd_req_desc_c_axuser_7_reg
    ,output reg [31:0] rd_req_desc_c_axuser_8_reg
    ,output reg [31:0] rd_req_desc_c_axuser_9_reg
    ,output reg [31:0] rd_req_desc_c_axuser_10_reg
    ,output reg [31:0] rd_req_desc_c_axuser_11_reg
    ,output reg [31:0] rd_req_desc_c_axuser_12_reg
    ,output reg [31:0] rd_req_desc_c_axuser_13_reg
    ,output reg [31:0] rd_req_desc_c_axuser_14_reg
    ,output reg [31:0] rd_req_desc_c_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_c_data_offset_reg
    ,output reg [31:0] rd_resp_desc_c_data_size_reg
    ,output reg [31:0] rd_resp_desc_c_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_c_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_c_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_c_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_c_resp_reg
    ,output reg [31:0] rd_resp_desc_c_xid_0_reg
    ,output reg [31:0] rd_resp_desc_c_xid_1_reg
    ,output reg [31:0] rd_resp_desc_c_xid_2_reg
    ,output reg [31:0] rd_resp_desc_c_xid_3_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_c_xuser_15_reg
    ,output reg [31:0] wr_req_desc_c_txn_type_reg
    ,output reg [31:0] wr_req_desc_c_size_reg
    ,output reg [31:0] wr_req_desc_c_data_offset_reg
    ,output reg [31:0] wr_req_desc_c_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_c_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_c_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_c_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_c_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_c_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_c_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_c_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_c_axsize_reg
    ,output reg [31:0] wr_req_desc_c_attr_reg
    ,output reg [31:0] wr_req_desc_c_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_c_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_c_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_c_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_c_axid_0_reg
    ,output reg [31:0] wr_req_desc_c_axid_1_reg
    ,output reg [31:0] wr_req_desc_c_axid_2_reg
    ,output reg [31:0] wr_req_desc_c_axid_3_reg
    ,output reg [31:0] wr_req_desc_c_axuser_0_reg
    ,output reg [31:0] wr_req_desc_c_axuser_1_reg
    ,output reg [31:0] wr_req_desc_c_axuser_2_reg
    ,output reg [31:0] wr_req_desc_c_axuser_3_reg
    ,output reg [31:0] wr_req_desc_c_axuser_4_reg
    ,output reg [31:0] wr_req_desc_c_axuser_5_reg
    ,output reg [31:0] wr_req_desc_c_axuser_6_reg
    ,output reg [31:0] wr_req_desc_c_axuser_7_reg
    ,output reg [31:0] wr_req_desc_c_axuser_8_reg
    ,output reg [31:0] wr_req_desc_c_axuser_9_reg
    ,output reg [31:0] wr_req_desc_c_axuser_10_reg
    ,output reg [31:0] wr_req_desc_c_axuser_11_reg
    ,output reg [31:0] wr_req_desc_c_axuser_12_reg
    ,output reg [31:0] wr_req_desc_c_axuser_13_reg
    ,output reg [31:0] wr_req_desc_c_axuser_14_reg
    ,output reg [31:0] wr_req_desc_c_axuser_15_reg
    ,output reg [31:0] wr_req_desc_c_wuser_0_reg
    ,output reg [31:0] wr_req_desc_c_wuser_1_reg
    ,output reg [31:0] wr_req_desc_c_wuser_2_reg
    ,output reg [31:0] wr_req_desc_c_wuser_3_reg
    ,output reg [31:0] wr_req_desc_c_wuser_4_reg
    ,output reg [31:0] wr_req_desc_c_wuser_5_reg
    ,output reg [31:0] wr_req_desc_c_wuser_6_reg
    ,output reg [31:0] wr_req_desc_c_wuser_7_reg
    ,output reg [31:0] wr_req_desc_c_wuser_8_reg
    ,output reg [31:0] wr_req_desc_c_wuser_9_reg
    ,output reg [31:0] wr_req_desc_c_wuser_10_reg
    ,output reg [31:0] wr_req_desc_c_wuser_11_reg
    ,output reg [31:0] wr_req_desc_c_wuser_12_reg
    ,output reg [31:0] wr_req_desc_c_wuser_13_reg
    ,output reg [31:0] wr_req_desc_c_wuser_14_reg
    ,output reg [31:0] wr_req_desc_c_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_c_resp_reg
    ,output reg [31:0] wr_resp_desc_c_xid_0_reg
    ,output reg [31:0] wr_resp_desc_c_xid_1_reg
    ,output reg [31:0] wr_resp_desc_c_xid_2_reg
    ,output reg [31:0] wr_resp_desc_c_xid_3_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_c_xuser_15_reg
    ,output reg [31:0] sn_req_desc_c_attr_reg
    ,output reg [31:0] sn_req_desc_c_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_c_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_c_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_c_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_c_resp_reg
    ,output reg [31:0] rd_req_desc_d_txn_type_reg
    ,output reg [31:0] rd_req_desc_d_size_reg
    ,output reg [31:0] rd_req_desc_d_axsize_reg
    ,output reg [31:0] rd_req_desc_d_attr_reg
    ,output reg [31:0] rd_req_desc_d_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_d_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_d_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_d_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_d_axid_0_reg
    ,output reg [31:0] rd_req_desc_d_axid_1_reg
    ,output reg [31:0] rd_req_desc_d_axid_2_reg
    ,output reg [31:0] rd_req_desc_d_axid_3_reg
    ,output reg [31:0] rd_req_desc_d_axuser_0_reg
    ,output reg [31:0] rd_req_desc_d_axuser_1_reg
    ,output reg [31:0] rd_req_desc_d_axuser_2_reg
    ,output reg [31:0] rd_req_desc_d_axuser_3_reg
    ,output reg [31:0] rd_req_desc_d_axuser_4_reg
    ,output reg [31:0] rd_req_desc_d_axuser_5_reg
    ,output reg [31:0] rd_req_desc_d_axuser_6_reg
    ,output reg [31:0] rd_req_desc_d_axuser_7_reg
    ,output reg [31:0] rd_req_desc_d_axuser_8_reg
    ,output reg [31:0] rd_req_desc_d_axuser_9_reg
    ,output reg [31:0] rd_req_desc_d_axuser_10_reg
    ,output reg [31:0] rd_req_desc_d_axuser_11_reg
    ,output reg [31:0] rd_req_desc_d_axuser_12_reg
    ,output reg [31:0] rd_req_desc_d_axuser_13_reg
    ,output reg [31:0] rd_req_desc_d_axuser_14_reg
    ,output reg [31:0] rd_req_desc_d_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_d_data_offset_reg
    ,output reg [31:0] rd_resp_desc_d_data_size_reg
    ,output reg [31:0] rd_resp_desc_d_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_d_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_d_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_d_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_d_resp_reg
    ,output reg [31:0] rd_resp_desc_d_xid_0_reg
    ,output reg [31:0] rd_resp_desc_d_xid_1_reg
    ,output reg [31:0] rd_resp_desc_d_xid_2_reg
    ,output reg [31:0] rd_resp_desc_d_xid_3_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_d_xuser_15_reg
    ,output reg [31:0] wr_req_desc_d_txn_type_reg
    ,output reg [31:0] wr_req_desc_d_size_reg
    ,output reg [31:0] wr_req_desc_d_data_offset_reg
    ,output reg [31:0] wr_req_desc_d_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_d_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_d_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_d_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_d_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_d_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_d_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_d_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_d_axsize_reg
    ,output reg [31:0] wr_req_desc_d_attr_reg
    ,output reg [31:0] wr_req_desc_d_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_d_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_d_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_d_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_d_axid_0_reg
    ,output reg [31:0] wr_req_desc_d_axid_1_reg
    ,output reg [31:0] wr_req_desc_d_axid_2_reg
    ,output reg [31:0] wr_req_desc_d_axid_3_reg
    ,output reg [31:0] wr_req_desc_d_axuser_0_reg
    ,output reg [31:0] wr_req_desc_d_axuser_1_reg
    ,output reg [31:0] wr_req_desc_d_axuser_2_reg
    ,output reg [31:0] wr_req_desc_d_axuser_3_reg
    ,output reg [31:0] wr_req_desc_d_axuser_4_reg
    ,output reg [31:0] wr_req_desc_d_axuser_5_reg
    ,output reg [31:0] wr_req_desc_d_axuser_6_reg
    ,output reg [31:0] wr_req_desc_d_axuser_7_reg
    ,output reg [31:0] wr_req_desc_d_axuser_8_reg
    ,output reg [31:0] wr_req_desc_d_axuser_9_reg
    ,output reg [31:0] wr_req_desc_d_axuser_10_reg
    ,output reg [31:0] wr_req_desc_d_axuser_11_reg
    ,output reg [31:0] wr_req_desc_d_axuser_12_reg
    ,output reg [31:0] wr_req_desc_d_axuser_13_reg
    ,output reg [31:0] wr_req_desc_d_axuser_14_reg
    ,output reg [31:0] wr_req_desc_d_axuser_15_reg
    ,output reg [31:0] wr_req_desc_d_wuser_0_reg
    ,output reg [31:0] wr_req_desc_d_wuser_1_reg
    ,output reg [31:0] wr_req_desc_d_wuser_2_reg
    ,output reg [31:0] wr_req_desc_d_wuser_3_reg
    ,output reg [31:0] wr_req_desc_d_wuser_4_reg
    ,output reg [31:0] wr_req_desc_d_wuser_5_reg
    ,output reg [31:0] wr_req_desc_d_wuser_6_reg
    ,output reg [31:0] wr_req_desc_d_wuser_7_reg
    ,output reg [31:0] wr_req_desc_d_wuser_8_reg
    ,output reg [31:0] wr_req_desc_d_wuser_9_reg
    ,output reg [31:0] wr_req_desc_d_wuser_10_reg
    ,output reg [31:0] wr_req_desc_d_wuser_11_reg
    ,output reg [31:0] wr_req_desc_d_wuser_12_reg
    ,output reg [31:0] wr_req_desc_d_wuser_13_reg
    ,output reg [31:0] wr_req_desc_d_wuser_14_reg
    ,output reg [31:0] wr_req_desc_d_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_d_resp_reg
    ,output reg [31:0] wr_resp_desc_d_xid_0_reg
    ,output reg [31:0] wr_resp_desc_d_xid_1_reg
    ,output reg [31:0] wr_resp_desc_d_xid_2_reg
    ,output reg [31:0] wr_resp_desc_d_xid_3_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_d_xuser_15_reg
    ,output reg [31:0] sn_req_desc_d_attr_reg
    ,output reg [31:0] sn_req_desc_d_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_d_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_d_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_d_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_d_resp_reg
    ,output reg [31:0] rd_req_desc_e_txn_type_reg
    ,output reg [31:0] rd_req_desc_e_size_reg
    ,output reg [31:0] rd_req_desc_e_axsize_reg
    ,output reg [31:0] rd_req_desc_e_attr_reg
    ,output reg [31:0] rd_req_desc_e_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_e_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_e_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_e_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_e_axid_0_reg
    ,output reg [31:0] rd_req_desc_e_axid_1_reg
    ,output reg [31:0] rd_req_desc_e_axid_2_reg
    ,output reg [31:0] rd_req_desc_e_axid_3_reg
    ,output reg [31:0] rd_req_desc_e_axuser_0_reg
    ,output reg [31:0] rd_req_desc_e_axuser_1_reg
    ,output reg [31:0] rd_req_desc_e_axuser_2_reg
    ,output reg [31:0] rd_req_desc_e_axuser_3_reg
    ,output reg [31:0] rd_req_desc_e_axuser_4_reg
    ,output reg [31:0] rd_req_desc_e_axuser_5_reg
    ,output reg [31:0] rd_req_desc_e_axuser_6_reg
    ,output reg [31:0] rd_req_desc_e_axuser_7_reg
    ,output reg [31:0] rd_req_desc_e_axuser_8_reg
    ,output reg [31:0] rd_req_desc_e_axuser_9_reg
    ,output reg [31:0] rd_req_desc_e_axuser_10_reg
    ,output reg [31:0] rd_req_desc_e_axuser_11_reg
    ,output reg [31:0] rd_req_desc_e_axuser_12_reg
    ,output reg [31:0] rd_req_desc_e_axuser_13_reg
    ,output reg [31:0] rd_req_desc_e_axuser_14_reg
    ,output reg [31:0] rd_req_desc_e_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_e_data_offset_reg
    ,output reg [31:0] rd_resp_desc_e_data_size_reg
    ,output reg [31:0] rd_resp_desc_e_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_e_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_e_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_e_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_e_resp_reg
    ,output reg [31:0] rd_resp_desc_e_xid_0_reg
    ,output reg [31:0] rd_resp_desc_e_xid_1_reg
    ,output reg [31:0] rd_resp_desc_e_xid_2_reg
    ,output reg [31:0] rd_resp_desc_e_xid_3_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_e_xuser_15_reg
    ,output reg [31:0] wr_req_desc_e_txn_type_reg
    ,output reg [31:0] wr_req_desc_e_size_reg
    ,output reg [31:0] wr_req_desc_e_data_offset_reg
    ,output reg [31:0] wr_req_desc_e_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_e_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_e_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_e_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_e_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_e_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_e_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_e_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_e_axsize_reg
    ,output reg [31:0] wr_req_desc_e_attr_reg
    ,output reg [31:0] wr_req_desc_e_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_e_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_e_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_e_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_e_axid_0_reg
    ,output reg [31:0] wr_req_desc_e_axid_1_reg
    ,output reg [31:0] wr_req_desc_e_axid_2_reg
    ,output reg [31:0] wr_req_desc_e_axid_3_reg
    ,output reg [31:0] wr_req_desc_e_axuser_0_reg
    ,output reg [31:0] wr_req_desc_e_axuser_1_reg
    ,output reg [31:0] wr_req_desc_e_axuser_2_reg
    ,output reg [31:0] wr_req_desc_e_axuser_3_reg
    ,output reg [31:0] wr_req_desc_e_axuser_4_reg
    ,output reg [31:0] wr_req_desc_e_axuser_5_reg
    ,output reg [31:0] wr_req_desc_e_axuser_6_reg
    ,output reg [31:0] wr_req_desc_e_axuser_7_reg
    ,output reg [31:0] wr_req_desc_e_axuser_8_reg
    ,output reg [31:0] wr_req_desc_e_axuser_9_reg
    ,output reg [31:0] wr_req_desc_e_axuser_10_reg
    ,output reg [31:0] wr_req_desc_e_axuser_11_reg
    ,output reg [31:0] wr_req_desc_e_axuser_12_reg
    ,output reg [31:0] wr_req_desc_e_axuser_13_reg
    ,output reg [31:0] wr_req_desc_e_axuser_14_reg
    ,output reg [31:0] wr_req_desc_e_axuser_15_reg
    ,output reg [31:0] wr_req_desc_e_wuser_0_reg
    ,output reg [31:0] wr_req_desc_e_wuser_1_reg
    ,output reg [31:0] wr_req_desc_e_wuser_2_reg
    ,output reg [31:0] wr_req_desc_e_wuser_3_reg
    ,output reg [31:0] wr_req_desc_e_wuser_4_reg
    ,output reg [31:0] wr_req_desc_e_wuser_5_reg
    ,output reg [31:0] wr_req_desc_e_wuser_6_reg
    ,output reg [31:0] wr_req_desc_e_wuser_7_reg
    ,output reg [31:0] wr_req_desc_e_wuser_8_reg
    ,output reg [31:0] wr_req_desc_e_wuser_9_reg
    ,output reg [31:0] wr_req_desc_e_wuser_10_reg
    ,output reg [31:0] wr_req_desc_e_wuser_11_reg
    ,output reg [31:0] wr_req_desc_e_wuser_12_reg
    ,output reg [31:0] wr_req_desc_e_wuser_13_reg
    ,output reg [31:0] wr_req_desc_e_wuser_14_reg
    ,output reg [31:0] wr_req_desc_e_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_e_resp_reg
    ,output reg [31:0] wr_resp_desc_e_xid_0_reg
    ,output reg [31:0] wr_resp_desc_e_xid_1_reg
    ,output reg [31:0] wr_resp_desc_e_xid_2_reg
    ,output reg [31:0] wr_resp_desc_e_xid_3_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_e_xuser_15_reg
    ,output reg [31:0] sn_req_desc_e_attr_reg
    ,output reg [31:0] sn_req_desc_e_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_e_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_e_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_e_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_e_resp_reg
    ,output reg [31:0] rd_req_desc_f_txn_type_reg
    ,output reg [31:0] rd_req_desc_f_size_reg
    ,output reg [31:0] rd_req_desc_f_axsize_reg
    ,output reg [31:0] rd_req_desc_f_attr_reg
    ,output reg [31:0] rd_req_desc_f_axaddr_0_reg
    ,output reg [31:0] rd_req_desc_f_axaddr_1_reg
    ,output reg [31:0] rd_req_desc_f_axaddr_2_reg
    ,output reg [31:0] rd_req_desc_f_axaddr_3_reg
    ,output reg [31:0] rd_req_desc_f_axid_0_reg
    ,output reg [31:0] rd_req_desc_f_axid_1_reg
    ,output reg [31:0] rd_req_desc_f_axid_2_reg
    ,output reg [31:0] rd_req_desc_f_axid_3_reg
    ,output reg [31:0] rd_req_desc_f_axuser_0_reg
    ,output reg [31:0] rd_req_desc_f_axuser_1_reg
    ,output reg [31:0] rd_req_desc_f_axuser_2_reg
    ,output reg [31:0] rd_req_desc_f_axuser_3_reg
    ,output reg [31:0] rd_req_desc_f_axuser_4_reg
    ,output reg [31:0] rd_req_desc_f_axuser_5_reg
    ,output reg [31:0] rd_req_desc_f_axuser_6_reg
    ,output reg [31:0] rd_req_desc_f_axuser_7_reg
    ,output reg [31:0] rd_req_desc_f_axuser_8_reg
    ,output reg [31:0] rd_req_desc_f_axuser_9_reg
    ,output reg [31:0] rd_req_desc_f_axuser_10_reg
    ,output reg [31:0] rd_req_desc_f_axuser_11_reg
    ,output reg [31:0] rd_req_desc_f_axuser_12_reg
    ,output reg [31:0] rd_req_desc_f_axuser_13_reg
    ,output reg [31:0] rd_req_desc_f_axuser_14_reg
    ,output reg [31:0] rd_req_desc_f_axuser_15_reg
    ,output reg [31:0] rd_resp_desc_f_data_offset_reg
    ,output reg [31:0] rd_resp_desc_f_data_size_reg
    ,output reg [31:0] rd_resp_desc_f_data_host_addr_0_reg
    ,output reg [31:0] rd_resp_desc_f_data_host_addr_1_reg
    ,output reg [31:0] rd_resp_desc_f_data_host_addr_2_reg
    ,output reg [31:0] rd_resp_desc_f_data_host_addr_3_reg
    ,output reg [31:0] rd_resp_desc_f_resp_reg
    ,output reg [31:0] rd_resp_desc_f_xid_0_reg
    ,output reg [31:0] rd_resp_desc_f_xid_1_reg
    ,output reg [31:0] rd_resp_desc_f_xid_2_reg
    ,output reg [31:0] rd_resp_desc_f_xid_3_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_0_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_1_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_2_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_3_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_4_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_5_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_6_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_7_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_8_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_9_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_10_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_11_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_12_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_13_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_14_reg
    ,output reg [31:0] rd_resp_desc_f_xuser_15_reg
    ,output reg [31:0] wr_req_desc_f_txn_type_reg
    ,output reg [31:0] wr_req_desc_f_size_reg
    ,output reg [31:0] wr_req_desc_f_data_offset_reg
    ,output reg [31:0] wr_req_desc_f_data_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_f_data_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_f_data_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_f_data_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_f_wstrb_host_addr_0_reg
    ,output reg [31:0] wr_req_desc_f_wstrb_host_addr_1_reg
    ,output reg [31:0] wr_req_desc_f_wstrb_host_addr_2_reg
    ,output reg [31:0] wr_req_desc_f_wstrb_host_addr_3_reg
    ,output reg [31:0] wr_req_desc_f_axsize_reg
    ,output reg [31:0] wr_req_desc_f_attr_reg
    ,output reg [31:0] wr_req_desc_f_axaddr_0_reg
    ,output reg [31:0] wr_req_desc_f_axaddr_1_reg
    ,output reg [31:0] wr_req_desc_f_axaddr_2_reg
    ,output reg [31:0] wr_req_desc_f_axaddr_3_reg
    ,output reg [31:0] wr_req_desc_f_axid_0_reg
    ,output reg [31:0] wr_req_desc_f_axid_1_reg
    ,output reg [31:0] wr_req_desc_f_axid_2_reg
    ,output reg [31:0] wr_req_desc_f_axid_3_reg
    ,output reg [31:0] wr_req_desc_f_axuser_0_reg
    ,output reg [31:0] wr_req_desc_f_axuser_1_reg
    ,output reg [31:0] wr_req_desc_f_axuser_2_reg
    ,output reg [31:0] wr_req_desc_f_axuser_3_reg
    ,output reg [31:0] wr_req_desc_f_axuser_4_reg
    ,output reg [31:0] wr_req_desc_f_axuser_5_reg
    ,output reg [31:0] wr_req_desc_f_axuser_6_reg
    ,output reg [31:0] wr_req_desc_f_axuser_7_reg
    ,output reg [31:0] wr_req_desc_f_axuser_8_reg
    ,output reg [31:0] wr_req_desc_f_axuser_9_reg
    ,output reg [31:0] wr_req_desc_f_axuser_10_reg
    ,output reg [31:0] wr_req_desc_f_axuser_11_reg
    ,output reg [31:0] wr_req_desc_f_axuser_12_reg
    ,output reg [31:0] wr_req_desc_f_axuser_13_reg
    ,output reg [31:0] wr_req_desc_f_axuser_14_reg
    ,output reg [31:0] wr_req_desc_f_axuser_15_reg
    ,output reg [31:0] wr_req_desc_f_wuser_0_reg
    ,output reg [31:0] wr_req_desc_f_wuser_1_reg
    ,output reg [31:0] wr_req_desc_f_wuser_2_reg
    ,output reg [31:0] wr_req_desc_f_wuser_3_reg
    ,output reg [31:0] wr_req_desc_f_wuser_4_reg
    ,output reg [31:0] wr_req_desc_f_wuser_5_reg
    ,output reg [31:0] wr_req_desc_f_wuser_6_reg
    ,output reg [31:0] wr_req_desc_f_wuser_7_reg
    ,output reg [31:0] wr_req_desc_f_wuser_8_reg
    ,output reg [31:0] wr_req_desc_f_wuser_9_reg
    ,output reg [31:0] wr_req_desc_f_wuser_10_reg
    ,output reg [31:0] wr_req_desc_f_wuser_11_reg
    ,output reg [31:0] wr_req_desc_f_wuser_12_reg
    ,output reg [31:0] wr_req_desc_f_wuser_13_reg
    ,output reg [31:0] wr_req_desc_f_wuser_14_reg
    ,output reg [31:0] wr_req_desc_f_wuser_15_reg
    ,output reg [31:0] wr_resp_desc_f_resp_reg
    ,output reg [31:0] wr_resp_desc_f_xid_0_reg
    ,output reg [31:0] wr_resp_desc_f_xid_1_reg
    ,output reg [31:0] wr_resp_desc_f_xid_2_reg
    ,output reg [31:0] wr_resp_desc_f_xid_3_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_0_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_1_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_2_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_3_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_4_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_5_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_6_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_7_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_8_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_9_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_10_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_11_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_12_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_13_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_14_reg
    ,output reg [31:0] wr_resp_desc_f_xuser_15_reg
    ,output reg [31:0] sn_req_desc_f_attr_reg
    ,output reg [31:0] sn_req_desc_f_acaddr_0_reg
    ,output reg [31:0] sn_req_desc_f_acaddr_1_reg
    ,output reg [31:0] sn_req_desc_f_acaddr_2_reg
    ,output reg [31:0] sn_req_desc_f_acaddr_3_reg
    ,output reg [31:0] sn_resp_desc_f_resp_reg
    
    ,input [31:0] uc2rb_intr_error_status_reg
    ,input [31:0] uc2rb_rd_req_fifo_pop_desc_reg
    ,input [31:0] uc2rb_rd_req_fifo_fill_level_reg
    ,input [31:0] uc2rb_rd_resp_fifo_free_level_reg
    ,input [31:0] uc2rb_rd_resp_intr_comp_status_reg
    ,input [31:0] uc2rb_wr_req_fifo_pop_desc_reg
    ,input [31:0] uc2rb_wr_req_fifo_fill_level_reg
    ,input [31:0] uc2rb_wr_resp_fifo_free_level_reg
    ,input [31:0] uc2rb_wr_resp_intr_comp_status_reg
    ,input [31:0] uc2rb_sn_req_fifo_free_level_reg
    ,input [31:0] uc2rb_sn_req_intr_comp_status_reg
    ,input [31:0] uc2rb_sn_resp_fifo_pop_desc_reg
    ,input [31:0] uc2rb_sn_resp_fifo_fill_level_reg
    ,input [31:0] uc2rb_sn_data_fifo_pop_desc_reg
    ,input [31:0] uc2rb_sn_data_fifo_fill_level_reg
    ,input [31:0] uc2rb_rd_req_desc_0_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_0_size_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_0_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_0_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_0_size_reg
    ,input [31:0] uc2rb_wr_req_desc_0_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_0_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_0_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_1_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_1_size_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_1_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_1_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_1_size_reg
    ,input [31:0] uc2rb_wr_req_desc_1_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_1_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_1_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_2_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_2_size_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_2_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_2_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_2_size_reg
    ,input [31:0] uc2rb_wr_req_desc_2_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_2_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_2_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_3_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_3_size_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_3_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_3_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_3_size_reg
    ,input [31:0] uc2rb_wr_req_desc_3_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_3_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_3_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_4_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_4_size_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_4_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_4_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_4_size_reg
    ,input [31:0] uc2rb_wr_req_desc_4_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_4_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_4_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_5_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_5_size_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_5_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_5_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_5_size_reg
    ,input [31:0] uc2rb_wr_req_desc_5_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_5_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_5_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_6_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_6_size_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_6_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_6_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_6_size_reg
    ,input [31:0] uc2rb_wr_req_desc_6_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_6_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_6_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_7_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_7_size_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_7_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_7_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_7_size_reg
    ,input [31:0] uc2rb_wr_req_desc_7_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_7_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_7_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_8_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_8_size_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_8_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_8_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_8_size_reg
    ,input [31:0] uc2rb_wr_req_desc_8_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_8_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_8_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_9_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_9_size_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_9_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_9_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_9_size_reg
    ,input [31:0] uc2rb_wr_req_desc_9_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_9_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_9_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_a_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_a_size_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_a_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_a_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_a_size_reg
    ,input [31:0] uc2rb_wr_req_desc_a_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_a_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_a_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_b_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_b_size_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_b_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_b_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_b_size_reg
    ,input [31:0] uc2rb_wr_req_desc_b_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_b_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_b_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_c_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_c_size_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_c_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_c_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_c_size_reg
    ,input [31:0] uc2rb_wr_req_desc_c_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_c_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_c_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_d_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_d_size_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_d_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_d_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_d_size_reg
    ,input [31:0] uc2rb_wr_req_desc_d_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_d_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_d_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_e_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_e_size_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_e_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_e_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_e_size_reg
    ,input [31:0] uc2rb_wr_req_desc_e_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_e_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_e_resp_reg
    ,input [31:0] uc2rb_rd_req_desc_f_txn_type_reg
    ,input [31:0] uc2rb_rd_req_desc_f_size_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axsize_reg
    ,input [31:0] uc2rb_rd_req_desc_f_attr_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_0_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_1_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_2_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_3_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axid_0_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axid_1_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axid_2_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axid_3_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_0_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_1_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_2_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_3_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_4_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_5_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_6_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_7_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_8_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_9_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_10_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_11_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_12_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_13_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_14_reg
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_f_txn_type_reg
    ,input [31:0] uc2rb_wr_req_desc_f_size_reg
    ,input [31:0] uc2rb_wr_req_desc_f_data_offset_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axsize_reg
    ,input [31:0] uc2rb_wr_req_desc_f_attr_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_0_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_1_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_2_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_3_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axid_0_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axid_1_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axid_2_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axid_3_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_15_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_0_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_1_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_2_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_3_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_4_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_5_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_6_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_7_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_8_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_9_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_10_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_11_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_12_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_13_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_14_reg
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_15_reg
    ,input [31:0] uc2rb_sn_resp_desc_f_resp_reg
    
    ,input [31:0] uc2rb_intr_error_status_reg_we
    ,input [31:0] uc2rb_rd_req_fifo_pop_desc_reg_we
    ,input [31:0] uc2rb_rd_req_fifo_fill_level_reg_we
    ,input [31:0] uc2rb_rd_resp_fifo_free_level_reg_we
    ,input [31:0] uc2rb_rd_resp_intr_comp_status_reg_we
    ,input [31:0] uc2rb_wr_req_fifo_pop_desc_reg_we
    ,input [31:0] uc2rb_wr_req_fifo_fill_level_reg_we
    ,input [31:0] uc2rb_wr_resp_fifo_free_level_reg_we
    ,input [31:0] uc2rb_wr_resp_intr_comp_status_reg_we
    ,input [31:0] uc2rb_sn_req_fifo_free_level_reg_we
    ,input [31:0] uc2rb_sn_req_intr_comp_status_reg_we
    ,input [31:0] uc2rb_sn_resp_fifo_pop_desc_reg_we
    ,input [31:0] uc2rb_sn_resp_fifo_fill_level_reg_we
    ,input [31:0] uc2rb_sn_data_fifo_pop_desc_reg_we
    ,input [31:0] uc2rb_sn_data_fifo_fill_level_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_0_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_0_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_0_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_1_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_1_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_1_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_2_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_2_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_2_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_3_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_3_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_3_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_4_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_4_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_4_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_5_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_5_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_5_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_6_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_6_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_6_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_7_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_7_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_7_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_8_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_8_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_8_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_9_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_9_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_9_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_a_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_a_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_a_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_b_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_b_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_b_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_c_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_c_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_c_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_d_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_d_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_d_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_e_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_e_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_e_resp_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_txn_type_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_size_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axsize_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_attr_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axaddr_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axid_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axid_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axid_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axid_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_0_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_1_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_2_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_3_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_4_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_5_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_6_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_7_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_8_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_9_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_10_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_11_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_12_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_13_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_14_reg_we
    ,input [31:0] uc2rb_rd_req_desc_f_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_txn_type_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_size_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_data_offset_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axsize_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_attr_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axaddr_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axid_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axid_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axid_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axid_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_axuser_15_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_0_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_1_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_2_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_3_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_4_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_5_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_6_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_7_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_8_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_9_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_10_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_11_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_12_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_13_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_14_reg_we
    ,input [31:0] uc2rb_wr_req_desc_f_wuser_15_reg_we
    ,input [31:0] uc2rb_sn_resp_desc_f_resp_reg_we
    
    
    // register interface between hm-rb
    ,input [31:0] hm2rb_intr_error_status_reg 
    ,input [31:0] hm2rb_intr_error_status_reg_we 
    
    // register interface between IH-rb
    
    ,input [31:0] ih2rb_c2h_intr_status_0_reg 
    ,input [31:0] ih2rb_c2h_intr_status_1_reg
    ,input [31:0] ih2rb_intr_c2h_toggle_status_0_reg 
    ,input [31:0] ih2rb_intr_c2h_toggle_status_1_reg 
    ,input [31:0] ih2rb_c2h_gpio_0_reg
    ,input [31:0] ih2rb_c2h_gpio_1_reg
    ,input [31:0] ih2rb_c2h_gpio_2_reg
    ,input [31:0] ih2rb_c2h_gpio_3_reg
    ,input [31:0] ih2rb_c2h_gpio_4_reg
    ,input [31:0] ih2rb_c2h_gpio_5_reg
    ,input [31:0] ih2rb_c2h_gpio_6_reg
    ,input [31:0] ih2rb_c2h_gpio_7_reg
    
    ,input [31:0] ih2rb_c2h_gpio_0_reg_we
    ,input [31:0] ih2rb_c2h_gpio_1_reg_we
    ,input [31:0] ih2rb_c2h_gpio_2_reg_we
    ,input [31:0] ih2rb_c2h_gpio_3_reg_we
    ,input [31:0] ih2rb_c2h_gpio_4_reg_we
    ,input [31:0] ih2rb_c2h_gpio_5_reg_we
    ,input [31:0] ih2rb_c2h_gpio_6_reg_we
    ,input [31:0] ih2rb_c2h_gpio_7_reg_we
    
    
    ,input [31:0] ih2rb_c2h_intr_status_0_reg_we 
    ,input [31:0] ih2rb_c2h_intr_status_1_reg_we
    ,input [31:0] ih2rb_intr_c2h_toggle_status_0_reg_we 
    ,input [31:0] ih2rb_intr_c2h_toggle_status_1_reg_we 

    );
   


   localparam S_ACE_USR_DATA_WIDTH = S_ACE_USR_XX_DATA_WIDTH;

   // BRIDGE_TYPE DEFINITION
   //0x0 : AXI3 Bridge in Master Mode
   //0x1 : AXI3 Bridge in Slave Mode
   //0x2 : AXI4 Bridge in Master Mode
   //0x3 : AXI4 Bridge in Slave Mode
   //0x4 : AXI4-lite Bridge in Master Mode
   //0x5 : AXI4-lite Bridge in Slave Mode
   //0x6 : Reserved
   //0x7 : Reserved
   //0x8 : ACE Bridge in Master Mode
   //0x9 : ACE Bridge in Slave Mode

   localparam BRIDGE_MSB = ((`CLOG2(XX_RAM_SIZE*8)) - 1 );
   localparam [0:0] LAST_BRIDGE_DECODE = LAST_BRIDGE;
   localparam [31:0] DWIDTH_DECODE = (S_ACE_USR_DATA_WIDTH==128)?3'h4:(S_ACE_USR_DATA_WIDTH==64)?3'h3:(S_ACE_USR_DATA_WIDTH==32)?3'h2:3'h4;
   localparam [31:0] IDWIDTH_DECODE = S_ACE_USR_ID_WIDTH;
   localparam [31:0] EXTEND_WSTRB_DECODE = EXTEND_WSTRB;
   localparam [31:0] ARUSER_WIDTH_DECODE = S_ACE_USR_ARUSER_WIDTH;        
   localparam [31:0] RUSER_WIDTH_DECODE  = S_ACE_USR_RUSER_WIDTH;         
   localparam [31:0] AWUSER_WIDTH_DECODE = S_ACE_USR_AWUSER_WIDTH;        
   localparam [31:0] WUSER_WIDTH_DECODE  = S_ACE_USR_WUSER_WIDTH;         
   localparam [31:0] BUSER_WIDTH_DECODE  = S_ACE_USR_BUSER_WIDTH;         
   localparam [31:0] XX_MAX_DESC_DECODE = XX_MAX_DESC;
   localparam [31:0] SN_MAX_DESC_DECODE = SN_MAX_DESC;

   

   localparam [31:0] BRIDGE_IDENTIFICATION_REG = 32'hC3A89FE1;
   localparam [31:0] LAST_BRIDGE_REG = { 31'h0, LAST_BRIDGE_DECODE[0] };
   localparam [31:0] VERSION_REG = 32'h0100;
   localparam [31:0] BRIDGE_TYPE_REG = 32'h0009;
   localparam [31:0] BRIDGE_CONFIG_REG = {19'b0,EXTEND_WSTRB_DECODE[0], IDWIDTH_DECODE[7:0],1'b0,DWIDTH_DECODE[2:0]};
   localparam [31:0] BRIDGE_RD_USER_CONFIG_REG = {  12'b0
                                                    , RUSER_WIDTH_DECODE[9:0]
                                                    , ARUSER_WIDTH_DECODE[9:0]
                                                    };
   localparam [31:0] BRIDGE_WR_USER_CONFIG_REG = {  2'b0
                                                    , BUSER_WIDTH_DECODE[9:0]
                                                    , WUSER_WIDTH_DECODE[9:0]
                                                    , AWUSER_WIDTH_DECODE[9:0]
                                                    };
   localparam [31:0] RD_MAX_DESC_REG = {16'h0, XX_MAX_DESC_DECODE[7:0], XX_MAX_DESC_DECODE[7:0]};
   localparam [31:0] WR_MAX_DESC_REG = {16'h0, XX_MAX_DESC_DECODE[7:0], XX_MAX_DESC_DECODE[7:0]};
   localparam [31:0] SN_MAX_DESC_REG = {8'h0, SN_MAX_DESC_DECODE[7:0], SN_MAX_DESC_DECODE[7:0], SN_MAX_DESC_DECODE[7:0]};
   
   
   reg [31:0] intr_error_clear_reg_clear;
   reg [31:0] intr_c2h_toggle_clear_0_reg_clear ;
   reg [31:0] intr_c2h_toggle_clear_1_reg_clear ;


   reg [31:0] rd_req_free_desc_reg_clear;
   reg [31:0] rd_resp_fifo_push_desc_reg_clear;
   reg [31:0] rd_resp_intr_comp_clear_reg_clear;
   reg [31:0] wr_req_free_desc_reg_clear;
   reg [31:0] wr_resp_fifo_push_desc_reg_clear;
   reg [31:0] wr_resp_intr_comp_clear_reg_clear;
   reg [31:0] sn_req_fifo_push_desc_reg_clear;
   reg [31:0] sn_req_intr_comp_clear_reg_clear;
   reg [31:0] sn_resp_free_desc_reg_clear;
   reg [31:0] sn_data_free_desc_reg_clear;



   reg 	      match_fifo_pop_desc; 
   reg [S_AXI_DATA_WIDTH-1:0] reg_data_out_pipeline; 
   
   reg [(`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8)))-1:0] wdata_ram_addr;
   reg 							       wdata_ram_rd_en;
   
   wire [S_ACE_USR_XX_DATA_WIDTH-1:0] 			       wdata_ram_data;                      
   wire [(S_ACE_USR_XX_DATA_WIDTH/8)-1:0] 		       wstrb_ram_data;
   
   reg 							       wdata_ram_data_ready;
   reg 							       wdata_ram_data_ready_1;

   reg 							       cddata_ram_data_ready;
   reg 							       cddata_ram_data_ready_1;
   reg 							       cddata_ram_data_ready_2; 
   
   wire [S_ACE_USR_SN_DATA_WIDTH-1:0] 			       cddata_ram_data;                         
   
   reg [(`CLOG2(SN_RAM_SIZE/(S_ACE_USR_SN_DATA_WIDTH/8)))-1:0] cddata_ram_addr;
   reg 							       cddata_ram_rd_en;
   
   reg [(`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8)))-1:0] wstrb_ram_addr;
   reg 							       wstrb_ram_rd_en;

   reg 							       rdata_ram_we;
   reg [(`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8)))-1:0] rdata_ram_addr;
   reg [S_ACE_USR_XX_DATA_WIDTH-1:0] 			       rdata_ram_data;
   reg [(S_ACE_USR_XX_DATA_WIDTH/8) -1:0] 		       rdata_ram_bwe;
   
   reg [(`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8)))-1:0] uc2rb_rd_addr_reg;



   // registering axi4lite signals
   reg [S_AXI_ADDR_WIDTH-1 : 0] 			       axi_awaddr;
   reg 							       axi_awready;
   reg 							       axi_wready;
   reg [1 : 0] 						       axi_bresp;
   reg 							       axi_bvalid;
   reg [S_AXI_ADDR_WIDTH-1 : 0] 			       axi_araddr;
   reg 							       axi_arready;
   reg [S_AXI_DATA_WIDTH-1 : 0] 			       axi_rdata;
   reg [1 : 0] 						       axi_rresp;
   reg 							       axi_rvalid;

   // example-specific design signals
   // local parameter for addressing 32 bit / 64 bit c_s_axi_data_width
   // addr_lsb is used for addressing 32/64 bit registers/memories
   // addr_lsb = 2 for 32 bits (n downto 2)
   // addr_lsb = 3 for 64 bits (n downto 3)
   localparam integer 					       addr_lsb = (S_AXI_DATA_WIDTH/32) + 1;
   localparam integer 					       opt_mem_addr_bits = 8;

   wire 						       reg_rd_en;
   wire 						       reg_wr_en;
   reg [S_AXI_DATA_WIDTH-1:0] 				       reg_data_out;



   reg 							       wdata_ram_data_ready_2; 
   reg 							       wstrb_ram_data_ready_2; 

   reg 							       wstrb_ram_data_ready;
   reg 							       wstrb_ram_data_ready_1;


   assign s_axi_awready    = axi_awready;
   assign s_axi_wready     = axi_wready;
   assign s_axi_bresp      = axi_bresp;
   assign s_axi_bvalid     = axi_bvalid;
   assign s_axi_arready    = axi_arready;
   assign s_axi_rdata      = axi_rdata;
   assign s_axi_rresp      = axi_rresp;
   assign s_axi_rvalid     = axi_rvalid;


 wire bnext;
   reg 	awready_state;

   localparam AWREADY_IDLE =0, WAIT_FOR_BNEXT = 1;
   
   
   //******************************************************************************/
   //AXI SLAVE STATE MACHINE
   //******************************************************************************/
   assign bnext = s_axi_bready & axi_bvalid;
      
   // implement axi_awready generation
   // axi_awready is asserted for one clk clock cycle when both
   // s_axi_awvalid and s_axi_wvalid are asserted. axi_awready is
   // de-asserted when reset is low.

   always @( posedge clk )
     begin
        if ( ~resetn  ) begin
           axi_awready <= 1'b0;
	   awready_state <= AWREADY_IDLE;
	end
        else
          begin
	     case(awready_state)
	       AWREADY_IDLE:
		 if (~axi_awready && s_axi_awvalid && s_axi_wvalid) begin
		    // slave is ready to accept write address when 
		    // there is a valid write address and write data
		    // on the write address and data bus. this design 
		    // expects no outstanding transactions. 
		    axi_awready <= 1'b1;
		    awready_state <= WAIT_FOR_BNEXT;
		 end
		 else begin
		    axi_awready <= 1'b0;
		    awready_state <= AWREADY_IDLE;
		 end // else: !if(~axi_awready && s_axi_awvalid && s_axi_wvalid)
	       WAIT_FOR_BNEXT:
		 if (bnext) begin
		    axi_awready <= 1'b0;
		    awready_state <= AWREADY_IDLE;
		 end
		 else begin
		    axi_awready <= 1'b0;
		    awready_state <= WAIT_FOR_BNEXT;
		 end
	       default:
		 awready_state <= awready_state;
	     endcase
	  end
     end // always @ ( posedge clk )
   

   // implement axi_awaddr latching
   // this process is used to latch the address when both 
   // s_axi_awvalid and s_axi_wvalid are valid. 

   always @( posedge clk )
     begin
        if ( ~resetn  )
          axi_awaddr <= 0;
        else
          begin    
             if (~axi_awready && s_axi_awvalid && s_axi_wvalid)
               // write address latching 
               axi_awaddr <= s_axi_awaddr;
          end 
     end       

   reg wready_state;

   localparam WREADY_IDLE=1,WREADY_ASSERTED=0;
   
   // implement axi_wready generation
   // axi_wready is asserted for one clk clock cycle when both
   // s_axi_awvalid and s_axi_wvalid are asserted. axi_wready is 
   // de-asserted when reset is low. 


   always @( posedge clk )
     begin
        if ( ~resetn  ) begin
           axi_wready <= 1'b0;
	   wready_state <= WREADY_IDLE;
	end
        else
          begin
	     case(wready_state)
	       WREADY_IDLE:
		 if (~axi_wready && s_axi_wvalid && s_axi_awvalid)
		   begin
		      // slave is ready to accept write data when 
		      // there is a valid write address and write data
		      // on the write address and data bus. this design 
		      // expects no outstanding transactions. 
		      axi_wready <= 1'b1;
		      wready_state <= WREADY_ASSERTED;
		   end
		 else begin
		    axi_wready <= 1'b0;
		    wready_state <= WREADY_IDLE;
		 end // else: !if(~axi_wready && s_axi_awvalid && s_axi_wvalid)
	       WREADY_ASSERTED:
		 if (bnext) begin
		    axi_wready <= 1'b0;
		    wready_state <= WREADY_IDLE;
		 end
		 else begin
		    axi_wready <= 1'b0;
		    wready_state <= WREADY_ASSERTED;
		 end
	       default:
		 wready_state <= wready_state;
	     endcase
	  end
     end // always @ ( posedge clk )

   // implement memory mapped register select and write logic generation
   // the write data is accepted and written to memory mapped registers when
   // axi_awready, s_axi_wvalid, axi_wready and s_axi_wvalid are asserted. write strobes are used to
   // select byte enables of slave registers while writing.
   // these registers are cleared when reset (active low) is applied.
   // slave register write enable is asserted when valid address and data are available
   // and the slave is ready to accept the write address and write data.
   assign reg_wr_en = axi_wready && s_axi_wvalid && axi_awready && s_axi_awvalid;   

   integer                                i;
   integer                                byte_index;

   always @( posedge clk )
     begin
        if ( ~resetn) 
          begin
             reset_reg                     <=32'hFFFFFFFF; 
          end
        else
          begin
             if ( reg_wr_en && (~|axi_awaddr[BRIDGE_MSB:6]) && (&axi_awaddr[5:2]) ) // Writing to RESET_REG
               begin
                  for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                    if ( s_axi_wstrb[byte_index] == 1 ) begin
                       reset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                    end  

               end
          end // else: !if( ~resetn)
     end // always @ ( posedge clk )
   
   
   //rw/rwso register write logic
   always @( posedge clk )
     begin
        if ( ~rst_n)
          begin
             
             mode_select_reg <= 32'h0;
             h2c_intr_0_reg <= 32'h0;
             h2c_intr_1_reg <= 32'h0;
             h2c_intr_2_reg <= 32'h0;
             h2c_intr_3_reg <= 32'h0;
             intr_c2h_toggle_clear_0_reg <= 32'h0;
             intr_c2h_toggle_enable_0_reg <= 32'h0;
             intr_c2h_toggle_clear_1_reg <= 32'h0;
             intr_c2h_toggle_enable_1_reg <= 32'h0;
             h2c_gpio_0_reg <= 32'h0;
             h2c_gpio_1_reg <= 32'h0;
             h2c_gpio_2_reg <= 32'h0;
             h2c_gpio_3_reg <= 32'h0;
             h2c_gpio_4_reg <= 32'h0;
             h2c_gpio_5_reg <= 32'h0;
             h2c_gpio_6_reg <= 32'h0;
             h2c_gpio_7_reg <= 32'h0;
             h2c_gpio_8_reg <= 32'h0;
             h2c_gpio_9_reg <= 32'h0;
             h2c_gpio_10_reg <= 32'h0;
             h2c_gpio_11_reg <= 32'h0;
             h2c_gpio_12_reg <= 32'h0;
             h2c_gpio_13_reg <= 32'h0;
             h2c_gpio_14_reg <= 32'h0;
             h2c_gpio_15_reg <= 32'h0;
             intr_error_clear_reg <= 32'h0;
             intr_error_enable_reg <= 32'h0;
             rd_req_free_desc_reg <= 32'h0;
             rd_resp_fifo_push_desc_reg <= 32'h0;
             rd_resp_intr_comp_clear_reg <= 32'h0;
             rd_resp_intr_comp_enable_reg <= 32'h0;
             wr_req_free_desc_reg <= 32'h0;
             wr_resp_fifo_push_desc_reg <= 32'h0;
             wr_resp_intr_comp_clear_reg <= 32'h0;
             wr_resp_intr_comp_enable_reg <= 32'h0;
             sn_req_fifo_push_desc_reg <= 32'h0;
             sn_req_intr_comp_clear_reg <= 32'h0;
             sn_req_intr_comp_enable_reg <= 32'h0;
             sn_resp_free_desc_reg <= 32'h0;
             sn_data_free_desc_reg <= 32'h0;
             intr_fifo_enable_reg <= 32'h0;
             rd_resp_desc_0_data_offset_reg <= 32'h0;
             rd_resp_desc_0_data_size_reg <= 32'h0;
             rd_resp_desc_0_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_0_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_0_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_0_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_0_resp_reg <= 32'h0;
             rd_resp_desc_0_xid_0_reg <= 32'h0;
             rd_resp_desc_0_xid_1_reg <= 32'h0;
             rd_resp_desc_0_xid_2_reg <= 32'h0;
             rd_resp_desc_0_xid_3_reg <= 32'h0;
             rd_resp_desc_0_xuser_0_reg <= 32'h0;
             rd_resp_desc_0_xuser_1_reg <= 32'h0;
             rd_resp_desc_0_xuser_2_reg <= 32'h0;
             rd_resp_desc_0_xuser_3_reg <= 32'h0;
             rd_resp_desc_0_xuser_4_reg <= 32'h0;
             rd_resp_desc_0_xuser_5_reg <= 32'h0;
             rd_resp_desc_0_xuser_6_reg <= 32'h0;
             rd_resp_desc_0_xuser_7_reg <= 32'h0;
             rd_resp_desc_0_xuser_8_reg <= 32'h0;
             rd_resp_desc_0_xuser_9_reg <= 32'h0;
             rd_resp_desc_0_xuser_10_reg <= 32'h0;
             rd_resp_desc_0_xuser_11_reg <= 32'h0;
             rd_resp_desc_0_xuser_12_reg <= 32'h0;
             rd_resp_desc_0_xuser_13_reg <= 32'h0;
             rd_resp_desc_0_xuser_14_reg <= 32'h0;
             rd_resp_desc_0_xuser_15_reg <= 32'h0;
             wr_req_desc_0_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_0_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_0_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_0_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_0_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_0_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_0_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_0_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_0_resp_reg <= 32'h0;
             wr_resp_desc_0_xid_0_reg <= 32'h0;
             wr_resp_desc_0_xid_1_reg <= 32'h0;
             wr_resp_desc_0_xid_2_reg <= 32'h0;
             wr_resp_desc_0_xid_3_reg <= 32'h0;
             wr_resp_desc_0_xuser_0_reg <= 32'h0;
             wr_resp_desc_0_xuser_1_reg <= 32'h0;
             wr_resp_desc_0_xuser_2_reg <= 32'h0;
             wr_resp_desc_0_xuser_3_reg <= 32'h0;
             wr_resp_desc_0_xuser_4_reg <= 32'h0;
             wr_resp_desc_0_xuser_5_reg <= 32'h0;
             wr_resp_desc_0_xuser_6_reg <= 32'h0;
             wr_resp_desc_0_xuser_7_reg <= 32'h0;
             wr_resp_desc_0_xuser_8_reg <= 32'h0;
             wr_resp_desc_0_xuser_9_reg <= 32'h0;
             wr_resp_desc_0_xuser_10_reg <= 32'h0;
             wr_resp_desc_0_xuser_11_reg <= 32'h0;
             wr_resp_desc_0_xuser_12_reg <= 32'h0;
             wr_resp_desc_0_xuser_13_reg <= 32'h0;
             wr_resp_desc_0_xuser_14_reg <= 32'h0;
             wr_resp_desc_0_xuser_15_reg <= 32'h0;
             sn_req_desc_0_attr_reg <= 32'h0;
             sn_req_desc_0_acaddr_0_reg <= 32'h0;
             sn_req_desc_0_acaddr_1_reg <= 32'h0;
             sn_req_desc_0_acaddr_2_reg <= 32'h0;
             sn_req_desc_0_acaddr_3_reg <= 32'h0;
             rd_resp_desc_1_data_offset_reg <= 32'h0;
             rd_resp_desc_1_data_size_reg <= 32'h0;
             rd_resp_desc_1_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_1_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_1_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_1_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_1_resp_reg <= 32'h0;
             rd_resp_desc_1_xid_0_reg <= 32'h0;
             rd_resp_desc_1_xid_1_reg <= 32'h0;
             rd_resp_desc_1_xid_2_reg <= 32'h0;
             rd_resp_desc_1_xid_3_reg <= 32'h0;
             rd_resp_desc_1_xuser_0_reg <= 32'h0;
             rd_resp_desc_1_xuser_1_reg <= 32'h0;
             rd_resp_desc_1_xuser_2_reg <= 32'h0;
             rd_resp_desc_1_xuser_3_reg <= 32'h0;
             rd_resp_desc_1_xuser_4_reg <= 32'h0;
             rd_resp_desc_1_xuser_5_reg <= 32'h0;
             rd_resp_desc_1_xuser_6_reg <= 32'h0;
             rd_resp_desc_1_xuser_7_reg <= 32'h0;
             rd_resp_desc_1_xuser_8_reg <= 32'h0;
             rd_resp_desc_1_xuser_9_reg <= 32'h0;
             rd_resp_desc_1_xuser_10_reg <= 32'h0;
             rd_resp_desc_1_xuser_11_reg <= 32'h0;
             rd_resp_desc_1_xuser_12_reg <= 32'h0;
             rd_resp_desc_1_xuser_13_reg <= 32'h0;
             rd_resp_desc_1_xuser_14_reg <= 32'h0;
             rd_resp_desc_1_xuser_15_reg <= 32'h0;
             wr_req_desc_1_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_1_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_1_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_1_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_1_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_1_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_1_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_1_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_1_resp_reg <= 32'h0;
             wr_resp_desc_1_xid_0_reg <= 32'h0;
             wr_resp_desc_1_xid_1_reg <= 32'h0;
             wr_resp_desc_1_xid_2_reg <= 32'h0;
             wr_resp_desc_1_xid_3_reg <= 32'h0;
             wr_resp_desc_1_xuser_0_reg <= 32'h0;
             wr_resp_desc_1_xuser_1_reg <= 32'h0;
             wr_resp_desc_1_xuser_2_reg <= 32'h0;
             wr_resp_desc_1_xuser_3_reg <= 32'h0;
             wr_resp_desc_1_xuser_4_reg <= 32'h0;
             wr_resp_desc_1_xuser_5_reg <= 32'h0;
             wr_resp_desc_1_xuser_6_reg <= 32'h0;
             wr_resp_desc_1_xuser_7_reg <= 32'h0;
             wr_resp_desc_1_xuser_8_reg <= 32'h0;
             wr_resp_desc_1_xuser_9_reg <= 32'h0;
             wr_resp_desc_1_xuser_10_reg <= 32'h0;
             wr_resp_desc_1_xuser_11_reg <= 32'h0;
             wr_resp_desc_1_xuser_12_reg <= 32'h0;
             wr_resp_desc_1_xuser_13_reg <= 32'h0;
             wr_resp_desc_1_xuser_14_reg <= 32'h0;
             wr_resp_desc_1_xuser_15_reg <= 32'h0;
             sn_req_desc_1_attr_reg <= 32'h0;
             sn_req_desc_1_acaddr_0_reg <= 32'h0;
             sn_req_desc_1_acaddr_1_reg <= 32'h0;
             sn_req_desc_1_acaddr_2_reg <= 32'h0;
             sn_req_desc_1_acaddr_3_reg <= 32'h0;
             rd_resp_desc_2_data_offset_reg <= 32'h0;
             rd_resp_desc_2_data_size_reg <= 32'h0;
             rd_resp_desc_2_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_2_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_2_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_2_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_2_resp_reg <= 32'h0;
             rd_resp_desc_2_xid_0_reg <= 32'h0;
             rd_resp_desc_2_xid_1_reg <= 32'h0;
             rd_resp_desc_2_xid_2_reg <= 32'h0;
             rd_resp_desc_2_xid_3_reg <= 32'h0;
             rd_resp_desc_2_xuser_0_reg <= 32'h0;
             rd_resp_desc_2_xuser_1_reg <= 32'h0;
             rd_resp_desc_2_xuser_2_reg <= 32'h0;
             rd_resp_desc_2_xuser_3_reg <= 32'h0;
             rd_resp_desc_2_xuser_4_reg <= 32'h0;
             rd_resp_desc_2_xuser_5_reg <= 32'h0;
             rd_resp_desc_2_xuser_6_reg <= 32'h0;
             rd_resp_desc_2_xuser_7_reg <= 32'h0;
             rd_resp_desc_2_xuser_8_reg <= 32'h0;
             rd_resp_desc_2_xuser_9_reg <= 32'h0;
             rd_resp_desc_2_xuser_10_reg <= 32'h0;
             rd_resp_desc_2_xuser_11_reg <= 32'h0;
             rd_resp_desc_2_xuser_12_reg <= 32'h0;
             rd_resp_desc_2_xuser_13_reg <= 32'h0;
             rd_resp_desc_2_xuser_14_reg <= 32'h0;
             rd_resp_desc_2_xuser_15_reg <= 32'h0;
             wr_req_desc_2_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_2_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_2_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_2_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_2_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_2_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_2_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_2_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_2_resp_reg <= 32'h0;
             wr_resp_desc_2_xid_0_reg <= 32'h0;
             wr_resp_desc_2_xid_1_reg <= 32'h0;
             wr_resp_desc_2_xid_2_reg <= 32'h0;
             wr_resp_desc_2_xid_3_reg <= 32'h0;
             wr_resp_desc_2_xuser_0_reg <= 32'h0;
             wr_resp_desc_2_xuser_1_reg <= 32'h0;
             wr_resp_desc_2_xuser_2_reg <= 32'h0;
             wr_resp_desc_2_xuser_3_reg <= 32'h0;
             wr_resp_desc_2_xuser_4_reg <= 32'h0;
             wr_resp_desc_2_xuser_5_reg <= 32'h0;
             wr_resp_desc_2_xuser_6_reg <= 32'h0;
             wr_resp_desc_2_xuser_7_reg <= 32'h0;
             wr_resp_desc_2_xuser_8_reg <= 32'h0;
             wr_resp_desc_2_xuser_9_reg <= 32'h0;
             wr_resp_desc_2_xuser_10_reg <= 32'h0;
             wr_resp_desc_2_xuser_11_reg <= 32'h0;
             wr_resp_desc_2_xuser_12_reg <= 32'h0;
             wr_resp_desc_2_xuser_13_reg <= 32'h0;
             wr_resp_desc_2_xuser_14_reg <= 32'h0;
             wr_resp_desc_2_xuser_15_reg <= 32'h0;
             sn_req_desc_2_attr_reg <= 32'h0;
             sn_req_desc_2_acaddr_0_reg <= 32'h0;
             sn_req_desc_2_acaddr_1_reg <= 32'h0;
             sn_req_desc_2_acaddr_2_reg <= 32'h0;
             sn_req_desc_2_acaddr_3_reg <= 32'h0;
             rd_resp_desc_3_data_offset_reg <= 32'h0;
             rd_resp_desc_3_data_size_reg <= 32'h0;
             rd_resp_desc_3_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_3_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_3_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_3_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_3_resp_reg <= 32'h0;
             rd_resp_desc_3_xid_0_reg <= 32'h0;
             rd_resp_desc_3_xid_1_reg <= 32'h0;
             rd_resp_desc_3_xid_2_reg <= 32'h0;
             rd_resp_desc_3_xid_3_reg <= 32'h0;
             rd_resp_desc_3_xuser_0_reg <= 32'h0;
             rd_resp_desc_3_xuser_1_reg <= 32'h0;
             rd_resp_desc_3_xuser_2_reg <= 32'h0;
             rd_resp_desc_3_xuser_3_reg <= 32'h0;
             rd_resp_desc_3_xuser_4_reg <= 32'h0;
             rd_resp_desc_3_xuser_5_reg <= 32'h0;
             rd_resp_desc_3_xuser_6_reg <= 32'h0;
             rd_resp_desc_3_xuser_7_reg <= 32'h0;
             rd_resp_desc_3_xuser_8_reg <= 32'h0;
             rd_resp_desc_3_xuser_9_reg <= 32'h0;
             rd_resp_desc_3_xuser_10_reg <= 32'h0;
             rd_resp_desc_3_xuser_11_reg <= 32'h0;
             rd_resp_desc_3_xuser_12_reg <= 32'h0;
             rd_resp_desc_3_xuser_13_reg <= 32'h0;
             rd_resp_desc_3_xuser_14_reg <= 32'h0;
             rd_resp_desc_3_xuser_15_reg <= 32'h0;
             wr_req_desc_3_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_3_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_3_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_3_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_3_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_3_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_3_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_3_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_3_resp_reg <= 32'h0;
             wr_resp_desc_3_xid_0_reg <= 32'h0;
             wr_resp_desc_3_xid_1_reg <= 32'h0;
             wr_resp_desc_3_xid_2_reg <= 32'h0;
             wr_resp_desc_3_xid_3_reg <= 32'h0;
             wr_resp_desc_3_xuser_0_reg <= 32'h0;
             wr_resp_desc_3_xuser_1_reg <= 32'h0;
             wr_resp_desc_3_xuser_2_reg <= 32'h0;
             wr_resp_desc_3_xuser_3_reg <= 32'h0;
             wr_resp_desc_3_xuser_4_reg <= 32'h0;
             wr_resp_desc_3_xuser_5_reg <= 32'h0;
             wr_resp_desc_3_xuser_6_reg <= 32'h0;
             wr_resp_desc_3_xuser_7_reg <= 32'h0;
             wr_resp_desc_3_xuser_8_reg <= 32'h0;
             wr_resp_desc_3_xuser_9_reg <= 32'h0;
             wr_resp_desc_3_xuser_10_reg <= 32'h0;
             wr_resp_desc_3_xuser_11_reg <= 32'h0;
             wr_resp_desc_3_xuser_12_reg <= 32'h0;
             wr_resp_desc_3_xuser_13_reg <= 32'h0;
             wr_resp_desc_3_xuser_14_reg <= 32'h0;
             wr_resp_desc_3_xuser_15_reg <= 32'h0;
             sn_req_desc_3_attr_reg <= 32'h0;
             sn_req_desc_3_acaddr_0_reg <= 32'h0;
             sn_req_desc_3_acaddr_1_reg <= 32'h0;
             sn_req_desc_3_acaddr_2_reg <= 32'h0;
             sn_req_desc_3_acaddr_3_reg <= 32'h0;
             rd_resp_desc_4_data_offset_reg <= 32'h0;
             rd_resp_desc_4_data_size_reg <= 32'h0;
             rd_resp_desc_4_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_4_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_4_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_4_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_4_resp_reg <= 32'h0;
             rd_resp_desc_4_xid_0_reg <= 32'h0;
             rd_resp_desc_4_xid_1_reg <= 32'h0;
             rd_resp_desc_4_xid_2_reg <= 32'h0;
             rd_resp_desc_4_xid_3_reg <= 32'h0;
             rd_resp_desc_4_xuser_0_reg <= 32'h0;
             rd_resp_desc_4_xuser_1_reg <= 32'h0;
             rd_resp_desc_4_xuser_2_reg <= 32'h0;
             rd_resp_desc_4_xuser_3_reg <= 32'h0;
             rd_resp_desc_4_xuser_4_reg <= 32'h0;
             rd_resp_desc_4_xuser_5_reg <= 32'h0;
             rd_resp_desc_4_xuser_6_reg <= 32'h0;
             rd_resp_desc_4_xuser_7_reg <= 32'h0;
             rd_resp_desc_4_xuser_8_reg <= 32'h0;
             rd_resp_desc_4_xuser_9_reg <= 32'h0;
             rd_resp_desc_4_xuser_10_reg <= 32'h0;
             rd_resp_desc_4_xuser_11_reg <= 32'h0;
             rd_resp_desc_4_xuser_12_reg <= 32'h0;
             rd_resp_desc_4_xuser_13_reg <= 32'h0;
             rd_resp_desc_4_xuser_14_reg <= 32'h0;
             rd_resp_desc_4_xuser_15_reg <= 32'h0;
             wr_req_desc_4_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_4_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_4_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_4_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_4_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_4_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_4_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_4_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_4_resp_reg <= 32'h0;
             wr_resp_desc_4_xid_0_reg <= 32'h0;
             wr_resp_desc_4_xid_1_reg <= 32'h0;
             wr_resp_desc_4_xid_2_reg <= 32'h0;
             wr_resp_desc_4_xid_3_reg <= 32'h0;
             wr_resp_desc_4_xuser_0_reg <= 32'h0;
             wr_resp_desc_4_xuser_1_reg <= 32'h0;
             wr_resp_desc_4_xuser_2_reg <= 32'h0;
             wr_resp_desc_4_xuser_3_reg <= 32'h0;
             wr_resp_desc_4_xuser_4_reg <= 32'h0;
             wr_resp_desc_4_xuser_5_reg <= 32'h0;
             wr_resp_desc_4_xuser_6_reg <= 32'h0;
             wr_resp_desc_4_xuser_7_reg <= 32'h0;
             wr_resp_desc_4_xuser_8_reg <= 32'h0;
             wr_resp_desc_4_xuser_9_reg <= 32'h0;
             wr_resp_desc_4_xuser_10_reg <= 32'h0;
             wr_resp_desc_4_xuser_11_reg <= 32'h0;
             wr_resp_desc_4_xuser_12_reg <= 32'h0;
             wr_resp_desc_4_xuser_13_reg <= 32'h0;
             wr_resp_desc_4_xuser_14_reg <= 32'h0;
             wr_resp_desc_4_xuser_15_reg <= 32'h0;
             sn_req_desc_4_attr_reg <= 32'h0;
             sn_req_desc_4_acaddr_0_reg <= 32'h0;
             sn_req_desc_4_acaddr_1_reg <= 32'h0;
             sn_req_desc_4_acaddr_2_reg <= 32'h0;
             sn_req_desc_4_acaddr_3_reg <= 32'h0;
             rd_resp_desc_5_data_offset_reg <= 32'h0;
             rd_resp_desc_5_data_size_reg <= 32'h0;
             rd_resp_desc_5_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_5_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_5_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_5_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_5_resp_reg <= 32'h0;
             rd_resp_desc_5_xid_0_reg <= 32'h0;
             rd_resp_desc_5_xid_1_reg <= 32'h0;
             rd_resp_desc_5_xid_2_reg <= 32'h0;
             rd_resp_desc_5_xid_3_reg <= 32'h0;
             rd_resp_desc_5_xuser_0_reg <= 32'h0;
             rd_resp_desc_5_xuser_1_reg <= 32'h0;
             rd_resp_desc_5_xuser_2_reg <= 32'h0;
             rd_resp_desc_5_xuser_3_reg <= 32'h0;
             rd_resp_desc_5_xuser_4_reg <= 32'h0;
             rd_resp_desc_5_xuser_5_reg <= 32'h0;
             rd_resp_desc_5_xuser_6_reg <= 32'h0;
             rd_resp_desc_5_xuser_7_reg <= 32'h0;
             rd_resp_desc_5_xuser_8_reg <= 32'h0;
             rd_resp_desc_5_xuser_9_reg <= 32'h0;
             rd_resp_desc_5_xuser_10_reg <= 32'h0;
             rd_resp_desc_5_xuser_11_reg <= 32'h0;
             rd_resp_desc_5_xuser_12_reg <= 32'h0;
             rd_resp_desc_5_xuser_13_reg <= 32'h0;
             rd_resp_desc_5_xuser_14_reg <= 32'h0;
             rd_resp_desc_5_xuser_15_reg <= 32'h0;
             wr_req_desc_5_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_5_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_5_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_5_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_5_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_5_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_5_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_5_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_5_resp_reg <= 32'h0;
             wr_resp_desc_5_xid_0_reg <= 32'h0;
             wr_resp_desc_5_xid_1_reg <= 32'h0;
             wr_resp_desc_5_xid_2_reg <= 32'h0;
             wr_resp_desc_5_xid_3_reg <= 32'h0;
             wr_resp_desc_5_xuser_0_reg <= 32'h0;
             wr_resp_desc_5_xuser_1_reg <= 32'h0;
             wr_resp_desc_5_xuser_2_reg <= 32'h0;
             wr_resp_desc_5_xuser_3_reg <= 32'h0;
             wr_resp_desc_5_xuser_4_reg <= 32'h0;
             wr_resp_desc_5_xuser_5_reg <= 32'h0;
             wr_resp_desc_5_xuser_6_reg <= 32'h0;
             wr_resp_desc_5_xuser_7_reg <= 32'h0;
             wr_resp_desc_5_xuser_8_reg <= 32'h0;
             wr_resp_desc_5_xuser_9_reg <= 32'h0;
             wr_resp_desc_5_xuser_10_reg <= 32'h0;
             wr_resp_desc_5_xuser_11_reg <= 32'h0;
             wr_resp_desc_5_xuser_12_reg <= 32'h0;
             wr_resp_desc_5_xuser_13_reg <= 32'h0;
             wr_resp_desc_5_xuser_14_reg <= 32'h0;
             wr_resp_desc_5_xuser_15_reg <= 32'h0;
             sn_req_desc_5_attr_reg <= 32'h0;
             sn_req_desc_5_acaddr_0_reg <= 32'h0;
             sn_req_desc_5_acaddr_1_reg <= 32'h0;
             sn_req_desc_5_acaddr_2_reg <= 32'h0;
             sn_req_desc_5_acaddr_3_reg <= 32'h0;
             rd_resp_desc_6_data_offset_reg <= 32'h0;
             rd_resp_desc_6_data_size_reg <= 32'h0;
             rd_resp_desc_6_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_6_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_6_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_6_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_6_resp_reg <= 32'h0;
             rd_resp_desc_6_xid_0_reg <= 32'h0;
             rd_resp_desc_6_xid_1_reg <= 32'h0;
             rd_resp_desc_6_xid_2_reg <= 32'h0;
             rd_resp_desc_6_xid_3_reg <= 32'h0;
             rd_resp_desc_6_xuser_0_reg <= 32'h0;
             rd_resp_desc_6_xuser_1_reg <= 32'h0;
             rd_resp_desc_6_xuser_2_reg <= 32'h0;
             rd_resp_desc_6_xuser_3_reg <= 32'h0;
             rd_resp_desc_6_xuser_4_reg <= 32'h0;
             rd_resp_desc_6_xuser_5_reg <= 32'h0;
             rd_resp_desc_6_xuser_6_reg <= 32'h0;
             rd_resp_desc_6_xuser_7_reg <= 32'h0;
             rd_resp_desc_6_xuser_8_reg <= 32'h0;
             rd_resp_desc_6_xuser_9_reg <= 32'h0;
             rd_resp_desc_6_xuser_10_reg <= 32'h0;
             rd_resp_desc_6_xuser_11_reg <= 32'h0;
             rd_resp_desc_6_xuser_12_reg <= 32'h0;
             rd_resp_desc_6_xuser_13_reg <= 32'h0;
             rd_resp_desc_6_xuser_14_reg <= 32'h0;
             rd_resp_desc_6_xuser_15_reg <= 32'h0;
             wr_req_desc_6_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_6_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_6_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_6_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_6_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_6_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_6_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_6_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_6_resp_reg <= 32'h0;
             wr_resp_desc_6_xid_0_reg <= 32'h0;
             wr_resp_desc_6_xid_1_reg <= 32'h0;
             wr_resp_desc_6_xid_2_reg <= 32'h0;
             wr_resp_desc_6_xid_3_reg <= 32'h0;
             wr_resp_desc_6_xuser_0_reg <= 32'h0;
             wr_resp_desc_6_xuser_1_reg <= 32'h0;
             wr_resp_desc_6_xuser_2_reg <= 32'h0;
             wr_resp_desc_6_xuser_3_reg <= 32'h0;
             wr_resp_desc_6_xuser_4_reg <= 32'h0;
             wr_resp_desc_6_xuser_5_reg <= 32'h0;
             wr_resp_desc_6_xuser_6_reg <= 32'h0;
             wr_resp_desc_6_xuser_7_reg <= 32'h0;
             wr_resp_desc_6_xuser_8_reg <= 32'h0;
             wr_resp_desc_6_xuser_9_reg <= 32'h0;
             wr_resp_desc_6_xuser_10_reg <= 32'h0;
             wr_resp_desc_6_xuser_11_reg <= 32'h0;
             wr_resp_desc_6_xuser_12_reg <= 32'h0;
             wr_resp_desc_6_xuser_13_reg <= 32'h0;
             wr_resp_desc_6_xuser_14_reg <= 32'h0;
             wr_resp_desc_6_xuser_15_reg <= 32'h0;
             sn_req_desc_6_attr_reg <= 32'h0;
             sn_req_desc_6_acaddr_0_reg <= 32'h0;
             sn_req_desc_6_acaddr_1_reg <= 32'h0;
             sn_req_desc_6_acaddr_2_reg <= 32'h0;
             sn_req_desc_6_acaddr_3_reg <= 32'h0;
             rd_resp_desc_7_data_offset_reg <= 32'h0;
             rd_resp_desc_7_data_size_reg <= 32'h0;
             rd_resp_desc_7_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_7_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_7_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_7_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_7_resp_reg <= 32'h0;
             rd_resp_desc_7_xid_0_reg <= 32'h0;
             rd_resp_desc_7_xid_1_reg <= 32'h0;
             rd_resp_desc_7_xid_2_reg <= 32'h0;
             rd_resp_desc_7_xid_3_reg <= 32'h0;
             rd_resp_desc_7_xuser_0_reg <= 32'h0;
             rd_resp_desc_7_xuser_1_reg <= 32'h0;
             rd_resp_desc_7_xuser_2_reg <= 32'h0;
             rd_resp_desc_7_xuser_3_reg <= 32'h0;
             rd_resp_desc_7_xuser_4_reg <= 32'h0;
             rd_resp_desc_7_xuser_5_reg <= 32'h0;
             rd_resp_desc_7_xuser_6_reg <= 32'h0;
             rd_resp_desc_7_xuser_7_reg <= 32'h0;
             rd_resp_desc_7_xuser_8_reg <= 32'h0;
             rd_resp_desc_7_xuser_9_reg <= 32'h0;
             rd_resp_desc_7_xuser_10_reg <= 32'h0;
             rd_resp_desc_7_xuser_11_reg <= 32'h0;
             rd_resp_desc_7_xuser_12_reg <= 32'h0;
             rd_resp_desc_7_xuser_13_reg <= 32'h0;
             rd_resp_desc_7_xuser_14_reg <= 32'h0;
             rd_resp_desc_7_xuser_15_reg <= 32'h0;
             wr_req_desc_7_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_7_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_7_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_7_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_7_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_7_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_7_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_7_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_7_resp_reg <= 32'h0;
             wr_resp_desc_7_xid_0_reg <= 32'h0;
             wr_resp_desc_7_xid_1_reg <= 32'h0;
             wr_resp_desc_7_xid_2_reg <= 32'h0;
             wr_resp_desc_7_xid_3_reg <= 32'h0;
             wr_resp_desc_7_xuser_0_reg <= 32'h0;
             wr_resp_desc_7_xuser_1_reg <= 32'h0;
             wr_resp_desc_7_xuser_2_reg <= 32'h0;
             wr_resp_desc_7_xuser_3_reg <= 32'h0;
             wr_resp_desc_7_xuser_4_reg <= 32'h0;
             wr_resp_desc_7_xuser_5_reg <= 32'h0;
             wr_resp_desc_7_xuser_6_reg <= 32'h0;
             wr_resp_desc_7_xuser_7_reg <= 32'h0;
             wr_resp_desc_7_xuser_8_reg <= 32'h0;
             wr_resp_desc_7_xuser_9_reg <= 32'h0;
             wr_resp_desc_7_xuser_10_reg <= 32'h0;
             wr_resp_desc_7_xuser_11_reg <= 32'h0;
             wr_resp_desc_7_xuser_12_reg <= 32'h0;
             wr_resp_desc_7_xuser_13_reg <= 32'h0;
             wr_resp_desc_7_xuser_14_reg <= 32'h0;
             wr_resp_desc_7_xuser_15_reg <= 32'h0;
             sn_req_desc_7_attr_reg <= 32'h0;
             sn_req_desc_7_acaddr_0_reg <= 32'h0;
             sn_req_desc_7_acaddr_1_reg <= 32'h0;
             sn_req_desc_7_acaddr_2_reg <= 32'h0;
             sn_req_desc_7_acaddr_3_reg <= 32'h0;
             rd_resp_desc_8_data_offset_reg <= 32'h0;
             rd_resp_desc_8_data_size_reg <= 32'h0;
             rd_resp_desc_8_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_8_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_8_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_8_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_8_resp_reg <= 32'h0;
             rd_resp_desc_8_xid_0_reg <= 32'h0;
             rd_resp_desc_8_xid_1_reg <= 32'h0;
             rd_resp_desc_8_xid_2_reg <= 32'h0;
             rd_resp_desc_8_xid_3_reg <= 32'h0;
             rd_resp_desc_8_xuser_0_reg <= 32'h0;
             rd_resp_desc_8_xuser_1_reg <= 32'h0;
             rd_resp_desc_8_xuser_2_reg <= 32'h0;
             rd_resp_desc_8_xuser_3_reg <= 32'h0;
             rd_resp_desc_8_xuser_4_reg <= 32'h0;
             rd_resp_desc_8_xuser_5_reg <= 32'h0;
             rd_resp_desc_8_xuser_6_reg <= 32'h0;
             rd_resp_desc_8_xuser_7_reg <= 32'h0;
             rd_resp_desc_8_xuser_8_reg <= 32'h0;
             rd_resp_desc_8_xuser_9_reg <= 32'h0;
             rd_resp_desc_8_xuser_10_reg <= 32'h0;
             rd_resp_desc_8_xuser_11_reg <= 32'h0;
             rd_resp_desc_8_xuser_12_reg <= 32'h0;
             rd_resp_desc_8_xuser_13_reg <= 32'h0;
             rd_resp_desc_8_xuser_14_reg <= 32'h0;
             rd_resp_desc_8_xuser_15_reg <= 32'h0;
             wr_req_desc_8_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_8_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_8_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_8_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_8_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_8_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_8_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_8_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_8_resp_reg <= 32'h0;
             wr_resp_desc_8_xid_0_reg <= 32'h0;
             wr_resp_desc_8_xid_1_reg <= 32'h0;
             wr_resp_desc_8_xid_2_reg <= 32'h0;
             wr_resp_desc_8_xid_3_reg <= 32'h0;
             wr_resp_desc_8_xuser_0_reg <= 32'h0;
             wr_resp_desc_8_xuser_1_reg <= 32'h0;
             wr_resp_desc_8_xuser_2_reg <= 32'h0;
             wr_resp_desc_8_xuser_3_reg <= 32'h0;
             wr_resp_desc_8_xuser_4_reg <= 32'h0;
             wr_resp_desc_8_xuser_5_reg <= 32'h0;
             wr_resp_desc_8_xuser_6_reg <= 32'h0;
             wr_resp_desc_8_xuser_7_reg <= 32'h0;
             wr_resp_desc_8_xuser_8_reg <= 32'h0;
             wr_resp_desc_8_xuser_9_reg <= 32'h0;
             wr_resp_desc_8_xuser_10_reg <= 32'h0;
             wr_resp_desc_8_xuser_11_reg <= 32'h0;
             wr_resp_desc_8_xuser_12_reg <= 32'h0;
             wr_resp_desc_8_xuser_13_reg <= 32'h0;
             wr_resp_desc_8_xuser_14_reg <= 32'h0;
             wr_resp_desc_8_xuser_15_reg <= 32'h0;
             sn_req_desc_8_attr_reg <= 32'h0;
             sn_req_desc_8_acaddr_0_reg <= 32'h0;
             sn_req_desc_8_acaddr_1_reg <= 32'h0;
             sn_req_desc_8_acaddr_2_reg <= 32'h0;
             sn_req_desc_8_acaddr_3_reg <= 32'h0;
             rd_resp_desc_9_data_offset_reg <= 32'h0;
             rd_resp_desc_9_data_size_reg <= 32'h0;
             rd_resp_desc_9_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_9_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_9_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_9_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_9_resp_reg <= 32'h0;
             rd_resp_desc_9_xid_0_reg <= 32'h0;
             rd_resp_desc_9_xid_1_reg <= 32'h0;
             rd_resp_desc_9_xid_2_reg <= 32'h0;
             rd_resp_desc_9_xid_3_reg <= 32'h0;
             rd_resp_desc_9_xuser_0_reg <= 32'h0;
             rd_resp_desc_9_xuser_1_reg <= 32'h0;
             rd_resp_desc_9_xuser_2_reg <= 32'h0;
             rd_resp_desc_9_xuser_3_reg <= 32'h0;
             rd_resp_desc_9_xuser_4_reg <= 32'h0;
             rd_resp_desc_9_xuser_5_reg <= 32'h0;
             rd_resp_desc_9_xuser_6_reg <= 32'h0;
             rd_resp_desc_9_xuser_7_reg <= 32'h0;
             rd_resp_desc_9_xuser_8_reg <= 32'h0;
             rd_resp_desc_9_xuser_9_reg <= 32'h0;
             rd_resp_desc_9_xuser_10_reg <= 32'h0;
             rd_resp_desc_9_xuser_11_reg <= 32'h0;
             rd_resp_desc_9_xuser_12_reg <= 32'h0;
             rd_resp_desc_9_xuser_13_reg <= 32'h0;
             rd_resp_desc_9_xuser_14_reg <= 32'h0;
             rd_resp_desc_9_xuser_15_reg <= 32'h0;
             wr_req_desc_9_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_9_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_9_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_9_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_9_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_9_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_9_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_9_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_9_resp_reg <= 32'h0;
             wr_resp_desc_9_xid_0_reg <= 32'h0;
             wr_resp_desc_9_xid_1_reg <= 32'h0;
             wr_resp_desc_9_xid_2_reg <= 32'h0;
             wr_resp_desc_9_xid_3_reg <= 32'h0;
             wr_resp_desc_9_xuser_0_reg <= 32'h0;
             wr_resp_desc_9_xuser_1_reg <= 32'h0;
             wr_resp_desc_9_xuser_2_reg <= 32'h0;
             wr_resp_desc_9_xuser_3_reg <= 32'h0;
             wr_resp_desc_9_xuser_4_reg <= 32'h0;
             wr_resp_desc_9_xuser_5_reg <= 32'h0;
             wr_resp_desc_9_xuser_6_reg <= 32'h0;
             wr_resp_desc_9_xuser_7_reg <= 32'h0;
             wr_resp_desc_9_xuser_8_reg <= 32'h0;
             wr_resp_desc_9_xuser_9_reg <= 32'h0;
             wr_resp_desc_9_xuser_10_reg <= 32'h0;
             wr_resp_desc_9_xuser_11_reg <= 32'h0;
             wr_resp_desc_9_xuser_12_reg <= 32'h0;
             wr_resp_desc_9_xuser_13_reg <= 32'h0;
             wr_resp_desc_9_xuser_14_reg <= 32'h0;
             wr_resp_desc_9_xuser_15_reg <= 32'h0;
             sn_req_desc_9_attr_reg <= 32'h0;
             sn_req_desc_9_acaddr_0_reg <= 32'h0;
             sn_req_desc_9_acaddr_1_reg <= 32'h0;
             sn_req_desc_9_acaddr_2_reg <= 32'h0;
             sn_req_desc_9_acaddr_3_reg <= 32'h0;
             rd_resp_desc_a_data_offset_reg <= 32'h0;
             rd_resp_desc_a_data_size_reg <= 32'h0;
             rd_resp_desc_a_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_a_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_a_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_a_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_a_resp_reg <= 32'h0;
             rd_resp_desc_a_xid_0_reg <= 32'h0;
             rd_resp_desc_a_xid_1_reg <= 32'h0;
             rd_resp_desc_a_xid_2_reg <= 32'h0;
             rd_resp_desc_a_xid_3_reg <= 32'h0;
             rd_resp_desc_a_xuser_0_reg <= 32'h0;
             rd_resp_desc_a_xuser_1_reg <= 32'h0;
             rd_resp_desc_a_xuser_2_reg <= 32'h0;
             rd_resp_desc_a_xuser_3_reg <= 32'h0;
             rd_resp_desc_a_xuser_4_reg <= 32'h0;
             rd_resp_desc_a_xuser_5_reg <= 32'h0;
             rd_resp_desc_a_xuser_6_reg <= 32'h0;
             rd_resp_desc_a_xuser_7_reg <= 32'h0;
             rd_resp_desc_a_xuser_8_reg <= 32'h0;
             rd_resp_desc_a_xuser_9_reg <= 32'h0;
             rd_resp_desc_a_xuser_10_reg <= 32'h0;
             rd_resp_desc_a_xuser_11_reg <= 32'h0;
             rd_resp_desc_a_xuser_12_reg <= 32'h0;
             rd_resp_desc_a_xuser_13_reg <= 32'h0;
             rd_resp_desc_a_xuser_14_reg <= 32'h0;
             rd_resp_desc_a_xuser_15_reg <= 32'h0;
             wr_req_desc_a_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_a_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_a_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_a_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_a_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_a_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_a_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_a_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_a_resp_reg <= 32'h0;
             wr_resp_desc_a_xid_0_reg <= 32'h0;
             wr_resp_desc_a_xid_1_reg <= 32'h0;
             wr_resp_desc_a_xid_2_reg <= 32'h0;
             wr_resp_desc_a_xid_3_reg <= 32'h0;
             wr_resp_desc_a_xuser_0_reg <= 32'h0;
             wr_resp_desc_a_xuser_1_reg <= 32'h0;
             wr_resp_desc_a_xuser_2_reg <= 32'h0;
             wr_resp_desc_a_xuser_3_reg <= 32'h0;
             wr_resp_desc_a_xuser_4_reg <= 32'h0;
             wr_resp_desc_a_xuser_5_reg <= 32'h0;
             wr_resp_desc_a_xuser_6_reg <= 32'h0;
             wr_resp_desc_a_xuser_7_reg <= 32'h0;
             wr_resp_desc_a_xuser_8_reg <= 32'h0;
             wr_resp_desc_a_xuser_9_reg <= 32'h0;
             wr_resp_desc_a_xuser_10_reg <= 32'h0;
             wr_resp_desc_a_xuser_11_reg <= 32'h0;
             wr_resp_desc_a_xuser_12_reg <= 32'h0;
             wr_resp_desc_a_xuser_13_reg <= 32'h0;
             wr_resp_desc_a_xuser_14_reg <= 32'h0;
             wr_resp_desc_a_xuser_15_reg <= 32'h0;
             sn_req_desc_a_attr_reg <= 32'h0;
             sn_req_desc_a_acaddr_0_reg <= 32'h0;
             sn_req_desc_a_acaddr_1_reg <= 32'h0;
             sn_req_desc_a_acaddr_2_reg <= 32'h0;
             sn_req_desc_a_acaddr_3_reg <= 32'h0;
             rd_resp_desc_b_data_offset_reg <= 32'h0;
             rd_resp_desc_b_data_size_reg <= 32'h0;
             rd_resp_desc_b_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_b_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_b_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_b_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_b_resp_reg <= 32'h0;
             rd_resp_desc_b_xid_0_reg <= 32'h0;
             rd_resp_desc_b_xid_1_reg <= 32'h0;
             rd_resp_desc_b_xid_2_reg <= 32'h0;
             rd_resp_desc_b_xid_3_reg <= 32'h0;
             rd_resp_desc_b_xuser_0_reg <= 32'h0;
             rd_resp_desc_b_xuser_1_reg <= 32'h0;
             rd_resp_desc_b_xuser_2_reg <= 32'h0;
             rd_resp_desc_b_xuser_3_reg <= 32'h0;
             rd_resp_desc_b_xuser_4_reg <= 32'h0;
             rd_resp_desc_b_xuser_5_reg <= 32'h0;
             rd_resp_desc_b_xuser_6_reg <= 32'h0;
             rd_resp_desc_b_xuser_7_reg <= 32'h0;
             rd_resp_desc_b_xuser_8_reg <= 32'h0;
             rd_resp_desc_b_xuser_9_reg <= 32'h0;
             rd_resp_desc_b_xuser_10_reg <= 32'h0;
             rd_resp_desc_b_xuser_11_reg <= 32'h0;
             rd_resp_desc_b_xuser_12_reg <= 32'h0;
             rd_resp_desc_b_xuser_13_reg <= 32'h0;
             rd_resp_desc_b_xuser_14_reg <= 32'h0;
             rd_resp_desc_b_xuser_15_reg <= 32'h0;
             wr_req_desc_b_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_b_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_b_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_b_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_b_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_b_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_b_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_b_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_b_resp_reg <= 32'h0;
             wr_resp_desc_b_xid_0_reg <= 32'h0;
             wr_resp_desc_b_xid_1_reg <= 32'h0;
             wr_resp_desc_b_xid_2_reg <= 32'h0;
             wr_resp_desc_b_xid_3_reg <= 32'h0;
             wr_resp_desc_b_xuser_0_reg <= 32'h0;
             wr_resp_desc_b_xuser_1_reg <= 32'h0;
             wr_resp_desc_b_xuser_2_reg <= 32'h0;
             wr_resp_desc_b_xuser_3_reg <= 32'h0;
             wr_resp_desc_b_xuser_4_reg <= 32'h0;
             wr_resp_desc_b_xuser_5_reg <= 32'h0;
             wr_resp_desc_b_xuser_6_reg <= 32'h0;
             wr_resp_desc_b_xuser_7_reg <= 32'h0;
             wr_resp_desc_b_xuser_8_reg <= 32'h0;
             wr_resp_desc_b_xuser_9_reg <= 32'h0;
             wr_resp_desc_b_xuser_10_reg <= 32'h0;
             wr_resp_desc_b_xuser_11_reg <= 32'h0;
             wr_resp_desc_b_xuser_12_reg <= 32'h0;
             wr_resp_desc_b_xuser_13_reg <= 32'h0;
             wr_resp_desc_b_xuser_14_reg <= 32'h0;
             wr_resp_desc_b_xuser_15_reg <= 32'h0;
             sn_req_desc_b_attr_reg <= 32'h0;
             sn_req_desc_b_acaddr_0_reg <= 32'h0;
             sn_req_desc_b_acaddr_1_reg <= 32'h0;
             sn_req_desc_b_acaddr_2_reg <= 32'h0;
             sn_req_desc_b_acaddr_3_reg <= 32'h0;
             rd_resp_desc_c_data_offset_reg <= 32'h0;
             rd_resp_desc_c_data_size_reg <= 32'h0;
             rd_resp_desc_c_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_c_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_c_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_c_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_c_resp_reg <= 32'h0;
             rd_resp_desc_c_xid_0_reg <= 32'h0;
             rd_resp_desc_c_xid_1_reg <= 32'h0;
             rd_resp_desc_c_xid_2_reg <= 32'h0;
             rd_resp_desc_c_xid_3_reg <= 32'h0;
             rd_resp_desc_c_xuser_0_reg <= 32'h0;
             rd_resp_desc_c_xuser_1_reg <= 32'h0;
             rd_resp_desc_c_xuser_2_reg <= 32'h0;
             rd_resp_desc_c_xuser_3_reg <= 32'h0;
             rd_resp_desc_c_xuser_4_reg <= 32'h0;
             rd_resp_desc_c_xuser_5_reg <= 32'h0;
             rd_resp_desc_c_xuser_6_reg <= 32'h0;
             rd_resp_desc_c_xuser_7_reg <= 32'h0;
             rd_resp_desc_c_xuser_8_reg <= 32'h0;
             rd_resp_desc_c_xuser_9_reg <= 32'h0;
             rd_resp_desc_c_xuser_10_reg <= 32'h0;
             rd_resp_desc_c_xuser_11_reg <= 32'h0;
             rd_resp_desc_c_xuser_12_reg <= 32'h0;
             rd_resp_desc_c_xuser_13_reg <= 32'h0;
             rd_resp_desc_c_xuser_14_reg <= 32'h0;
             rd_resp_desc_c_xuser_15_reg <= 32'h0;
             wr_req_desc_c_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_c_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_c_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_c_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_c_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_c_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_c_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_c_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_c_resp_reg <= 32'h0;
             wr_resp_desc_c_xid_0_reg <= 32'h0;
             wr_resp_desc_c_xid_1_reg <= 32'h0;
             wr_resp_desc_c_xid_2_reg <= 32'h0;
             wr_resp_desc_c_xid_3_reg <= 32'h0;
             wr_resp_desc_c_xuser_0_reg <= 32'h0;
             wr_resp_desc_c_xuser_1_reg <= 32'h0;
             wr_resp_desc_c_xuser_2_reg <= 32'h0;
             wr_resp_desc_c_xuser_3_reg <= 32'h0;
             wr_resp_desc_c_xuser_4_reg <= 32'h0;
             wr_resp_desc_c_xuser_5_reg <= 32'h0;
             wr_resp_desc_c_xuser_6_reg <= 32'h0;
             wr_resp_desc_c_xuser_7_reg <= 32'h0;
             wr_resp_desc_c_xuser_8_reg <= 32'h0;
             wr_resp_desc_c_xuser_9_reg <= 32'h0;
             wr_resp_desc_c_xuser_10_reg <= 32'h0;
             wr_resp_desc_c_xuser_11_reg <= 32'h0;
             wr_resp_desc_c_xuser_12_reg <= 32'h0;
             wr_resp_desc_c_xuser_13_reg <= 32'h0;
             wr_resp_desc_c_xuser_14_reg <= 32'h0;
             wr_resp_desc_c_xuser_15_reg <= 32'h0;
             sn_req_desc_c_attr_reg <= 32'h0;
             sn_req_desc_c_acaddr_0_reg <= 32'h0;
             sn_req_desc_c_acaddr_1_reg <= 32'h0;
             sn_req_desc_c_acaddr_2_reg <= 32'h0;
             sn_req_desc_c_acaddr_3_reg <= 32'h0;
             rd_resp_desc_d_data_offset_reg <= 32'h0;
             rd_resp_desc_d_data_size_reg <= 32'h0;
             rd_resp_desc_d_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_d_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_d_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_d_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_d_resp_reg <= 32'h0;
             rd_resp_desc_d_xid_0_reg <= 32'h0;
             rd_resp_desc_d_xid_1_reg <= 32'h0;
             rd_resp_desc_d_xid_2_reg <= 32'h0;
             rd_resp_desc_d_xid_3_reg <= 32'h0;
             rd_resp_desc_d_xuser_0_reg <= 32'h0;
             rd_resp_desc_d_xuser_1_reg <= 32'h0;
             rd_resp_desc_d_xuser_2_reg <= 32'h0;
             rd_resp_desc_d_xuser_3_reg <= 32'h0;
             rd_resp_desc_d_xuser_4_reg <= 32'h0;
             rd_resp_desc_d_xuser_5_reg <= 32'h0;
             rd_resp_desc_d_xuser_6_reg <= 32'h0;
             rd_resp_desc_d_xuser_7_reg <= 32'h0;
             rd_resp_desc_d_xuser_8_reg <= 32'h0;
             rd_resp_desc_d_xuser_9_reg <= 32'h0;
             rd_resp_desc_d_xuser_10_reg <= 32'h0;
             rd_resp_desc_d_xuser_11_reg <= 32'h0;
             rd_resp_desc_d_xuser_12_reg <= 32'h0;
             rd_resp_desc_d_xuser_13_reg <= 32'h0;
             rd_resp_desc_d_xuser_14_reg <= 32'h0;
             rd_resp_desc_d_xuser_15_reg <= 32'h0;
             wr_req_desc_d_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_d_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_d_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_d_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_d_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_d_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_d_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_d_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_d_resp_reg <= 32'h0;
             wr_resp_desc_d_xid_0_reg <= 32'h0;
             wr_resp_desc_d_xid_1_reg <= 32'h0;
             wr_resp_desc_d_xid_2_reg <= 32'h0;
             wr_resp_desc_d_xid_3_reg <= 32'h0;
             wr_resp_desc_d_xuser_0_reg <= 32'h0;
             wr_resp_desc_d_xuser_1_reg <= 32'h0;
             wr_resp_desc_d_xuser_2_reg <= 32'h0;
             wr_resp_desc_d_xuser_3_reg <= 32'h0;
             wr_resp_desc_d_xuser_4_reg <= 32'h0;
             wr_resp_desc_d_xuser_5_reg <= 32'h0;
             wr_resp_desc_d_xuser_6_reg <= 32'h0;
             wr_resp_desc_d_xuser_7_reg <= 32'h0;
             wr_resp_desc_d_xuser_8_reg <= 32'h0;
             wr_resp_desc_d_xuser_9_reg <= 32'h0;
             wr_resp_desc_d_xuser_10_reg <= 32'h0;
             wr_resp_desc_d_xuser_11_reg <= 32'h0;
             wr_resp_desc_d_xuser_12_reg <= 32'h0;
             wr_resp_desc_d_xuser_13_reg <= 32'h0;
             wr_resp_desc_d_xuser_14_reg <= 32'h0;
             wr_resp_desc_d_xuser_15_reg <= 32'h0;
             sn_req_desc_d_attr_reg <= 32'h0;
             sn_req_desc_d_acaddr_0_reg <= 32'h0;
             sn_req_desc_d_acaddr_1_reg <= 32'h0;
             sn_req_desc_d_acaddr_2_reg <= 32'h0;
             sn_req_desc_d_acaddr_3_reg <= 32'h0;
             rd_resp_desc_e_data_offset_reg <= 32'h0;
             rd_resp_desc_e_data_size_reg <= 32'h0;
             rd_resp_desc_e_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_e_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_e_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_e_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_e_resp_reg <= 32'h0;
             rd_resp_desc_e_xid_0_reg <= 32'h0;
             rd_resp_desc_e_xid_1_reg <= 32'h0;
             rd_resp_desc_e_xid_2_reg <= 32'h0;
             rd_resp_desc_e_xid_3_reg <= 32'h0;
             rd_resp_desc_e_xuser_0_reg <= 32'h0;
             rd_resp_desc_e_xuser_1_reg <= 32'h0;
             rd_resp_desc_e_xuser_2_reg <= 32'h0;
             rd_resp_desc_e_xuser_3_reg <= 32'h0;
             rd_resp_desc_e_xuser_4_reg <= 32'h0;
             rd_resp_desc_e_xuser_5_reg <= 32'h0;
             rd_resp_desc_e_xuser_6_reg <= 32'h0;
             rd_resp_desc_e_xuser_7_reg <= 32'h0;
             rd_resp_desc_e_xuser_8_reg <= 32'h0;
             rd_resp_desc_e_xuser_9_reg <= 32'h0;
             rd_resp_desc_e_xuser_10_reg <= 32'h0;
             rd_resp_desc_e_xuser_11_reg <= 32'h0;
             rd_resp_desc_e_xuser_12_reg <= 32'h0;
             rd_resp_desc_e_xuser_13_reg <= 32'h0;
             rd_resp_desc_e_xuser_14_reg <= 32'h0;
             rd_resp_desc_e_xuser_15_reg <= 32'h0;
             wr_req_desc_e_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_e_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_e_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_e_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_e_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_e_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_e_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_e_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_e_resp_reg <= 32'h0;
             wr_resp_desc_e_xid_0_reg <= 32'h0;
             wr_resp_desc_e_xid_1_reg <= 32'h0;
             wr_resp_desc_e_xid_2_reg <= 32'h0;
             wr_resp_desc_e_xid_3_reg <= 32'h0;
             wr_resp_desc_e_xuser_0_reg <= 32'h0;
             wr_resp_desc_e_xuser_1_reg <= 32'h0;
             wr_resp_desc_e_xuser_2_reg <= 32'h0;
             wr_resp_desc_e_xuser_3_reg <= 32'h0;
             wr_resp_desc_e_xuser_4_reg <= 32'h0;
             wr_resp_desc_e_xuser_5_reg <= 32'h0;
             wr_resp_desc_e_xuser_6_reg <= 32'h0;
             wr_resp_desc_e_xuser_7_reg <= 32'h0;
             wr_resp_desc_e_xuser_8_reg <= 32'h0;
             wr_resp_desc_e_xuser_9_reg <= 32'h0;
             wr_resp_desc_e_xuser_10_reg <= 32'h0;
             wr_resp_desc_e_xuser_11_reg <= 32'h0;
             wr_resp_desc_e_xuser_12_reg <= 32'h0;
             wr_resp_desc_e_xuser_13_reg <= 32'h0;
             wr_resp_desc_e_xuser_14_reg <= 32'h0;
             wr_resp_desc_e_xuser_15_reg <= 32'h0;
             sn_req_desc_e_attr_reg <= 32'h0;
             sn_req_desc_e_acaddr_0_reg <= 32'h0;
             sn_req_desc_e_acaddr_1_reg <= 32'h0;
             sn_req_desc_e_acaddr_2_reg <= 32'h0;
             sn_req_desc_e_acaddr_3_reg <= 32'h0;
             rd_resp_desc_f_data_offset_reg <= 32'h0;
             rd_resp_desc_f_data_size_reg <= 32'h0;
             rd_resp_desc_f_data_host_addr_0_reg <= 32'h0;
             rd_resp_desc_f_data_host_addr_1_reg <= 32'h0;
             rd_resp_desc_f_data_host_addr_2_reg <= 32'h0;
             rd_resp_desc_f_data_host_addr_3_reg <= 32'h0;
             rd_resp_desc_f_resp_reg <= 32'h0;
             rd_resp_desc_f_xid_0_reg <= 32'h0;
             rd_resp_desc_f_xid_1_reg <= 32'h0;
             rd_resp_desc_f_xid_2_reg <= 32'h0;
             rd_resp_desc_f_xid_3_reg <= 32'h0;
             rd_resp_desc_f_xuser_0_reg <= 32'h0;
             rd_resp_desc_f_xuser_1_reg <= 32'h0;
             rd_resp_desc_f_xuser_2_reg <= 32'h0;
             rd_resp_desc_f_xuser_3_reg <= 32'h0;
             rd_resp_desc_f_xuser_4_reg <= 32'h0;
             rd_resp_desc_f_xuser_5_reg <= 32'h0;
             rd_resp_desc_f_xuser_6_reg <= 32'h0;
             rd_resp_desc_f_xuser_7_reg <= 32'h0;
             rd_resp_desc_f_xuser_8_reg <= 32'h0;
             rd_resp_desc_f_xuser_9_reg <= 32'h0;
             rd_resp_desc_f_xuser_10_reg <= 32'h0;
             rd_resp_desc_f_xuser_11_reg <= 32'h0;
             rd_resp_desc_f_xuser_12_reg <= 32'h0;
             rd_resp_desc_f_xuser_13_reg <= 32'h0;
             rd_resp_desc_f_xuser_14_reg <= 32'h0;
             rd_resp_desc_f_xuser_15_reg <= 32'h0;
             wr_req_desc_f_data_host_addr_0_reg <= 32'h0;
             wr_req_desc_f_data_host_addr_1_reg <= 32'h0;
             wr_req_desc_f_data_host_addr_2_reg <= 32'h0;
             wr_req_desc_f_data_host_addr_3_reg <= 32'h0;
             wr_req_desc_f_wstrb_host_addr_0_reg <= 32'h0;
             wr_req_desc_f_wstrb_host_addr_1_reg <= 32'h0;
             wr_req_desc_f_wstrb_host_addr_2_reg <= 32'h0;
             wr_req_desc_f_wstrb_host_addr_3_reg <= 32'h0;
             wr_resp_desc_f_resp_reg <= 32'h0;
             wr_resp_desc_f_xid_0_reg <= 32'h0;
             wr_resp_desc_f_xid_1_reg <= 32'h0;
             wr_resp_desc_f_xid_2_reg <= 32'h0;
             wr_resp_desc_f_xid_3_reg <= 32'h0;
             wr_resp_desc_f_xuser_0_reg <= 32'h0;
             wr_resp_desc_f_xuser_1_reg <= 32'h0;
             wr_resp_desc_f_xuser_2_reg <= 32'h0;
             wr_resp_desc_f_xuser_3_reg <= 32'h0;
             wr_resp_desc_f_xuser_4_reg <= 32'h0;
             wr_resp_desc_f_xuser_5_reg <= 32'h0;
             wr_resp_desc_f_xuser_6_reg <= 32'h0;
             wr_resp_desc_f_xuser_7_reg <= 32'h0;
             wr_resp_desc_f_xuser_8_reg <= 32'h0;
             wr_resp_desc_f_xuser_9_reg <= 32'h0;
             wr_resp_desc_f_xuser_10_reg <= 32'h0;
             wr_resp_desc_f_xuser_11_reg <= 32'h0;
             wr_resp_desc_f_xuser_12_reg <= 32'h0;
             wr_resp_desc_f_xuser_13_reg <= 32'h0;
             wr_resp_desc_f_xuser_14_reg <= 32'h0;
             wr_resp_desc_f_xuser_15_reg <= 32'h0;
             sn_req_desc_f_attr_reg <= 32'h0;
             sn_req_desc_f_acaddr_0_reg <= 32'h0;
             sn_req_desc_f_acaddr_1_reg <= 32'h0;
             sn_req_desc_f_acaddr_2_reg <= 32'h0;
             sn_req_desc_f_acaddr_3_reg <= 32'h0;
             
             
          end
        else begin
           if (reg_wr_en)
             begin
                case (axi_awaddr[BRIDGE_MSB:0])  
                  
                  `MODE_SELECT_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         mode_select_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_INTR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_intr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_INTR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_intr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_INTR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_intr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_INTR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_intr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_C2H_TOGGLE_CLEAR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_c2h_toggle_clear_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_C2H_TOGGLE_ENABLE_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_c2h_toggle_enable_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_C2H_TOGGLE_CLEAR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_c2h_toggle_clear_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_C2H_TOGGLE_ENABLE_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_c2h_toggle_enable_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `H2C_GPIO_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         h2c_gpio_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_ERROR_CLEAR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_error_clear_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_ERROR_ENABLE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_error_enable_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_REQ_FREE_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_req_free_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_FIFO_PUSH_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_fifo_push_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_INTR_COMP_CLEAR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_intr_comp_clear_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_INTR_COMP_ENABLE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_intr_comp_enable_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_FREE_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_free_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_FIFO_PUSH_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_fifo_push_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_INTR_COMP_CLEAR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_intr_comp_clear_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_INTR_COMP_ENABLE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_intr_comp_enable_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_FIFO_PUSH_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_fifo_push_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_INTR_COMP_CLEAR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_intr_comp_clear_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_INTR_COMP_ENABLE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_intr_comp_enable_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_RESP_FREE_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_resp_free_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_DATA_FREE_DESC_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_data_free_desc_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `INTR_FIFO_ENABLE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         intr_fifo_enable_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_0_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_0_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_0_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_0_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_0_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_0_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_0_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_0_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_0_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_0_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_0_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_0_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_0_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_0_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_0_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_0_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_1_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_1_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_1_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_1_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_1_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_1_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_1_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_1_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_1_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_1_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_1_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_1_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_1_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_1_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_1_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_1_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_2_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_2_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_2_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_2_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_2_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_2_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_2_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_2_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_2_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_2_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_2_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_2_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_2_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_2_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_2_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_2_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_3_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_3_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_3_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_3_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_3_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_3_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_3_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_3_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_3_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_3_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_3_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_3_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_3_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_3_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_3_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_3_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_4_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_4_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_4_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_4_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_4_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_4_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_4_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_4_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_4_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_4_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_4_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_4_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_4_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_4_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_4_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_4_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_5_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_5_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_5_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_5_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_5_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_5_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_5_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_5_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_5_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_5_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_5_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_5_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_5_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_5_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_5_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_5_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_6_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_6_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_6_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_6_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_6_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_6_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_6_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_6_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_6_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_6_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_6_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_6_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_6_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_6_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_6_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_6_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_7_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_7_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_7_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_7_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_7_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_7_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_7_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_7_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_7_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_7_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_7_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_7_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_7_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_7_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_7_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_7_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_8_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_8_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_8_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_8_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_8_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_8_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_8_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_8_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_8_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_8_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_8_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_8_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_8_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_8_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_8_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_8_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_9_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_9_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_9_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_9_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_9_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_9_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_9_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_9_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_9_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_9_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_9_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_9_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_9_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_9_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_9_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_9_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_A_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_a_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_A_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_a_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_A_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_a_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_A_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_a_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_A_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_a_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_A_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_a_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_A_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_a_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_A_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_a_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_B_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_b_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_B_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_b_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_B_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_b_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_B_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_b_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_B_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_b_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_B_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_b_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_B_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_b_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_B_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_b_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_C_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_c_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_C_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_c_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_C_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_c_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_C_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_c_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_C_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_c_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_C_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_c_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_C_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_c_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_C_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_c_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_D_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_d_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_D_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_d_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_D_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_d_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_D_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_d_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_D_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_d_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_D_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_d_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_D_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_d_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_D_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_d_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_E_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_e_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_E_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_e_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_E_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_e_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_E_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_e_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_E_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_e_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_E_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_e_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_E_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_e_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_E_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_e_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_DATA_OFFSET_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_data_offset_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_DATA_SIZE_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_data_size_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `RD_RESP_DESC_F_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         rd_resp_desc_f_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_DATA_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_data_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_DATA_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_data_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_DATA_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_data_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_DATA_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_data_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_WSTRB_HOST_ADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_wstrb_host_addr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_WSTRB_HOST_ADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_wstrb_host_addr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_WSTRB_HOST_ADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_wstrb_host_addr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_REQ_DESC_F_WSTRB_HOST_ADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_req_desc_f_wstrb_host_addr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_RESP_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_resp_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XID_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xid_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XID_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xid_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XID_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xid_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XID_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xid_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_4_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_4_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_5_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_5_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_6_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_6_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_7_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_7_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_8_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_8_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_9_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_9_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_10_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_10_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_11_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_11_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_12_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_12_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_13_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_13_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_14_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_14_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `WR_RESP_DESC_F_XUSER_15_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         wr_resp_desc_f_xuser_15_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_F_ATTR_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_f_attr_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_F_ACADDR_0_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_f_acaddr_0_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_F_ACADDR_1_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_f_acaddr_1_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_F_ACADDR_2_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_f_acaddr_2_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
                  `SN_REQ_DESC_F_ACADDR_3_REG_ADDR:
                    for ( byte_index = 0; byte_index <= (S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
                      if ( s_axi_wstrb[byte_index] == 1 ) begin
                         sn_req_desc_f_acaddr_3_reg[(byte_index*8) +: 8] <= s_axi_wdata[(byte_index*8) +: 8];
                      end
		  
		  

                endcase // case (axi_awaddr[16:0])
             end // if (reg_wr_en)
           else
             for (i = 0; i < 32 ; i = i + 1) begin


                if (intr_c2h_toggle_clear_0_reg_clear[i])begin
                   intr_c2h_toggle_clear_0_reg[i] <= 1'h0;
                end
                if (intr_c2h_toggle_clear_1_reg_clear[i])begin
                   intr_c2h_toggle_clear_1_reg[i] <= 1'h0;
                end
                if (intr_error_clear_reg_clear[i])begin
                   intr_error_clear_reg[i] <= 1'h0;
                end
                if (rd_req_free_desc_reg_clear[i])begin
                   rd_req_free_desc_reg[i] <= 1'h0;
                end
                if (rd_resp_fifo_push_desc_reg_clear[i])begin
                   rd_resp_fifo_push_desc_reg[i] <= 1'h0;
                end
                if (rd_resp_intr_comp_clear_reg_clear[i])begin
                   rd_resp_intr_comp_clear_reg[i] <= 1'h0;
                end
                if (wr_req_free_desc_reg_clear[i])begin
                   wr_req_free_desc_reg[i] <= 1'h0;
                end
                if (wr_resp_fifo_push_desc_reg_clear[i])begin
                   wr_resp_fifo_push_desc_reg[i] <= 1'h0;
                end
                if (wr_resp_intr_comp_clear_reg_clear[i])begin
                   wr_resp_intr_comp_clear_reg[i] <= 1'h0;
                end
                if (sn_req_fifo_push_desc_reg_clear[i])begin
                   sn_req_fifo_push_desc_reg[i] <= 1'h0;
                end
                if (sn_req_intr_comp_clear_reg_clear[i])begin
                   sn_req_intr_comp_clear_reg[i] <= 1'h0;
                end
                if (sn_resp_free_desc_reg_clear[i])begin
                   sn_resp_free_desc_reg[i] <= 1'h0;
                end
                if (sn_data_free_desc_reg_clear[i])begin
                   sn_data_free_desc_reg[i] <= 1'h0;
                end


             end
           
        end // else: !if( ~rst_n)
     end // always @ ( posedge clk )




   // Implement write response logic generation
   // The write response and response valid signals are asserted by the slave 
   // when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
   // This marks the acceptance of address and indicates the status of 
   // write transaction.

   always @( posedge clk )
     begin
        if ( resetn == 1'b0 )
          begin
             axi_bvalid  <= 0;
             axi_bresp   <= 2'b0;
          end 
        else
          begin    
             if (axi_awready && s_axi_awvalid && ~axi_bvalid && axi_wready && s_axi_wvalid)
               begin
                  // indicates a valid write response is available
                  axi_bvalid <= 1'b1;
                  axi_bresp  <= 2'b0; // 'OKAY' response 
               end                   // work error responses in future
             else
               begin
                  if (s_axi_bready && axi_bvalid) 
                    //check if bready is asserted while bvalid is high) 
                    //(there is a possibility that bready is always asserted high)   
                    axi_bvalid <= 1'b0; 
               end // else: !if(axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
          end // else: !if( S_AXI_ARESETN == 1'b0 )
     end // always @ ( posedge clk )
   
   


   // Implement axi_arready generation
   // axi_arready is asserted for one S_AXI_ACLK clock cycle when
   // S_AXI_ARVALID is asserted. axi_awready is 
   // de-asserted when reset (active low) is asserted. 
   // The read address is also latched when S_AXI_ARVALID is 
   // asserted. axi_araddr is reset to zero on reset assertion.

   always @( posedge clk )
     begin
        if ( resetn == 1'b0 )
          begin
             axi_araddr  <= {S_AXI_ADDR_WIDTH{1'b0}};
          end 
        else
          begin    
             if (~axi_arready && s_axi_arvalid)
               begin
                  // read address latching
                  axi_araddr  <= s_axi_araddr;
               end
             else
               begin
                  axi_araddr  <= axi_araddr;
               end
          end 
     end       


   //

   wire arvalid_pending_pulse;
   reg  arvalid_pending_0;
   reg  arvalid_pending_1 ;
   reg  arvalid_reg;
   
   always@(posedge clk)
     begin
	if ( resetn == 1'b0 )
	  begin
             arvalid_reg <= 1'b0;
             arvalid_pending_0 <= 1'b0;
             arvalid_pending_1 <= 1'b0;
	  end 
	else
	  begin
             arvalid_reg <= s_axi_arvalid;
             arvalid_pending_0 <= ~axi_arready && s_axi_arvalid;
             arvalid_pending_1 <= arvalid_pending_0;
	  end
     end // always@ (posedge clk)
   
   
   assign arvalid_pending_pulse = (arvalid_pending_0 & ~arvalid_pending_1);
   //
   
   
   always @( posedge clk )
     begin
        if ( resetn == 1'b0 )
          begin
             axi_arready <= 1'b0;
          end 
        else
          begin    
             if (~axi_arready)begin
                if (arvalid_pending_0) begin
                   if (~axi_araddr[BRIDGE_MSB] && axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2])begin    // read is targeted to WDATA RAM
                      axi_arready <= wdata_ram_data_ready_2;
                   end
                   else begin
                      if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && ~axi_araddr[BRIDGE_MSB-2])begin    // read is targeted to WSTRB RAM
                         axi_arready <= wstrb_ram_data_ready_2;
                      end
                      //else if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && ~axi_araddr[BRIDGE_MSB-2])begin    // read is targeted to CDDATA RAM
                      else if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2] && ~(|axi_araddr[BRIDGE_MSB-3:BRIDGE_MSB-6])) begin    // read is targeted to CDDATA RAM
                         axi_arready <= cddata_ram_data_ready_2;
                      end
                      else begin    // read is targeted to regs
			 //                           axi_arready <= 1'b1;     // indicates that the slave has acceped the valid read address
                         axi_arready <= arvalid_pending_1;     // indicates that the slave has acceped the valid read address
                      end
                   end
                end
                else 
                  axi_arready <= 1'b0;
             end
             else
               axi_arready <= 1'b0;
          end
     end // always @ ( posedge clk )
   

   
   // Implement memory mapped register select and read logic generation
   // Slave register read enable is asserted when valid address is available
   // and the slave is ready to accept the read address.
   assign reg_rd_en = axi_arready & s_axi_arvalid & ~axi_rvalid;


   reg [S_AXI_DATA_WIDTH-1:0]             reg_data_out_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_1;

   reg 					  reg_block_hit_0;
   reg 					  reg_block_hit_1;
   

   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_1;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_2;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_3;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_4;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_5;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_6;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_7;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_8;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_9;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_a;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_b;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_c;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_d;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_e;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_req_desc_f;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_1;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_2;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_3;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_4;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_5;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_6;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_7;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_8;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_9;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_a;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_b;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_c;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_d;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_e;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_rd_resp_desc_f;
   
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_1;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_2;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_3;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_4;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_5;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_6;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_7;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_8;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_9;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_a;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_b;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_c;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_d;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_e;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_req_desc_f;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_1;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_2;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_3;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_4;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_5;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_6;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_7;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_8;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_9;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_a;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_b;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_c;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_d;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_e;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_wr_resp_desc_f;

   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_1;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_2;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_3;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_4;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_5;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_6;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_7;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_8;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_9;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_a;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_b;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_c;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_d;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_e;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_req_desc_f;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_0;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_1;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_2;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_3;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_4;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_5;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_6;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_7;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_8;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_9;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_a;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_b;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_c;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_d;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_e;
   reg [S_AXI_DATA_WIDTH-1:0] 		  reg_data_out_sn_resp_desc_f;

   reg [15:0] 				  reg_block_hit_rd_req_desc;  //width = XX_MAX_DESC 
   reg [15:0] 				  reg_block_hit_rd_resp_desc; //width = XX_MAX_DESC   
   reg [15:0] 				  reg_block_hit_wr_req_desc;  //width = XX_MAX_DESC 
   reg [15:0] 				  reg_block_hit_wr_resp_desc; //width = XX_MAX_DESC  
   reg [15:0] 				  reg_block_hit_sn_req_desc;  //width = SN_MAX_DESC 
   reg [15:0] 				  reg_block_hit_sn_resp_desc; //width = SN_MAX_DESC  


   always @( posedge clk ) begin

      if (~resetn) begin
         reg_block_hit_rd_req_desc <= 'b0;
      end else begin
         
         if (~|axi_araddr[BRIDGE_MSB:16] && (axi_araddr[15:12]==4'h3) ) begin //access to rd-req-desc reg block   (16 descriptors)
            for (i=0; i<=15; i=i+1) begin : for_reg_block_hit_rd_req_desc
               if(i==axi_araddr[11:8]) begin
                  reg_block_hit_rd_req_desc[i] <= 'b1;
               end else begin
                  reg_block_hit_rd_req_desc[i] <= 'b0;
               end
            end
         end else begin
            reg_block_hit_rd_req_desc <= 'b0;
         end

      end

   end
   
   always @( posedge clk ) begin

      if (~resetn) begin
         reg_block_hit_rd_resp_desc <= 'b0;
      end else begin
         
         if (~|axi_araddr[BRIDGE_MSB:16] && (axi_araddr[15:12]==4'h4) ) begin //access to rd-resp-desc reg block   (16 descriptors)
            for (i=0; i<=15; i=i+1) begin : for_reg_block_hit_rd_resp_desc
               if(i==axi_araddr[11:8]) begin
                  reg_block_hit_rd_resp_desc[i] <= 'b1;
               end else begin
                  reg_block_hit_rd_resp_desc[i] <= 'b0;
               end
            end
         end else begin
            reg_block_hit_rd_resp_desc <= 'b0;
         end

      end

   end
   
   always @( posedge clk ) begin

      if (~resetn) begin
         reg_block_hit_wr_req_desc <= 'b0;
      end else begin
         
         if (~|axi_araddr[BRIDGE_MSB:16] && (axi_araddr[15:12]==4'h5) ) begin //access to wr-req-desc reg block   (16 descriptors)
            for (i=0; i<=15; i=i+1) begin : for_reg_block_hit_wr_req_desc
               if(i==axi_araddr[11:8]) begin
                  reg_block_hit_wr_req_desc[i] <= 'b1;
               end else begin
                  reg_block_hit_wr_req_desc[i] <= 'b0;
               end
            end
         end else begin
            reg_block_hit_wr_req_desc <= 'b0;
         end

      end

   end
   
   always @( posedge clk ) begin

      if (~resetn) begin
         reg_block_hit_wr_resp_desc <= 'b0;
      end else begin
         
         if (~|axi_araddr[BRIDGE_MSB:16] && (axi_araddr[15:12]==4'h6) ) begin //access to wr-resp-desc reg block   (16 descriptors)
            for (i=0; i<=15; i=i+1) begin : for_reg_block_hit_wr_resp_desc
               if(i==axi_araddr[11:8]) begin
                  reg_block_hit_wr_resp_desc[i] <= 'b1;
               end else begin
                  reg_block_hit_wr_resp_desc[i] <= 'b0;
               end
            end
         end else begin
            reg_block_hit_wr_resp_desc <= 'b0;
         end

      end

   end
   
   always @( posedge clk ) begin

      if (~resetn) begin
         reg_block_hit_sn_req_desc <= 'b0;
      end else begin
         
         if (~|axi_araddr[BRIDGE_MSB:16] && (axi_araddr[15:12]==4'h7) && (axi_araddr[11:9]==4'h0) ) begin //access to sn-req-desc reg block   (16 descriptors)
            for (i=0; i<=15; i=i+1) begin : for_reg_block_hit_sn_req_desc
               if((2*i)==axi_araddr[8:4]) begin
                  reg_block_hit_sn_req_desc[i] <= 'b1;
               end else begin
                  reg_block_hit_sn_req_desc[i] <= 'b0;
               end
            end
         end else begin
            reg_block_hit_sn_req_desc <= 'b0;
         end

      end

   end
   
   always @( posedge clk ) begin

      if (~resetn) begin
         reg_block_hit_sn_resp_desc <= 'b0;
      end else begin
         
         if (~|axi_araddr[BRIDGE_MSB:16] && (axi_araddr[15:12]==4'h7) && (axi_araddr[11:9]==4'h1) ) begin //access to sn-req-desc reg block   (16 descriptors)
            for (i=0; i<=15; i=i+1) begin : for_reg_block_hit_sn_resp_desc
               if((2*i)==axi_araddr[8:4]) begin
                  reg_block_hit_sn_resp_desc[i] <= 'b1;
               end else begin
                  reg_block_hit_sn_resp_desc[i] <= 'b0;
               end
            end
         end else begin
            reg_block_hit_sn_resp_desc <= 'b0;
         end

      end

   end
   
   

   always @( posedge clk )
     begin
	if (~resetn)
          begin
             reg_block_hit_0 <= 1'b0;
          end
	else
          begin
             if ( (~|axi_araddr[BRIDGE_MSB:10]) && (~&axi_araddr[9:8]) ) //access to reg block 0
               begin
                  reg_block_hit_0 <= 1'b1;                 

               end
             else
               begin
                  reg_block_hit_0 <= 1'b0;
               end
          end
     end


   always @( posedge clk )
     begin
	if (~resetn)
          begin
             reg_block_hit_1 <= 1'b0;
          end
	else
          begin
             if ( (~|axi_araddr[BRIDGE_MSB:10]) && (&axi_araddr[9:8]) ) //access to reg block 1
               begin
                  reg_block_hit_1 <= 1'b1;                 

               end
             else
               begin
                  reg_block_hit_1 <= 1'b0;
               end
          end
     end



   always @( posedge clk )
     begin
	if (~resetn)
          begin
             reg_data_out_0 <= 32'b0;
          end
	else
          begin

             case ({7'b0000000,axi_araddr[9:0]}) 
               
               //Register reads expect desc
               
               `BRIDGE_IDENTIFICATION_REG_ADDR : reg_data_out_0 <= bridge_identification_reg;
               `LAST_BRIDGE_REG_ADDR : reg_data_out_0 <= last_bridge_reg;
               `VERSION_REG_ADDR : reg_data_out_0 <= version_reg;
               `BRIDGE_TYPE_REG_ADDR : reg_data_out_0 <= bridge_type_reg;
               `MODE_SELECT_REG_ADDR : reg_data_out_0 <= mode_select_reg;
               `RESET_REG_ADDR : reg_data_out_0 <= reset_reg;
               `H2C_INTR_0_REG_ADDR : reg_data_out_0 <= h2c_intr_0_reg;
               `H2C_INTR_1_REG_ADDR : reg_data_out_0 <= h2c_intr_1_reg;
               `H2C_INTR_2_REG_ADDR : reg_data_out_0 <= h2c_intr_2_reg;
               `H2C_INTR_3_REG_ADDR : reg_data_out_0 <= h2c_intr_3_reg;
               `C2H_INTR_STATUS_0_REG_ADDR : reg_data_out_0 <= c2h_intr_status_0_reg;
               `INTR_C2H_TOGGLE_STATUS_0_REG_ADDR : reg_data_out_0 <= intr_c2h_toggle_status_0_reg;
               `INTR_C2H_TOGGLE_CLEAR_0_REG_ADDR : reg_data_out_0 <= intr_c2h_toggle_clear_0_reg;
               `INTR_C2H_TOGGLE_ENABLE_0_REG_ADDR : reg_data_out_0 <= intr_c2h_toggle_enable_0_reg;
               `C2H_INTR_STATUS_1_REG_ADDR : reg_data_out_0 <= c2h_intr_status_1_reg;
               `INTR_C2H_TOGGLE_STATUS_1_REG_ADDR : reg_data_out_0 <= intr_c2h_toggle_status_1_reg;
               `INTR_C2H_TOGGLE_CLEAR_1_REG_ADDR : reg_data_out_0 <= intr_c2h_toggle_clear_1_reg;
               `INTR_C2H_TOGGLE_ENABLE_1_REG_ADDR : reg_data_out_0 <= intr_c2h_toggle_enable_1_reg;
               `C2H_GPIO_0_REG_ADDR : reg_data_out_0 <= c2h_gpio_0_reg;
               `C2H_GPIO_1_REG_ADDR : reg_data_out_0 <= c2h_gpio_1_reg;
               `C2H_GPIO_2_REG_ADDR : reg_data_out_0 <= c2h_gpio_2_reg;
               `C2H_GPIO_3_REG_ADDR : reg_data_out_0 <= c2h_gpio_3_reg;
               `C2H_GPIO_4_REG_ADDR : reg_data_out_0 <= c2h_gpio_4_reg;
               `C2H_GPIO_5_REG_ADDR : reg_data_out_0 <= c2h_gpio_5_reg;
               `C2H_GPIO_6_REG_ADDR : reg_data_out_0 <= c2h_gpio_6_reg;
               `C2H_GPIO_7_REG_ADDR : reg_data_out_0 <= c2h_gpio_7_reg;
               `C2H_GPIO_8_REG_ADDR : reg_data_out_0 <= c2h_gpio_8_reg;
               `C2H_GPIO_9_REG_ADDR : reg_data_out_0 <= c2h_gpio_9_reg;
               `C2H_GPIO_10_REG_ADDR : reg_data_out_0 <= c2h_gpio_10_reg;
               `C2H_GPIO_11_REG_ADDR : reg_data_out_0 <= c2h_gpio_11_reg;
               `C2H_GPIO_12_REG_ADDR : reg_data_out_0 <= c2h_gpio_12_reg;
               `C2H_GPIO_13_REG_ADDR : reg_data_out_0 <= c2h_gpio_13_reg;
               `C2H_GPIO_14_REG_ADDR : reg_data_out_0 <= c2h_gpio_14_reg;
               `C2H_GPIO_15_REG_ADDR : reg_data_out_0 <= c2h_gpio_15_reg;
               `H2C_GPIO_0_REG_ADDR : reg_data_out_0 <= h2c_gpio_0_reg;
               `H2C_GPIO_1_REG_ADDR : reg_data_out_0 <= h2c_gpio_1_reg;
               `H2C_GPIO_2_REG_ADDR : reg_data_out_0 <= h2c_gpio_2_reg;
               `H2C_GPIO_3_REG_ADDR : reg_data_out_0 <= h2c_gpio_3_reg;
               `H2C_GPIO_4_REG_ADDR : reg_data_out_0 <= h2c_gpio_4_reg;
               `H2C_GPIO_5_REG_ADDR : reg_data_out_0 <= h2c_gpio_5_reg;
               `H2C_GPIO_6_REG_ADDR : reg_data_out_0 <= h2c_gpio_6_reg;
               `H2C_GPIO_7_REG_ADDR : reg_data_out_0 <= h2c_gpio_7_reg;
               `H2C_GPIO_8_REG_ADDR : reg_data_out_0 <= h2c_gpio_8_reg;
               `H2C_GPIO_9_REG_ADDR : reg_data_out_0 <= h2c_gpio_9_reg;
               `H2C_GPIO_10_REG_ADDR : reg_data_out_0 <= h2c_gpio_10_reg;
               `H2C_GPIO_11_REG_ADDR : reg_data_out_0 <= h2c_gpio_11_reg;
               `H2C_GPIO_12_REG_ADDR : reg_data_out_0 <= h2c_gpio_12_reg;
               `H2C_GPIO_13_REG_ADDR : reg_data_out_0 <= h2c_gpio_13_reg;
               `H2C_GPIO_14_REG_ADDR : reg_data_out_0 <= h2c_gpio_14_reg;
               `H2C_GPIO_15_REG_ADDR : reg_data_out_0 <= h2c_gpio_15_reg;
               `BRIDGE_CONFIG_REG_ADDR : reg_data_out_0 <= bridge_config_reg;
               `INTR_STATUS_REG_ADDR : reg_data_out_0 <= intr_status_reg;
               `INTR_ERROR_STATUS_REG_ADDR : reg_data_out_0 <= intr_error_status_reg;
               `INTR_ERROR_CLEAR_REG_ADDR : reg_data_out_0 <= intr_error_clear_reg;
               `INTR_ERROR_ENABLE_REG_ADDR : reg_data_out_0 <= intr_error_enable_reg;
               `BRIDGE_RD_USER_CONFIG_REG_ADDR : reg_data_out_0 <= bridge_rd_user_config_reg;
               `BRIDGE_WR_USER_CONFIG_REG_ADDR : reg_data_out_0 <= bridge_wr_user_config_reg;
               `RD_MAX_DESC_REG_ADDR : reg_data_out_0 <= rd_max_desc_reg;
               `WR_MAX_DESC_REG_ADDR : reg_data_out_0 <= wr_max_desc_reg;
               `SN_MAX_DESC_REG_ADDR : reg_data_out_0 <= sn_max_desc_reg;
               
               default                                  :reg_data_out_0 <= 32'b0      ;        
             endcase
          end
     end


   always @( posedge clk )
     begin
	if (~resetn)
          begin
             reg_data_out_1 <= 32'b0;
          end
	else
          begin

             case ({9'b000000011,axi_araddr[7:0]}) 
               
               //Register reads expect desc
               
               `RD_REQ_FREE_DESC_REG_ADDR : reg_data_out_1 <= rd_req_free_desc_reg;
               `RD_REQ_FIFO_POP_DESC_REG_ADDR : reg_data_out_1 <= rd_req_fifo_pop_desc_reg;
               `RD_REQ_FIFO_FILL_LEVEL_REG_ADDR : reg_data_out_1 <= rd_req_fifo_fill_level_reg;
               `RD_RESP_FIFO_PUSH_DESC_REG_ADDR : reg_data_out_1 <= rd_resp_fifo_push_desc_reg;
               `RD_RESP_FIFO_FREE_LEVEL_REG_ADDR : reg_data_out_1 <= rd_resp_fifo_free_level_reg;
               `RD_RESP_INTR_COMP_STATUS_REG_ADDR : reg_data_out_1 <= rd_resp_intr_comp_status_reg;
               `RD_RESP_INTR_COMP_CLEAR_REG_ADDR : reg_data_out_1 <= rd_resp_intr_comp_clear_reg;
               `RD_RESP_INTR_COMP_ENABLE_REG_ADDR : reg_data_out_1 <= rd_resp_intr_comp_enable_reg;
               `WR_REQ_FREE_DESC_REG_ADDR : reg_data_out_1 <= wr_req_free_desc_reg;
               `WR_REQ_FIFO_POP_DESC_REG_ADDR : reg_data_out_1 <= wr_req_fifo_pop_desc_reg;
               `WR_REQ_FIFO_FILL_LEVEL_REG_ADDR : reg_data_out_1 <= wr_req_fifo_fill_level_reg;
               `WR_RESP_FIFO_PUSH_DESC_REG_ADDR : reg_data_out_1 <= wr_resp_fifo_push_desc_reg;
               `WR_RESP_FIFO_FREE_LEVEL_REG_ADDR : reg_data_out_1 <= wr_resp_fifo_free_level_reg;
               `WR_RESP_INTR_COMP_STATUS_REG_ADDR : reg_data_out_1 <= wr_resp_intr_comp_status_reg;
               `WR_RESP_INTR_COMP_CLEAR_REG_ADDR : reg_data_out_1 <= wr_resp_intr_comp_clear_reg;
               `WR_RESP_INTR_COMP_ENABLE_REG_ADDR : reg_data_out_1 <= wr_resp_intr_comp_enable_reg;
               `SN_REQ_FIFO_PUSH_DESC_REG_ADDR : reg_data_out_1 <= sn_req_fifo_push_desc_reg;
               `SN_REQ_FIFO_FREE_LEVEL_REG_ADDR : reg_data_out_1 <= sn_req_fifo_free_level_reg;
               `SN_REQ_INTR_COMP_STATUS_REG_ADDR : reg_data_out_1 <= sn_req_intr_comp_status_reg;
               `SN_REQ_INTR_COMP_CLEAR_REG_ADDR : reg_data_out_1 <= sn_req_intr_comp_clear_reg;
               `SN_REQ_INTR_COMP_ENABLE_REG_ADDR : reg_data_out_1 <= sn_req_intr_comp_enable_reg;
               `SN_RESP_FREE_DESC_REG_ADDR : reg_data_out_1 <= sn_resp_free_desc_reg;
               `SN_RESP_FIFO_POP_DESC_REG_ADDR : reg_data_out_1 <= sn_resp_fifo_pop_desc_reg;
               `SN_RESP_FIFO_FILL_LEVEL_REG_ADDR : reg_data_out_1 <= sn_resp_fifo_fill_level_reg;
               `SN_DATA_FREE_DESC_REG_ADDR : reg_data_out_1 <= sn_data_free_desc_reg;
               `SN_DATA_FIFO_POP_DESC_REG_ADDR : reg_data_out_1 <= sn_data_fifo_pop_desc_reg;
               `SN_DATA_FIFO_FILL_LEVEL_REG_ADDR : reg_data_out_1 <= sn_data_fifo_fill_level_reg;
               `INTR_FIFO_ENABLE_REG_ADDR : reg_data_out_1 <= intr_fifo_enable_reg;
               
               
               default                                  :reg_data_out_1 <= 32'b0      ;        
             endcase
          end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_0 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_0_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_txn_type_reg;
               (`RD_REQ_DESC_0_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_size_reg;
               (`RD_REQ_DESC_0_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axsize_reg;
               (`RD_REQ_DESC_0_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_attr_reg;
               (`RD_REQ_DESC_0_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axaddr_0_reg;
               (`RD_REQ_DESC_0_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axaddr_1_reg;
               (`RD_REQ_DESC_0_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axaddr_2_reg;
               (`RD_REQ_DESC_0_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axaddr_3_reg;
               (`RD_REQ_DESC_0_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axid_0_reg;
               (`RD_REQ_DESC_0_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axid_1_reg;
               (`RD_REQ_DESC_0_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axid_2_reg;
               (`RD_REQ_DESC_0_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axid_3_reg;
               (`RD_REQ_DESC_0_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_0_reg;
               (`RD_REQ_DESC_0_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_1_reg;
               (`RD_REQ_DESC_0_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_2_reg;
               (`RD_REQ_DESC_0_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_3_reg;
               (`RD_REQ_DESC_0_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_4_reg;
               (`RD_REQ_DESC_0_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_5_reg;
               (`RD_REQ_DESC_0_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_6_reg;
               (`RD_REQ_DESC_0_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_7_reg;
               (`RD_REQ_DESC_0_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_8_reg;
               (`RD_REQ_DESC_0_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_9_reg;
               (`RD_REQ_DESC_0_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_10_reg;
               (`RD_REQ_DESC_0_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_11_reg;
               (`RD_REQ_DESC_0_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_12_reg;
               (`RD_REQ_DESC_0_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_13_reg;
               (`RD_REQ_DESC_0_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_14_reg;
               (`RD_REQ_DESC_0_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_0 <= rd_req_desc_0_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_0 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_1 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_1_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_txn_type_reg;
               (`RD_REQ_DESC_1_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_size_reg;
               (`RD_REQ_DESC_1_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axsize_reg;
               (`RD_REQ_DESC_1_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_attr_reg;
               (`RD_REQ_DESC_1_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axaddr_0_reg;
               (`RD_REQ_DESC_1_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axaddr_1_reg;
               (`RD_REQ_DESC_1_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axaddr_2_reg;
               (`RD_REQ_DESC_1_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axaddr_3_reg;
               (`RD_REQ_DESC_1_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axid_0_reg;
               (`RD_REQ_DESC_1_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axid_1_reg;
               (`RD_REQ_DESC_1_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axid_2_reg;
               (`RD_REQ_DESC_1_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axid_3_reg;
               (`RD_REQ_DESC_1_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_0_reg;
               (`RD_REQ_DESC_1_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_1_reg;
               (`RD_REQ_DESC_1_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_2_reg;
               (`RD_REQ_DESC_1_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_3_reg;
               (`RD_REQ_DESC_1_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_4_reg;
               (`RD_REQ_DESC_1_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_5_reg;
               (`RD_REQ_DESC_1_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_6_reg;
               (`RD_REQ_DESC_1_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_7_reg;
               (`RD_REQ_DESC_1_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_8_reg;
               (`RD_REQ_DESC_1_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_9_reg;
               (`RD_REQ_DESC_1_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_10_reg;
               (`RD_REQ_DESC_1_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_11_reg;
               (`RD_REQ_DESC_1_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_12_reg;
               (`RD_REQ_DESC_1_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_13_reg;
               (`RD_REQ_DESC_1_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_14_reg;
               (`RD_REQ_DESC_1_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_1 <= rd_req_desc_1_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_1 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_2 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_2_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_txn_type_reg;
               (`RD_REQ_DESC_2_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_size_reg;
               (`RD_REQ_DESC_2_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axsize_reg;
               (`RD_REQ_DESC_2_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_attr_reg;
               (`RD_REQ_DESC_2_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axaddr_0_reg;
               (`RD_REQ_DESC_2_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axaddr_1_reg;
               (`RD_REQ_DESC_2_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axaddr_2_reg;
               (`RD_REQ_DESC_2_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axaddr_3_reg;
               (`RD_REQ_DESC_2_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axid_0_reg;
               (`RD_REQ_DESC_2_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axid_1_reg;
               (`RD_REQ_DESC_2_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axid_2_reg;
               (`RD_REQ_DESC_2_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axid_3_reg;
               (`RD_REQ_DESC_2_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_0_reg;
               (`RD_REQ_DESC_2_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_1_reg;
               (`RD_REQ_DESC_2_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_2_reg;
               (`RD_REQ_DESC_2_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_3_reg;
               (`RD_REQ_DESC_2_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_4_reg;
               (`RD_REQ_DESC_2_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_5_reg;
               (`RD_REQ_DESC_2_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_6_reg;
               (`RD_REQ_DESC_2_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_7_reg;
               (`RD_REQ_DESC_2_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_8_reg;
               (`RD_REQ_DESC_2_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_9_reg;
               (`RD_REQ_DESC_2_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_10_reg;
               (`RD_REQ_DESC_2_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_11_reg;
               (`RD_REQ_DESC_2_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_12_reg;
               (`RD_REQ_DESC_2_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_13_reg;
               (`RD_REQ_DESC_2_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_14_reg;
               (`RD_REQ_DESC_2_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_2 <= rd_req_desc_2_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_2 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_3 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_3_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_txn_type_reg;
               (`RD_REQ_DESC_3_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_size_reg;
               (`RD_REQ_DESC_3_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axsize_reg;
               (`RD_REQ_DESC_3_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_attr_reg;
               (`RD_REQ_DESC_3_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axaddr_0_reg;
               (`RD_REQ_DESC_3_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axaddr_1_reg;
               (`RD_REQ_DESC_3_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axaddr_2_reg;
               (`RD_REQ_DESC_3_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axaddr_3_reg;
               (`RD_REQ_DESC_3_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axid_0_reg;
               (`RD_REQ_DESC_3_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axid_1_reg;
               (`RD_REQ_DESC_3_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axid_2_reg;
               (`RD_REQ_DESC_3_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axid_3_reg;
               (`RD_REQ_DESC_3_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_0_reg;
               (`RD_REQ_DESC_3_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_1_reg;
               (`RD_REQ_DESC_3_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_2_reg;
               (`RD_REQ_DESC_3_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_3_reg;
               (`RD_REQ_DESC_3_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_4_reg;
               (`RD_REQ_DESC_3_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_5_reg;
               (`RD_REQ_DESC_3_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_6_reg;
               (`RD_REQ_DESC_3_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_7_reg;
               (`RD_REQ_DESC_3_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_8_reg;
               (`RD_REQ_DESC_3_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_9_reg;
               (`RD_REQ_DESC_3_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_10_reg;
               (`RD_REQ_DESC_3_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_11_reg;
               (`RD_REQ_DESC_3_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_12_reg;
               (`RD_REQ_DESC_3_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_13_reg;
               (`RD_REQ_DESC_3_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_14_reg;
               (`RD_REQ_DESC_3_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_3 <= rd_req_desc_3_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_3 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_4 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_4_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_txn_type_reg;
               (`RD_REQ_DESC_4_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_size_reg;
               (`RD_REQ_DESC_4_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axsize_reg;
               (`RD_REQ_DESC_4_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_attr_reg;
               (`RD_REQ_DESC_4_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axaddr_0_reg;
               (`RD_REQ_DESC_4_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axaddr_1_reg;
               (`RD_REQ_DESC_4_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axaddr_2_reg;
               (`RD_REQ_DESC_4_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axaddr_3_reg;
               (`RD_REQ_DESC_4_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axid_0_reg;
               (`RD_REQ_DESC_4_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axid_1_reg;
               (`RD_REQ_DESC_4_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axid_2_reg;
               (`RD_REQ_DESC_4_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axid_3_reg;
               (`RD_REQ_DESC_4_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_0_reg;
               (`RD_REQ_DESC_4_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_1_reg;
               (`RD_REQ_DESC_4_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_2_reg;
               (`RD_REQ_DESC_4_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_3_reg;
               (`RD_REQ_DESC_4_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_4_reg;
               (`RD_REQ_DESC_4_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_5_reg;
               (`RD_REQ_DESC_4_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_6_reg;
               (`RD_REQ_DESC_4_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_7_reg;
               (`RD_REQ_DESC_4_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_8_reg;
               (`RD_REQ_DESC_4_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_9_reg;
               (`RD_REQ_DESC_4_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_10_reg;
               (`RD_REQ_DESC_4_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_11_reg;
               (`RD_REQ_DESC_4_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_12_reg;
               (`RD_REQ_DESC_4_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_13_reg;
               (`RD_REQ_DESC_4_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_14_reg;
               (`RD_REQ_DESC_4_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_4 <= rd_req_desc_4_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_4 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_5 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_5_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_txn_type_reg;
               (`RD_REQ_DESC_5_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_size_reg;
               (`RD_REQ_DESC_5_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axsize_reg;
               (`RD_REQ_DESC_5_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_attr_reg;
               (`RD_REQ_DESC_5_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axaddr_0_reg;
               (`RD_REQ_DESC_5_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axaddr_1_reg;
               (`RD_REQ_DESC_5_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axaddr_2_reg;
               (`RD_REQ_DESC_5_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axaddr_3_reg;
               (`RD_REQ_DESC_5_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axid_0_reg;
               (`RD_REQ_DESC_5_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axid_1_reg;
               (`RD_REQ_DESC_5_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axid_2_reg;
               (`RD_REQ_DESC_5_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axid_3_reg;
               (`RD_REQ_DESC_5_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_0_reg;
               (`RD_REQ_DESC_5_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_1_reg;
               (`RD_REQ_DESC_5_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_2_reg;
               (`RD_REQ_DESC_5_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_3_reg;
               (`RD_REQ_DESC_5_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_4_reg;
               (`RD_REQ_DESC_5_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_5_reg;
               (`RD_REQ_DESC_5_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_6_reg;
               (`RD_REQ_DESC_5_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_7_reg;
               (`RD_REQ_DESC_5_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_8_reg;
               (`RD_REQ_DESC_5_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_9_reg;
               (`RD_REQ_DESC_5_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_10_reg;
               (`RD_REQ_DESC_5_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_11_reg;
               (`RD_REQ_DESC_5_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_12_reg;
               (`RD_REQ_DESC_5_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_13_reg;
               (`RD_REQ_DESC_5_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_14_reg;
               (`RD_REQ_DESC_5_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_5 <= rd_req_desc_5_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_5 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_6 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_6_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_txn_type_reg;
               (`RD_REQ_DESC_6_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_size_reg;
               (`RD_REQ_DESC_6_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axsize_reg;
               (`RD_REQ_DESC_6_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_attr_reg;
               (`RD_REQ_DESC_6_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axaddr_0_reg;
               (`RD_REQ_DESC_6_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axaddr_1_reg;
               (`RD_REQ_DESC_6_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axaddr_2_reg;
               (`RD_REQ_DESC_6_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axaddr_3_reg;
               (`RD_REQ_DESC_6_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axid_0_reg;
               (`RD_REQ_DESC_6_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axid_1_reg;
               (`RD_REQ_DESC_6_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axid_2_reg;
               (`RD_REQ_DESC_6_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axid_3_reg;
               (`RD_REQ_DESC_6_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_0_reg;
               (`RD_REQ_DESC_6_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_1_reg;
               (`RD_REQ_DESC_6_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_2_reg;
               (`RD_REQ_DESC_6_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_3_reg;
               (`RD_REQ_DESC_6_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_4_reg;
               (`RD_REQ_DESC_6_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_5_reg;
               (`RD_REQ_DESC_6_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_6_reg;
               (`RD_REQ_DESC_6_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_7_reg;
               (`RD_REQ_DESC_6_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_8_reg;
               (`RD_REQ_DESC_6_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_9_reg;
               (`RD_REQ_DESC_6_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_10_reg;
               (`RD_REQ_DESC_6_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_11_reg;
               (`RD_REQ_DESC_6_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_12_reg;
               (`RD_REQ_DESC_6_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_13_reg;
               (`RD_REQ_DESC_6_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_14_reg;
               (`RD_REQ_DESC_6_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_6 <= rd_req_desc_6_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_6 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_7 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_7_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_txn_type_reg;
               (`RD_REQ_DESC_7_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_size_reg;
               (`RD_REQ_DESC_7_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axsize_reg;
               (`RD_REQ_DESC_7_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_attr_reg;
               (`RD_REQ_DESC_7_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axaddr_0_reg;
               (`RD_REQ_DESC_7_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axaddr_1_reg;
               (`RD_REQ_DESC_7_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axaddr_2_reg;
               (`RD_REQ_DESC_7_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axaddr_3_reg;
               (`RD_REQ_DESC_7_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axid_0_reg;
               (`RD_REQ_DESC_7_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axid_1_reg;
               (`RD_REQ_DESC_7_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axid_2_reg;
               (`RD_REQ_DESC_7_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axid_3_reg;
               (`RD_REQ_DESC_7_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_0_reg;
               (`RD_REQ_DESC_7_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_1_reg;
               (`RD_REQ_DESC_7_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_2_reg;
               (`RD_REQ_DESC_7_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_3_reg;
               (`RD_REQ_DESC_7_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_4_reg;
               (`RD_REQ_DESC_7_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_5_reg;
               (`RD_REQ_DESC_7_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_6_reg;
               (`RD_REQ_DESC_7_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_7_reg;
               (`RD_REQ_DESC_7_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_8_reg;
               (`RD_REQ_DESC_7_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_9_reg;
               (`RD_REQ_DESC_7_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_10_reg;
               (`RD_REQ_DESC_7_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_11_reg;
               (`RD_REQ_DESC_7_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_12_reg;
               (`RD_REQ_DESC_7_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_13_reg;
               (`RD_REQ_DESC_7_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_14_reg;
               (`RD_REQ_DESC_7_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_7 <= rd_req_desc_7_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_7 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_8 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_8_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_txn_type_reg;
               (`RD_REQ_DESC_8_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_size_reg;
               (`RD_REQ_DESC_8_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axsize_reg;
               (`RD_REQ_DESC_8_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_attr_reg;
               (`RD_REQ_DESC_8_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axaddr_0_reg;
               (`RD_REQ_DESC_8_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axaddr_1_reg;
               (`RD_REQ_DESC_8_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axaddr_2_reg;
               (`RD_REQ_DESC_8_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axaddr_3_reg;
               (`RD_REQ_DESC_8_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axid_0_reg;
               (`RD_REQ_DESC_8_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axid_1_reg;
               (`RD_REQ_DESC_8_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axid_2_reg;
               (`RD_REQ_DESC_8_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axid_3_reg;
               (`RD_REQ_DESC_8_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_0_reg;
               (`RD_REQ_DESC_8_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_1_reg;
               (`RD_REQ_DESC_8_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_2_reg;
               (`RD_REQ_DESC_8_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_3_reg;
               (`RD_REQ_DESC_8_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_4_reg;
               (`RD_REQ_DESC_8_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_5_reg;
               (`RD_REQ_DESC_8_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_6_reg;
               (`RD_REQ_DESC_8_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_7_reg;
               (`RD_REQ_DESC_8_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_8_reg;
               (`RD_REQ_DESC_8_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_9_reg;
               (`RD_REQ_DESC_8_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_10_reg;
               (`RD_REQ_DESC_8_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_11_reg;
               (`RD_REQ_DESC_8_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_12_reg;
               (`RD_REQ_DESC_8_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_13_reg;
               (`RD_REQ_DESC_8_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_14_reg;
               (`RD_REQ_DESC_8_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_8 <= rd_req_desc_8_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_8 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_9 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_9_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_txn_type_reg;
               (`RD_REQ_DESC_9_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_size_reg;
               (`RD_REQ_DESC_9_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axsize_reg;
               (`RD_REQ_DESC_9_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_attr_reg;
               (`RD_REQ_DESC_9_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axaddr_0_reg;
               (`RD_REQ_DESC_9_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axaddr_1_reg;
               (`RD_REQ_DESC_9_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axaddr_2_reg;
               (`RD_REQ_DESC_9_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axaddr_3_reg;
               (`RD_REQ_DESC_9_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axid_0_reg;
               (`RD_REQ_DESC_9_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axid_1_reg;
               (`RD_REQ_DESC_9_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axid_2_reg;
               (`RD_REQ_DESC_9_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axid_3_reg;
               (`RD_REQ_DESC_9_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_0_reg;
               (`RD_REQ_DESC_9_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_1_reg;
               (`RD_REQ_DESC_9_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_2_reg;
               (`RD_REQ_DESC_9_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_3_reg;
               (`RD_REQ_DESC_9_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_4_reg;
               (`RD_REQ_DESC_9_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_5_reg;
               (`RD_REQ_DESC_9_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_6_reg;
               (`RD_REQ_DESC_9_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_7_reg;
               (`RD_REQ_DESC_9_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_8_reg;
               (`RD_REQ_DESC_9_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_9_reg;
               (`RD_REQ_DESC_9_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_10_reg;
               (`RD_REQ_DESC_9_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_11_reg;
               (`RD_REQ_DESC_9_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_12_reg;
               (`RD_REQ_DESC_9_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_13_reg;
               (`RD_REQ_DESC_9_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_14_reg;
               (`RD_REQ_DESC_9_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_9 <= rd_req_desc_9_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_9 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_a <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_A_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_txn_type_reg;
               (`RD_REQ_DESC_A_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_size_reg;
               (`RD_REQ_DESC_A_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axsize_reg;
               (`RD_REQ_DESC_A_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_attr_reg;
               (`RD_REQ_DESC_A_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axaddr_0_reg;
               (`RD_REQ_DESC_A_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axaddr_1_reg;
               (`RD_REQ_DESC_A_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axaddr_2_reg;
               (`RD_REQ_DESC_A_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axaddr_3_reg;
               (`RD_REQ_DESC_A_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axid_0_reg;
               (`RD_REQ_DESC_A_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axid_1_reg;
               (`RD_REQ_DESC_A_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axid_2_reg;
               (`RD_REQ_DESC_A_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axid_3_reg;
               (`RD_REQ_DESC_A_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_0_reg;
               (`RD_REQ_DESC_A_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_1_reg;
               (`RD_REQ_DESC_A_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_2_reg;
               (`RD_REQ_DESC_A_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_3_reg;
               (`RD_REQ_DESC_A_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_4_reg;
               (`RD_REQ_DESC_A_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_5_reg;
               (`RD_REQ_DESC_A_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_6_reg;
               (`RD_REQ_DESC_A_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_7_reg;
               (`RD_REQ_DESC_A_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_8_reg;
               (`RD_REQ_DESC_A_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_9_reg;
               (`RD_REQ_DESC_A_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_10_reg;
               (`RD_REQ_DESC_A_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_11_reg;
               (`RD_REQ_DESC_A_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_12_reg;
               (`RD_REQ_DESC_A_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_13_reg;
               (`RD_REQ_DESC_A_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_14_reg;
               (`RD_REQ_DESC_A_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_a <= rd_req_desc_a_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_a <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_b <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_B_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_txn_type_reg;
               (`RD_REQ_DESC_B_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_size_reg;
               (`RD_REQ_DESC_B_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axsize_reg;
               (`RD_REQ_DESC_B_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_attr_reg;
               (`RD_REQ_DESC_B_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axaddr_0_reg;
               (`RD_REQ_DESC_B_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axaddr_1_reg;
               (`RD_REQ_DESC_B_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axaddr_2_reg;
               (`RD_REQ_DESC_B_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axaddr_3_reg;
               (`RD_REQ_DESC_B_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axid_0_reg;
               (`RD_REQ_DESC_B_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axid_1_reg;
               (`RD_REQ_DESC_B_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axid_2_reg;
               (`RD_REQ_DESC_B_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axid_3_reg;
               (`RD_REQ_DESC_B_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_0_reg;
               (`RD_REQ_DESC_B_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_1_reg;
               (`RD_REQ_DESC_B_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_2_reg;
               (`RD_REQ_DESC_B_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_3_reg;
               (`RD_REQ_DESC_B_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_4_reg;
               (`RD_REQ_DESC_B_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_5_reg;
               (`RD_REQ_DESC_B_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_6_reg;
               (`RD_REQ_DESC_B_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_7_reg;
               (`RD_REQ_DESC_B_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_8_reg;
               (`RD_REQ_DESC_B_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_9_reg;
               (`RD_REQ_DESC_B_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_10_reg;
               (`RD_REQ_DESC_B_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_11_reg;
               (`RD_REQ_DESC_B_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_12_reg;
               (`RD_REQ_DESC_B_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_13_reg;
               (`RD_REQ_DESC_B_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_14_reg;
               (`RD_REQ_DESC_B_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_b <= rd_req_desc_b_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_b <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_c <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_C_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_txn_type_reg;
               (`RD_REQ_DESC_C_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_size_reg;
               (`RD_REQ_DESC_C_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axsize_reg;
               (`RD_REQ_DESC_C_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_attr_reg;
               (`RD_REQ_DESC_C_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axaddr_0_reg;
               (`RD_REQ_DESC_C_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axaddr_1_reg;
               (`RD_REQ_DESC_C_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axaddr_2_reg;
               (`RD_REQ_DESC_C_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axaddr_3_reg;
               (`RD_REQ_DESC_C_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axid_0_reg;
               (`RD_REQ_DESC_C_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axid_1_reg;
               (`RD_REQ_DESC_C_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axid_2_reg;
               (`RD_REQ_DESC_C_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axid_3_reg;
               (`RD_REQ_DESC_C_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_0_reg;
               (`RD_REQ_DESC_C_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_1_reg;
               (`RD_REQ_DESC_C_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_2_reg;
               (`RD_REQ_DESC_C_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_3_reg;
               (`RD_REQ_DESC_C_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_4_reg;
               (`RD_REQ_DESC_C_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_5_reg;
               (`RD_REQ_DESC_C_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_6_reg;
               (`RD_REQ_DESC_C_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_7_reg;
               (`RD_REQ_DESC_C_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_8_reg;
               (`RD_REQ_DESC_C_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_9_reg;
               (`RD_REQ_DESC_C_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_10_reg;
               (`RD_REQ_DESC_C_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_11_reg;
               (`RD_REQ_DESC_C_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_12_reg;
               (`RD_REQ_DESC_C_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_13_reg;
               (`RD_REQ_DESC_C_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_14_reg;
               (`RD_REQ_DESC_C_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_c <= rd_req_desc_c_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_c <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_d <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_D_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_txn_type_reg;
               (`RD_REQ_DESC_D_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_size_reg;
               (`RD_REQ_DESC_D_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axsize_reg;
               (`RD_REQ_DESC_D_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_attr_reg;
               (`RD_REQ_DESC_D_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axaddr_0_reg;
               (`RD_REQ_DESC_D_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axaddr_1_reg;
               (`RD_REQ_DESC_D_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axaddr_2_reg;
               (`RD_REQ_DESC_D_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axaddr_3_reg;
               (`RD_REQ_DESC_D_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axid_0_reg;
               (`RD_REQ_DESC_D_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axid_1_reg;
               (`RD_REQ_DESC_D_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axid_2_reg;
               (`RD_REQ_DESC_D_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axid_3_reg;
               (`RD_REQ_DESC_D_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_0_reg;
               (`RD_REQ_DESC_D_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_1_reg;
               (`RD_REQ_DESC_D_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_2_reg;
               (`RD_REQ_DESC_D_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_3_reg;
               (`RD_REQ_DESC_D_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_4_reg;
               (`RD_REQ_DESC_D_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_5_reg;
               (`RD_REQ_DESC_D_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_6_reg;
               (`RD_REQ_DESC_D_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_7_reg;
               (`RD_REQ_DESC_D_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_8_reg;
               (`RD_REQ_DESC_D_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_9_reg;
               (`RD_REQ_DESC_D_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_10_reg;
               (`RD_REQ_DESC_D_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_11_reg;
               (`RD_REQ_DESC_D_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_12_reg;
               (`RD_REQ_DESC_D_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_13_reg;
               (`RD_REQ_DESC_D_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_14_reg;
               (`RD_REQ_DESC_D_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_d <= rd_req_desc_d_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_d <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_e <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_E_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_txn_type_reg;
               (`RD_REQ_DESC_E_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_size_reg;
               (`RD_REQ_DESC_E_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axsize_reg;
               (`RD_REQ_DESC_E_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_attr_reg;
               (`RD_REQ_DESC_E_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axaddr_0_reg;
               (`RD_REQ_DESC_E_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axaddr_1_reg;
               (`RD_REQ_DESC_E_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axaddr_2_reg;
               (`RD_REQ_DESC_E_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axaddr_3_reg;
               (`RD_REQ_DESC_E_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axid_0_reg;
               (`RD_REQ_DESC_E_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axid_1_reg;
               (`RD_REQ_DESC_E_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axid_2_reg;
               (`RD_REQ_DESC_E_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axid_3_reg;
               (`RD_REQ_DESC_E_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_0_reg;
               (`RD_REQ_DESC_E_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_1_reg;
               (`RD_REQ_DESC_E_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_2_reg;
               (`RD_REQ_DESC_E_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_3_reg;
               (`RD_REQ_DESC_E_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_4_reg;
               (`RD_REQ_DESC_E_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_5_reg;
               (`RD_REQ_DESC_E_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_6_reg;
               (`RD_REQ_DESC_E_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_7_reg;
               (`RD_REQ_DESC_E_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_8_reg;
               (`RD_REQ_DESC_E_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_9_reg;
               (`RD_REQ_DESC_E_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_10_reg;
               (`RD_REQ_DESC_E_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_11_reg;
               (`RD_REQ_DESC_E_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_12_reg;
               (`RD_REQ_DESC_E_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_13_reg;
               (`RD_REQ_DESC_E_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_14_reg;
               (`RD_REQ_DESC_E_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_e <= rd_req_desc_e_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_e <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_req_desc_f <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_REQ_DESC_F_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_txn_type_reg;
               (`RD_REQ_DESC_F_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_size_reg;
               (`RD_REQ_DESC_F_AXSIZE_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axsize_reg;
               (`RD_REQ_DESC_F_ATTR_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_attr_reg;
               (`RD_REQ_DESC_F_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axaddr_0_reg;
               (`RD_REQ_DESC_F_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axaddr_1_reg;
               (`RD_REQ_DESC_F_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axaddr_2_reg;
               (`RD_REQ_DESC_F_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axaddr_3_reg;
               (`RD_REQ_DESC_F_AXID_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axid_0_reg;
               (`RD_REQ_DESC_F_AXID_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axid_1_reg;
               (`RD_REQ_DESC_F_AXID_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axid_2_reg;
               (`RD_REQ_DESC_F_AXID_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axid_3_reg;
               (`RD_REQ_DESC_F_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_0_reg;
               (`RD_REQ_DESC_F_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_1_reg;
               (`RD_REQ_DESC_F_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_2_reg;
               (`RD_REQ_DESC_F_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_3_reg;
               (`RD_REQ_DESC_F_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_4_reg;
               (`RD_REQ_DESC_F_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_5_reg;
               (`RD_REQ_DESC_F_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_6_reg;
               (`RD_REQ_DESC_F_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_7_reg;
               (`RD_REQ_DESC_F_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_8_reg;
               (`RD_REQ_DESC_F_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_9_reg;
               (`RD_REQ_DESC_F_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_10_reg;
               (`RD_REQ_DESC_F_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_11_reg;
               (`RD_REQ_DESC_F_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_12_reg;
               (`RD_REQ_DESC_F_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_13_reg;
               (`RD_REQ_DESC_F_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_14_reg;
               (`RD_REQ_DESC_F_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_req_desc_f <= rd_req_desc_f_axuser_15_reg;
               default                                  :reg_data_out_rd_req_desc_f <= 32'b0      ;        
             endcase
	  end
     end




   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_0 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_0_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_data_offset_reg;
               (`RD_RESP_DESC_0_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_data_size_reg;
               (`RD_RESP_DESC_0_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_data_host_addr_0_reg;
               (`RD_RESP_DESC_0_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_data_host_addr_1_reg;
               (`RD_RESP_DESC_0_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_data_host_addr_2_reg;
               (`RD_RESP_DESC_0_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_data_host_addr_3_reg;
               (`RD_RESP_DESC_0_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_resp_reg;
               (`RD_RESP_DESC_0_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xid_0_reg;
               (`RD_RESP_DESC_0_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xid_1_reg;
               (`RD_RESP_DESC_0_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xid_2_reg;
               (`RD_RESP_DESC_0_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xid_3_reg;
               (`RD_RESP_DESC_0_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_0_reg;
               (`RD_RESP_DESC_0_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_1_reg;
               (`RD_RESP_DESC_0_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_2_reg;
               (`RD_RESP_DESC_0_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_3_reg;
               (`RD_RESP_DESC_0_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_4_reg;
               (`RD_RESP_DESC_0_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_5_reg;
               (`RD_RESP_DESC_0_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_6_reg;
               (`RD_RESP_DESC_0_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_7_reg;
               (`RD_RESP_DESC_0_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_8_reg;
               (`RD_RESP_DESC_0_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_9_reg;
               (`RD_RESP_DESC_0_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_10_reg;
               (`RD_RESP_DESC_0_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_11_reg;
               (`RD_RESP_DESC_0_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_12_reg;
               (`RD_RESP_DESC_0_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_13_reg;
               (`RD_RESP_DESC_0_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_14_reg;
               (`RD_RESP_DESC_0_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_0 <= rd_resp_desc_0_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_0 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_1 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_1_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_data_offset_reg;
               (`RD_RESP_DESC_1_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_data_size_reg;
               (`RD_RESP_DESC_1_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_data_host_addr_0_reg;
               (`RD_RESP_DESC_1_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_data_host_addr_1_reg;
               (`RD_RESP_DESC_1_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_data_host_addr_2_reg;
               (`RD_RESP_DESC_1_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_data_host_addr_3_reg;
               (`RD_RESP_DESC_1_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_resp_reg;
               (`RD_RESP_DESC_1_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xid_0_reg;
               (`RD_RESP_DESC_1_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xid_1_reg;
               (`RD_RESP_DESC_1_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xid_2_reg;
               (`RD_RESP_DESC_1_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xid_3_reg;
               (`RD_RESP_DESC_1_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_0_reg;
               (`RD_RESP_DESC_1_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_1_reg;
               (`RD_RESP_DESC_1_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_2_reg;
               (`RD_RESP_DESC_1_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_3_reg;
               (`RD_RESP_DESC_1_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_4_reg;
               (`RD_RESP_DESC_1_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_5_reg;
               (`RD_RESP_DESC_1_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_6_reg;
               (`RD_RESP_DESC_1_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_7_reg;
               (`RD_RESP_DESC_1_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_8_reg;
               (`RD_RESP_DESC_1_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_9_reg;
               (`RD_RESP_DESC_1_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_10_reg;
               (`RD_RESP_DESC_1_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_11_reg;
               (`RD_RESP_DESC_1_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_12_reg;
               (`RD_RESP_DESC_1_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_13_reg;
               (`RD_RESP_DESC_1_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_14_reg;
               (`RD_RESP_DESC_1_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_1 <= rd_resp_desc_1_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_1 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_2 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_2_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_data_offset_reg;
               (`RD_RESP_DESC_2_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_data_size_reg;
               (`RD_RESP_DESC_2_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_data_host_addr_0_reg;
               (`RD_RESP_DESC_2_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_data_host_addr_1_reg;
               (`RD_RESP_DESC_2_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_data_host_addr_2_reg;
               (`RD_RESP_DESC_2_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_data_host_addr_3_reg;
               (`RD_RESP_DESC_2_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_resp_reg;
               (`RD_RESP_DESC_2_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xid_0_reg;
               (`RD_RESP_DESC_2_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xid_1_reg;
               (`RD_RESP_DESC_2_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xid_2_reg;
               (`RD_RESP_DESC_2_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xid_3_reg;
               (`RD_RESP_DESC_2_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_0_reg;
               (`RD_RESP_DESC_2_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_1_reg;
               (`RD_RESP_DESC_2_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_2_reg;
               (`RD_RESP_DESC_2_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_3_reg;
               (`RD_RESP_DESC_2_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_4_reg;
               (`RD_RESP_DESC_2_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_5_reg;
               (`RD_RESP_DESC_2_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_6_reg;
               (`RD_RESP_DESC_2_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_7_reg;
               (`RD_RESP_DESC_2_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_8_reg;
               (`RD_RESP_DESC_2_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_9_reg;
               (`RD_RESP_DESC_2_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_10_reg;
               (`RD_RESP_DESC_2_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_11_reg;
               (`RD_RESP_DESC_2_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_12_reg;
               (`RD_RESP_DESC_2_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_13_reg;
               (`RD_RESP_DESC_2_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_14_reg;
               (`RD_RESP_DESC_2_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_2 <= rd_resp_desc_2_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_2 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_3 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_3_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_data_offset_reg;
               (`RD_RESP_DESC_3_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_data_size_reg;
               (`RD_RESP_DESC_3_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_data_host_addr_0_reg;
               (`RD_RESP_DESC_3_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_data_host_addr_1_reg;
               (`RD_RESP_DESC_3_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_data_host_addr_2_reg;
               (`RD_RESP_DESC_3_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_data_host_addr_3_reg;
               (`RD_RESP_DESC_3_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_resp_reg;
               (`RD_RESP_DESC_3_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xid_0_reg;
               (`RD_RESP_DESC_3_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xid_1_reg;
               (`RD_RESP_DESC_3_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xid_2_reg;
               (`RD_RESP_DESC_3_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xid_3_reg;
               (`RD_RESP_DESC_3_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_0_reg;
               (`RD_RESP_DESC_3_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_1_reg;
               (`RD_RESP_DESC_3_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_2_reg;
               (`RD_RESP_DESC_3_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_3_reg;
               (`RD_RESP_DESC_3_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_4_reg;
               (`RD_RESP_DESC_3_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_5_reg;
               (`RD_RESP_DESC_3_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_6_reg;
               (`RD_RESP_DESC_3_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_7_reg;
               (`RD_RESP_DESC_3_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_8_reg;
               (`RD_RESP_DESC_3_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_9_reg;
               (`RD_RESP_DESC_3_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_10_reg;
               (`RD_RESP_DESC_3_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_11_reg;
               (`RD_RESP_DESC_3_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_12_reg;
               (`RD_RESP_DESC_3_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_13_reg;
               (`RD_RESP_DESC_3_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_14_reg;
               (`RD_RESP_DESC_3_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_3 <= rd_resp_desc_3_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_3 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_4 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_4_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_data_offset_reg;
               (`RD_RESP_DESC_4_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_data_size_reg;
               (`RD_RESP_DESC_4_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_data_host_addr_0_reg;
               (`RD_RESP_DESC_4_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_data_host_addr_1_reg;
               (`RD_RESP_DESC_4_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_data_host_addr_2_reg;
               (`RD_RESP_DESC_4_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_data_host_addr_3_reg;
               (`RD_RESP_DESC_4_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_resp_reg;
               (`RD_RESP_DESC_4_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xid_0_reg;
               (`RD_RESP_DESC_4_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xid_1_reg;
               (`RD_RESP_DESC_4_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xid_2_reg;
               (`RD_RESP_DESC_4_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xid_3_reg;
               (`RD_RESP_DESC_4_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_0_reg;
               (`RD_RESP_DESC_4_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_1_reg;
               (`RD_RESP_DESC_4_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_2_reg;
               (`RD_RESP_DESC_4_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_3_reg;
               (`RD_RESP_DESC_4_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_4_reg;
               (`RD_RESP_DESC_4_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_5_reg;
               (`RD_RESP_DESC_4_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_6_reg;
               (`RD_RESP_DESC_4_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_7_reg;
               (`RD_RESP_DESC_4_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_8_reg;
               (`RD_RESP_DESC_4_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_9_reg;
               (`RD_RESP_DESC_4_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_10_reg;
               (`RD_RESP_DESC_4_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_11_reg;
               (`RD_RESP_DESC_4_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_12_reg;
               (`RD_RESP_DESC_4_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_13_reg;
               (`RD_RESP_DESC_4_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_14_reg;
               (`RD_RESP_DESC_4_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_4 <= rd_resp_desc_4_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_4 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_5 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_5_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_data_offset_reg;
               (`RD_RESP_DESC_5_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_data_size_reg;
               (`RD_RESP_DESC_5_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_data_host_addr_0_reg;
               (`RD_RESP_DESC_5_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_data_host_addr_1_reg;
               (`RD_RESP_DESC_5_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_data_host_addr_2_reg;
               (`RD_RESP_DESC_5_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_data_host_addr_3_reg;
               (`RD_RESP_DESC_5_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_resp_reg;
               (`RD_RESP_DESC_5_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xid_0_reg;
               (`RD_RESP_DESC_5_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xid_1_reg;
               (`RD_RESP_DESC_5_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xid_2_reg;
               (`RD_RESP_DESC_5_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xid_3_reg;
               (`RD_RESP_DESC_5_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_0_reg;
               (`RD_RESP_DESC_5_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_1_reg;
               (`RD_RESP_DESC_5_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_2_reg;
               (`RD_RESP_DESC_5_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_3_reg;
               (`RD_RESP_DESC_5_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_4_reg;
               (`RD_RESP_DESC_5_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_5_reg;
               (`RD_RESP_DESC_5_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_6_reg;
               (`RD_RESP_DESC_5_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_7_reg;
               (`RD_RESP_DESC_5_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_8_reg;
               (`RD_RESP_DESC_5_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_9_reg;
               (`RD_RESP_DESC_5_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_10_reg;
               (`RD_RESP_DESC_5_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_11_reg;
               (`RD_RESP_DESC_5_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_12_reg;
               (`RD_RESP_DESC_5_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_13_reg;
               (`RD_RESP_DESC_5_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_14_reg;
               (`RD_RESP_DESC_5_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_5 <= rd_resp_desc_5_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_5 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_6 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_6_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_data_offset_reg;
               (`RD_RESP_DESC_6_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_data_size_reg;
               (`RD_RESP_DESC_6_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_data_host_addr_0_reg;
               (`RD_RESP_DESC_6_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_data_host_addr_1_reg;
               (`RD_RESP_DESC_6_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_data_host_addr_2_reg;
               (`RD_RESP_DESC_6_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_data_host_addr_3_reg;
               (`RD_RESP_DESC_6_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_resp_reg;
               (`RD_RESP_DESC_6_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xid_0_reg;
               (`RD_RESP_DESC_6_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xid_1_reg;
               (`RD_RESP_DESC_6_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xid_2_reg;
               (`RD_RESP_DESC_6_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xid_3_reg;
               (`RD_RESP_DESC_6_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_0_reg;
               (`RD_RESP_DESC_6_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_1_reg;
               (`RD_RESP_DESC_6_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_2_reg;
               (`RD_RESP_DESC_6_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_3_reg;
               (`RD_RESP_DESC_6_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_4_reg;
               (`RD_RESP_DESC_6_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_5_reg;
               (`RD_RESP_DESC_6_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_6_reg;
               (`RD_RESP_DESC_6_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_7_reg;
               (`RD_RESP_DESC_6_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_8_reg;
               (`RD_RESP_DESC_6_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_9_reg;
               (`RD_RESP_DESC_6_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_10_reg;
               (`RD_RESP_DESC_6_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_11_reg;
               (`RD_RESP_DESC_6_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_12_reg;
               (`RD_RESP_DESC_6_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_13_reg;
               (`RD_RESP_DESC_6_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_14_reg;
               (`RD_RESP_DESC_6_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_6 <= rd_resp_desc_6_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_6 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_7 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_7_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_data_offset_reg;
               (`RD_RESP_DESC_7_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_data_size_reg;
               (`RD_RESP_DESC_7_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_data_host_addr_0_reg;
               (`RD_RESP_DESC_7_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_data_host_addr_1_reg;
               (`RD_RESP_DESC_7_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_data_host_addr_2_reg;
               (`RD_RESP_DESC_7_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_data_host_addr_3_reg;
               (`RD_RESP_DESC_7_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_resp_reg;
               (`RD_RESP_DESC_7_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xid_0_reg;
               (`RD_RESP_DESC_7_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xid_1_reg;
               (`RD_RESP_DESC_7_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xid_2_reg;
               (`RD_RESP_DESC_7_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xid_3_reg;
               (`RD_RESP_DESC_7_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_0_reg;
               (`RD_RESP_DESC_7_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_1_reg;
               (`RD_RESP_DESC_7_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_2_reg;
               (`RD_RESP_DESC_7_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_3_reg;
               (`RD_RESP_DESC_7_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_4_reg;
               (`RD_RESP_DESC_7_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_5_reg;
               (`RD_RESP_DESC_7_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_6_reg;
               (`RD_RESP_DESC_7_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_7_reg;
               (`RD_RESP_DESC_7_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_8_reg;
               (`RD_RESP_DESC_7_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_9_reg;
               (`RD_RESP_DESC_7_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_10_reg;
               (`RD_RESP_DESC_7_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_11_reg;
               (`RD_RESP_DESC_7_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_12_reg;
               (`RD_RESP_DESC_7_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_13_reg;
               (`RD_RESP_DESC_7_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_14_reg;
               (`RD_RESP_DESC_7_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_7 <= rd_resp_desc_7_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_7 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_8 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_8_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_data_offset_reg;
               (`RD_RESP_DESC_8_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_data_size_reg;
               (`RD_RESP_DESC_8_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_data_host_addr_0_reg;
               (`RD_RESP_DESC_8_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_data_host_addr_1_reg;
               (`RD_RESP_DESC_8_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_data_host_addr_2_reg;
               (`RD_RESP_DESC_8_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_data_host_addr_3_reg;
               (`RD_RESP_DESC_8_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_resp_reg;
               (`RD_RESP_DESC_8_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xid_0_reg;
               (`RD_RESP_DESC_8_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xid_1_reg;
               (`RD_RESP_DESC_8_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xid_2_reg;
               (`RD_RESP_DESC_8_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xid_3_reg;
               (`RD_RESP_DESC_8_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_0_reg;
               (`RD_RESP_DESC_8_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_1_reg;
               (`RD_RESP_DESC_8_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_2_reg;
               (`RD_RESP_DESC_8_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_3_reg;
               (`RD_RESP_DESC_8_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_4_reg;
               (`RD_RESP_DESC_8_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_5_reg;
               (`RD_RESP_DESC_8_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_6_reg;
               (`RD_RESP_DESC_8_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_7_reg;
               (`RD_RESP_DESC_8_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_8_reg;
               (`RD_RESP_DESC_8_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_9_reg;
               (`RD_RESP_DESC_8_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_10_reg;
               (`RD_RESP_DESC_8_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_11_reg;
               (`RD_RESP_DESC_8_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_12_reg;
               (`RD_RESP_DESC_8_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_13_reg;
               (`RD_RESP_DESC_8_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_14_reg;
               (`RD_RESP_DESC_8_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_8 <= rd_resp_desc_8_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_8 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_9 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_9_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_data_offset_reg;
               (`RD_RESP_DESC_9_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_data_size_reg;
               (`RD_RESP_DESC_9_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_data_host_addr_0_reg;
               (`RD_RESP_DESC_9_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_data_host_addr_1_reg;
               (`RD_RESP_DESC_9_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_data_host_addr_2_reg;
               (`RD_RESP_DESC_9_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_data_host_addr_3_reg;
               (`RD_RESP_DESC_9_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_resp_reg;
               (`RD_RESP_DESC_9_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xid_0_reg;
               (`RD_RESP_DESC_9_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xid_1_reg;
               (`RD_RESP_DESC_9_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xid_2_reg;
               (`RD_RESP_DESC_9_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xid_3_reg;
               (`RD_RESP_DESC_9_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_0_reg;
               (`RD_RESP_DESC_9_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_1_reg;
               (`RD_RESP_DESC_9_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_2_reg;
               (`RD_RESP_DESC_9_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_3_reg;
               (`RD_RESP_DESC_9_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_4_reg;
               (`RD_RESP_DESC_9_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_5_reg;
               (`RD_RESP_DESC_9_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_6_reg;
               (`RD_RESP_DESC_9_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_7_reg;
               (`RD_RESP_DESC_9_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_8_reg;
               (`RD_RESP_DESC_9_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_9_reg;
               (`RD_RESP_DESC_9_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_10_reg;
               (`RD_RESP_DESC_9_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_11_reg;
               (`RD_RESP_DESC_9_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_12_reg;
               (`RD_RESP_DESC_9_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_13_reg;
               (`RD_RESP_DESC_9_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_14_reg;
               (`RD_RESP_DESC_9_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_9 <= rd_resp_desc_9_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_9 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_a <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_A_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_data_offset_reg;
               (`RD_RESP_DESC_A_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_data_size_reg;
               (`RD_RESP_DESC_A_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_data_host_addr_0_reg;
               (`RD_RESP_DESC_A_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_data_host_addr_1_reg;
               (`RD_RESP_DESC_A_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_data_host_addr_2_reg;
               (`RD_RESP_DESC_A_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_data_host_addr_3_reg;
               (`RD_RESP_DESC_A_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_resp_reg;
               (`RD_RESP_DESC_A_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xid_0_reg;
               (`RD_RESP_DESC_A_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xid_1_reg;
               (`RD_RESP_DESC_A_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xid_2_reg;
               (`RD_RESP_DESC_A_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xid_3_reg;
               (`RD_RESP_DESC_A_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_0_reg;
               (`RD_RESP_DESC_A_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_1_reg;
               (`RD_RESP_DESC_A_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_2_reg;
               (`RD_RESP_DESC_A_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_3_reg;
               (`RD_RESP_DESC_A_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_4_reg;
               (`RD_RESP_DESC_A_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_5_reg;
               (`RD_RESP_DESC_A_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_6_reg;
               (`RD_RESP_DESC_A_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_7_reg;
               (`RD_RESP_DESC_A_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_8_reg;
               (`RD_RESP_DESC_A_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_9_reg;
               (`RD_RESP_DESC_A_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_10_reg;
               (`RD_RESP_DESC_A_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_11_reg;
               (`RD_RESP_DESC_A_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_12_reg;
               (`RD_RESP_DESC_A_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_13_reg;
               (`RD_RESP_DESC_A_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_14_reg;
               (`RD_RESP_DESC_A_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_a <= rd_resp_desc_a_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_a <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_b <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_B_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_data_offset_reg;
               (`RD_RESP_DESC_B_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_data_size_reg;
               (`RD_RESP_DESC_B_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_data_host_addr_0_reg;
               (`RD_RESP_DESC_B_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_data_host_addr_1_reg;
               (`RD_RESP_DESC_B_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_data_host_addr_2_reg;
               (`RD_RESP_DESC_B_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_data_host_addr_3_reg;
               (`RD_RESP_DESC_B_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_resp_reg;
               (`RD_RESP_DESC_B_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xid_0_reg;
               (`RD_RESP_DESC_B_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xid_1_reg;
               (`RD_RESP_DESC_B_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xid_2_reg;
               (`RD_RESP_DESC_B_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xid_3_reg;
               (`RD_RESP_DESC_B_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_0_reg;
               (`RD_RESP_DESC_B_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_1_reg;
               (`RD_RESP_DESC_B_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_2_reg;
               (`RD_RESP_DESC_B_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_3_reg;
               (`RD_RESP_DESC_B_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_4_reg;
               (`RD_RESP_DESC_B_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_5_reg;
               (`RD_RESP_DESC_B_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_6_reg;
               (`RD_RESP_DESC_B_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_7_reg;
               (`RD_RESP_DESC_B_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_8_reg;
               (`RD_RESP_DESC_B_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_9_reg;
               (`RD_RESP_DESC_B_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_10_reg;
               (`RD_RESP_DESC_B_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_11_reg;
               (`RD_RESP_DESC_B_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_12_reg;
               (`RD_RESP_DESC_B_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_13_reg;
               (`RD_RESP_DESC_B_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_14_reg;
               (`RD_RESP_DESC_B_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_b <= rd_resp_desc_b_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_b <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_c <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_C_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_data_offset_reg;
               (`RD_RESP_DESC_C_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_data_size_reg;
               (`RD_RESP_DESC_C_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_data_host_addr_0_reg;
               (`RD_RESP_DESC_C_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_data_host_addr_1_reg;
               (`RD_RESP_DESC_C_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_data_host_addr_2_reg;
               (`RD_RESP_DESC_C_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_data_host_addr_3_reg;
               (`RD_RESP_DESC_C_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_resp_reg;
               (`RD_RESP_DESC_C_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xid_0_reg;
               (`RD_RESP_DESC_C_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xid_1_reg;
               (`RD_RESP_DESC_C_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xid_2_reg;
               (`RD_RESP_DESC_C_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xid_3_reg;
               (`RD_RESP_DESC_C_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_0_reg;
               (`RD_RESP_DESC_C_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_1_reg;
               (`RD_RESP_DESC_C_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_2_reg;
               (`RD_RESP_DESC_C_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_3_reg;
               (`RD_RESP_DESC_C_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_4_reg;
               (`RD_RESP_DESC_C_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_5_reg;
               (`RD_RESP_DESC_C_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_6_reg;
               (`RD_RESP_DESC_C_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_7_reg;
               (`RD_RESP_DESC_C_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_8_reg;
               (`RD_RESP_DESC_C_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_9_reg;
               (`RD_RESP_DESC_C_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_10_reg;
               (`RD_RESP_DESC_C_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_11_reg;
               (`RD_RESP_DESC_C_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_12_reg;
               (`RD_RESP_DESC_C_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_13_reg;
               (`RD_RESP_DESC_C_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_14_reg;
               (`RD_RESP_DESC_C_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_c <= rd_resp_desc_c_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_c <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_d <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_D_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_data_offset_reg;
               (`RD_RESP_DESC_D_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_data_size_reg;
               (`RD_RESP_DESC_D_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_data_host_addr_0_reg;
               (`RD_RESP_DESC_D_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_data_host_addr_1_reg;
               (`RD_RESP_DESC_D_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_data_host_addr_2_reg;
               (`RD_RESP_DESC_D_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_data_host_addr_3_reg;
               (`RD_RESP_DESC_D_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_resp_reg;
               (`RD_RESP_DESC_D_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xid_0_reg;
               (`RD_RESP_DESC_D_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xid_1_reg;
               (`RD_RESP_DESC_D_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xid_2_reg;
               (`RD_RESP_DESC_D_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xid_3_reg;
               (`RD_RESP_DESC_D_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_0_reg;
               (`RD_RESP_DESC_D_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_1_reg;
               (`RD_RESP_DESC_D_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_2_reg;
               (`RD_RESP_DESC_D_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_3_reg;
               (`RD_RESP_DESC_D_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_4_reg;
               (`RD_RESP_DESC_D_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_5_reg;
               (`RD_RESP_DESC_D_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_6_reg;
               (`RD_RESP_DESC_D_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_7_reg;
               (`RD_RESP_DESC_D_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_8_reg;
               (`RD_RESP_DESC_D_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_9_reg;
               (`RD_RESP_DESC_D_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_10_reg;
               (`RD_RESP_DESC_D_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_11_reg;
               (`RD_RESP_DESC_D_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_12_reg;
               (`RD_RESP_DESC_D_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_13_reg;
               (`RD_RESP_DESC_D_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_14_reg;
               (`RD_RESP_DESC_D_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_d <= rd_resp_desc_d_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_d <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_e <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_E_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_data_offset_reg;
               (`RD_RESP_DESC_E_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_data_size_reg;
               (`RD_RESP_DESC_E_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_data_host_addr_0_reg;
               (`RD_RESP_DESC_E_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_data_host_addr_1_reg;
               (`RD_RESP_DESC_E_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_data_host_addr_2_reg;
               (`RD_RESP_DESC_E_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_data_host_addr_3_reg;
               (`RD_RESP_DESC_E_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_resp_reg;
               (`RD_RESP_DESC_E_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xid_0_reg;
               (`RD_RESP_DESC_E_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xid_1_reg;
               (`RD_RESP_DESC_E_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xid_2_reg;
               (`RD_RESP_DESC_E_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xid_3_reg;
               (`RD_RESP_DESC_E_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_0_reg;
               (`RD_RESP_DESC_E_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_1_reg;
               (`RD_RESP_DESC_E_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_2_reg;
               (`RD_RESP_DESC_E_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_3_reg;
               (`RD_RESP_DESC_E_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_4_reg;
               (`RD_RESP_DESC_E_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_5_reg;
               (`RD_RESP_DESC_E_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_6_reg;
               (`RD_RESP_DESC_E_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_7_reg;
               (`RD_RESP_DESC_E_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_8_reg;
               (`RD_RESP_DESC_E_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_9_reg;
               (`RD_RESP_DESC_E_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_10_reg;
               (`RD_RESP_DESC_E_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_11_reg;
               (`RD_RESP_DESC_E_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_12_reg;
               (`RD_RESP_DESC_E_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_13_reg;
               (`RD_RESP_DESC_E_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_14_reg;
               (`RD_RESP_DESC_E_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_e <= rd_resp_desc_e_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_e <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_rd_resp_desc_f <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`RD_RESP_DESC_F_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_data_offset_reg;
               (`RD_RESP_DESC_F_DATA_SIZE_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_data_size_reg;
               (`RD_RESP_DESC_F_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_data_host_addr_0_reg;
               (`RD_RESP_DESC_F_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_data_host_addr_1_reg;
               (`RD_RESP_DESC_F_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_data_host_addr_2_reg;
               (`RD_RESP_DESC_F_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_data_host_addr_3_reg;
               (`RD_RESP_DESC_F_RESP_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_resp_reg;
               (`RD_RESP_DESC_F_XID_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xid_0_reg;
               (`RD_RESP_DESC_F_XID_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xid_1_reg;
               (`RD_RESP_DESC_F_XID_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xid_2_reg;
               (`RD_RESP_DESC_F_XID_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xid_3_reg;
               (`RD_RESP_DESC_F_XUSER_0_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_0_reg;
               (`RD_RESP_DESC_F_XUSER_1_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_1_reg;
               (`RD_RESP_DESC_F_XUSER_2_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_2_reg;
               (`RD_RESP_DESC_F_XUSER_3_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_3_reg;
               (`RD_RESP_DESC_F_XUSER_4_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_4_reg;
               (`RD_RESP_DESC_F_XUSER_5_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_5_reg;
               (`RD_RESP_DESC_F_XUSER_6_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_6_reg;
               (`RD_RESP_DESC_F_XUSER_7_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_7_reg;
               (`RD_RESP_DESC_F_XUSER_8_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_8_reg;
               (`RD_RESP_DESC_F_XUSER_9_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_9_reg;
               (`RD_RESP_DESC_F_XUSER_10_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_10_reg;
               (`RD_RESP_DESC_F_XUSER_11_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_11_reg;
               (`RD_RESP_DESC_F_XUSER_12_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_12_reg;
               (`RD_RESP_DESC_F_XUSER_13_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_13_reg;
               (`RD_RESP_DESC_F_XUSER_14_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_14_reg;
               (`RD_RESP_DESC_F_XUSER_15_REG_ADDR&'hFF) :reg_data_out_rd_resp_desc_f <= rd_resp_desc_f_xuser_15_reg;
               default                                  :reg_data_out_rd_resp_desc_f <= 32'b0      ;        
             endcase
	  end
     end




   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_0 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_0_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_txn_type_reg;
               (`WR_REQ_DESC_0_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_size_reg;
               (`WR_REQ_DESC_0_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_data_offset_reg;
               (`WR_REQ_DESC_0_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_data_host_addr_0_reg;
               (`WR_REQ_DESC_0_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_data_host_addr_1_reg;
               (`WR_REQ_DESC_0_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_data_host_addr_2_reg;
               (`WR_REQ_DESC_0_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_data_host_addr_3_reg;
               (`WR_REQ_DESC_0_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_0_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_0_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_0_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_0_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axsize_reg;
               (`WR_REQ_DESC_0_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_attr_reg;
               (`WR_REQ_DESC_0_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axaddr_0_reg;
               (`WR_REQ_DESC_0_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axaddr_1_reg;
               (`WR_REQ_DESC_0_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axaddr_2_reg;
               (`WR_REQ_DESC_0_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axaddr_3_reg;
               (`WR_REQ_DESC_0_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axid_0_reg;
               (`WR_REQ_DESC_0_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axid_1_reg;
               (`WR_REQ_DESC_0_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axid_2_reg;
               (`WR_REQ_DESC_0_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axid_3_reg;
               (`WR_REQ_DESC_0_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_0_reg;
               (`WR_REQ_DESC_0_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_1_reg;
               (`WR_REQ_DESC_0_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_2_reg;
               (`WR_REQ_DESC_0_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_3_reg;
               (`WR_REQ_DESC_0_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_4_reg;
               (`WR_REQ_DESC_0_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_5_reg;
               (`WR_REQ_DESC_0_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_6_reg;
               (`WR_REQ_DESC_0_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_7_reg;
               (`WR_REQ_DESC_0_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_8_reg;
               (`WR_REQ_DESC_0_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_9_reg;
               (`WR_REQ_DESC_0_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_10_reg;
               (`WR_REQ_DESC_0_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_11_reg;
               (`WR_REQ_DESC_0_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_12_reg;
               (`WR_REQ_DESC_0_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_13_reg;
               (`WR_REQ_DESC_0_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_14_reg;
               (`WR_REQ_DESC_0_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_axuser_15_reg;
               (`WR_REQ_DESC_0_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_0_reg;
               (`WR_REQ_DESC_0_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_1_reg;
               (`WR_REQ_DESC_0_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_2_reg;
               (`WR_REQ_DESC_0_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_3_reg;
               (`WR_REQ_DESC_0_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_4_reg;
               (`WR_REQ_DESC_0_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_5_reg;
               (`WR_REQ_DESC_0_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_6_reg;
               (`WR_REQ_DESC_0_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_7_reg;
               (`WR_REQ_DESC_0_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_8_reg;
               (`WR_REQ_DESC_0_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_9_reg;
               (`WR_REQ_DESC_0_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_10_reg;
               (`WR_REQ_DESC_0_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_11_reg;
               (`WR_REQ_DESC_0_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_12_reg;
               (`WR_REQ_DESC_0_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_13_reg;
               (`WR_REQ_DESC_0_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_14_reg;
               (`WR_REQ_DESC_0_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_0 <= wr_req_desc_0_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_0 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_1 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_1_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_txn_type_reg;
               (`WR_REQ_DESC_1_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_size_reg;
               (`WR_REQ_DESC_1_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_data_offset_reg;
               (`WR_REQ_DESC_1_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_data_host_addr_0_reg;
               (`WR_REQ_DESC_1_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_data_host_addr_1_reg;
               (`WR_REQ_DESC_1_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_data_host_addr_2_reg;
               (`WR_REQ_DESC_1_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_data_host_addr_3_reg;
               (`WR_REQ_DESC_1_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_1_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_1_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_1_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_1_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axsize_reg;
               (`WR_REQ_DESC_1_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_attr_reg;
               (`WR_REQ_DESC_1_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axaddr_0_reg;
               (`WR_REQ_DESC_1_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axaddr_1_reg;
               (`WR_REQ_DESC_1_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axaddr_2_reg;
               (`WR_REQ_DESC_1_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axaddr_3_reg;
               (`WR_REQ_DESC_1_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axid_0_reg;
               (`WR_REQ_DESC_1_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axid_1_reg;
               (`WR_REQ_DESC_1_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axid_2_reg;
               (`WR_REQ_DESC_1_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axid_3_reg;
               (`WR_REQ_DESC_1_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_0_reg;
               (`WR_REQ_DESC_1_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_1_reg;
               (`WR_REQ_DESC_1_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_2_reg;
               (`WR_REQ_DESC_1_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_3_reg;
               (`WR_REQ_DESC_1_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_4_reg;
               (`WR_REQ_DESC_1_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_5_reg;
               (`WR_REQ_DESC_1_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_6_reg;
               (`WR_REQ_DESC_1_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_7_reg;
               (`WR_REQ_DESC_1_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_8_reg;
               (`WR_REQ_DESC_1_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_9_reg;
               (`WR_REQ_DESC_1_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_10_reg;
               (`WR_REQ_DESC_1_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_11_reg;
               (`WR_REQ_DESC_1_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_12_reg;
               (`WR_REQ_DESC_1_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_13_reg;
               (`WR_REQ_DESC_1_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_14_reg;
               (`WR_REQ_DESC_1_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_axuser_15_reg;
               (`WR_REQ_DESC_1_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_0_reg;
               (`WR_REQ_DESC_1_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_1_reg;
               (`WR_REQ_DESC_1_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_2_reg;
               (`WR_REQ_DESC_1_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_3_reg;
               (`WR_REQ_DESC_1_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_4_reg;
               (`WR_REQ_DESC_1_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_5_reg;
               (`WR_REQ_DESC_1_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_6_reg;
               (`WR_REQ_DESC_1_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_7_reg;
               (`WR_REQ_DESC_1_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_8_reg;
               (`WR_REQ_DESC_1_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_9_reg;
               (`WR_REQ_DESC_1_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_10_reg;
               (`WR_REQ_DESC_1_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_11_reg;
               (`WR_REQ_DESC_1_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_12_reg;
               (`WR_REQ_DESC_1_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_13_reg;
               (`WR_REQ_DESC_1_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_14_reg;
               (`WR_REQ_DESC_1_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_1 <= wr_req_desc_1_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_1 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_2 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_2_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_txn_type_reg;
               (`WR_REQ_DESC_2_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_size_reg;
               (`WR_REQ_DESC_2_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_data_offset_reg;
               (`WR_REQ_DESC_2_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_data_host_addr_0_reg;
               (`WR_REQ_DESC_2_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_data_host_addr_1_reg;
               (`WR_REQ_DESC_2_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_data_host_addr_2_reg;
               (`WR_REQ_DESC_2_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_data_host_addr_3_reg;
               (`WR_REQ_DESC_2_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_2_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_2_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_2_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_2_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axsize_reg;
               (`WR_REQ_DESC_2_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_attr_reg;
               (`WR_REQ_DESC_2_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axaddr_0_reg;
               (`WR_REQ_DESC_2_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axaddr_1_reg;
               (`WR_REQ_DESC_2_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axaddr_2_reg;
               (`WR_REQ_DESC_2_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axaddr_3_reg;
               (`WR_REQ_DESC_2_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axid_0_reg;
               (`WR_REQ_DESC_2_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axid_1_reg;
               (`WR_REQ_DESC_2_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axid_2_reg;
               (`WR_REQ_DESC_2_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axid_3_reg;
               (`WR_REQ_DESC_2_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_0_reg;
               (`WR_REQ_DESC_2_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_1_reg;
               (`WR_REQ_DESC_2_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_2_reg;
               (`WR_REQ_DESC_2_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_3_reg;
               (`WR_REQ_DESC_2_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_4_reg;
               (`WR_REQ_DESC_2_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_5_reg;
               (`WR_REQ_DESC_2_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_6_reg;
               (`WR_REQ_DESC_2_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_7_reg;
               (`WR_REQ_DESC_2_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_8_reg;
               (`WR_REQ_DESC_2_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_9_reg;
               (`WR_REQ_DESC_2_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_10_reg;
               (`WR_REQ_DESC_2_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_11_reg;
               (`WR_REQ_DESC_2_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_12_reg;
               (`WR_REQ_DESC_2_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_13_reg;
               (`WR_REQ_DESC_2_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_14_reg;
               (`WR_REQ_DESC_2_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_axuser_15_reg;
               (`WR_REQ_DESC_2_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_0_reg;
               (`WR_REQ_DESC_2_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_1_reg;
               (`WR_REQ_DESC_2_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_2_reg;
               (`WR_REQ_DESC_2_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_3_reg;
               (`WR_REQ_DESC_2_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_4_reg;
               (`WR_REQ_DESC_2_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_5_reg;
               (`WR_REQ_DESC_2_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_6_reg;
               (`WR_REQ_DESC_2_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_7_reg;
               (`WR_REQ_DESC_2_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_8_reg;
               (`WR_REQ_DESC_2_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_9_reg;
               (`WR_REQ_DESC_2_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_10_reg;
               (`WR_REQ_DESC_2_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_11_reg;
               (`WR_REQ_DESC_2_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_12_reg;
               (`WR_REQ_DESC_2_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_13_reg;
               (`WR_REQ_DESC_2_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_14_reg;
               (`WR_REQ_DESC_2_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_2 <= wr_req_desc_2_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_2 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_3 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_3_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_txn_type_reg;
               (`WR_REQ_DESC_3_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_size_reg;
               (`WR_REQ_DESC_3_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_data_offset_reg;
               (`WR_REQ_DESC_3_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_data_host_addr_0_reg;
               (`WR_REQ_DESC_3_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_data_host_addr_1_reg;
               (`WR_REQ_DESC_3_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_data_host_addr_2_reg;
               (`WR_REQ_DESC_3_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_data_host_addr_3_reg;
               (`WR_REQ_DESC_3_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_3_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_3_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_3_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_3_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axsize_reg;
               (`WR_REQ_DESC_3_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_attr_reg;
               (`WR_REQ_DESC_3_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axaddr_0_reg;
               (`WR_REQ_DESC_3_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axaddr_1_reg;
               (`WR_REQ_DESC_3_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axaddr_2_reg;
               (`WR_REQ_DESC_3_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axaddr_3_reg;
               (`WR_REQ_DESC_3_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axid_0_reg;
               (`WR_REQ_DESC_3_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axid_1_reg;
               (`WR_REQ_DESC_3_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axid_2_reg;
               (`WR_REQ_DESC_3_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axid_3_reg;
               (`WR_REQ_DESC_3_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_0_reg;
               (`WR_REQ_DESC_3_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_1_reg;
               (`WR_REQ_DESC_3_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_2_reg;
               (`WR_REQ_DESC_3_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_3_reg;
               (`WR_REQ_DESC_3_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_4_reg;
               (`WR_REQ_DESC_3_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_5_reg;
               (`WR_REQ_DESC_3_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_6_reg;
               (`WR_REQ_DESC_3_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_7_reg;
               (`WR_REQ_DESC_3_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_8_reg;
               (`WR_REQ_DESC_3_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_9_reg;
               (`WR_REQ_DESC_3_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_10_reg;
               (`WR_REQ_DESC_3_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_11_reg;
               (`WR_REQ_DESC_3_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_12_reg;
               (`WR_REQ_DESC_3_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_13_reg;
               (`WR_REQ_DESC_3_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_14_reg;
               (`WR_REQ_DESC_3_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_axuser_15_reg;
               (`WR_REQ_DESC_3_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_0_reg;
               (`WR_REQ_DESC_3_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_1_reg;
               (`WR_REQ_DESC_3_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_2_reg;
               (`WR_REQ_DESC_3_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_3_reg;
               (`WR_REQ_DESC_3_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_4_reg;
               (`WR_REQ_DESC_3_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_5_reg;
               (`WR_REQ_DESC_3_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_6_reg;
               (`WR_REQ_DESC_3_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_7_reg;
               (`WR_REQ_DESC_3_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_8_reg;
               (`WR_REQ_DESC_3_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_9_reg;
               (`WR_REQ_DESC_3_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_10_reg;
               (`WR_REQ_DESC_3_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_11_reg;
               (`WR_REQ_DESC_3_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_12_reg;
               (`WR_REQ_DESC_3_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_13_reg;
               (`WR_REQ_DESC_3_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_14_reg;
               (`WR_REQ_DESC_3_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_3 <= wr_req_desc_3_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_3 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_4 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_4_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_txn_type_reg;
               (`WR_REQ_DESC_4_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_size_reg;
               (`WR_REQ_DESC_4_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_data_offset_reg;
               (`WR_REQ_DESC_4_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_data_host_addr_0_reg;
               (`WR_REQ_DESC_4_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_data_host_addr_1_reg;
               (`WR_REQ_DESC_4_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_data_host_addr_2_reg;
               (`WR_REQ_DESC_4_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_data_host_addr_3_reg;
               (`WR_REQ_DESC_4_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_4_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_4_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_4_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_4_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axsize_reg;
               (`WR_REQ_DESC_4_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_attr_reg;
               (`WR_REQ_DESC_4_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axaddr_0_reg;
               (`WR_REQ_DESC_4_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axaddr_1_reg;
               (`WR_REQ_DESC_4_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axaddr_2_reg;
               (`WR_REQ_DESC_4_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axaddr_3_reg;
               (`WR_REQ_DESC_4_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axid_0_reg;
               (`WR_REQ_DESC_4_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axid_1_reg;
               (`WR_REQ_DESC_4_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axid_2_reg;
               (`WR_REQ_DESC_4_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axid_3_reg;
               (`WR_REQ_DESC_4_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_0_reg;
               (`WR_REQ_DESC_4_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_1_reg;
               (`WR_REQ_DESC_4_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_2_reg;
               (`WR_REQ_DESC_4_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_3_reg;
               (`WR_REQ_DESC_4_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_4_reg;
               (`WR_REQ_DESC_4_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_5_reg;
               (`WR_REQ_DESC_4_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_6_reg;
               (`WR_REQ_DESC_4_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_7_reg;
               (`WR_REQ_DESC_4_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_8_reg;
               (`WR_REQ_DESC_4_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_9_reg;
               (`WR_REQ_DESC_4_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_10_reg;
               (`WR_REQ_DESC_4_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_11_reg;
               (`WR_REQ_DESC_4_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_12_reg;
               (`WR_REQ_DESC_4_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_13_reg;
               (`WR_REQ_DESC_4_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_14_reg;
               (`WR_REQ_DESC_4_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_axuser_15_reg;
               (`WR_REQ_DESC_4_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_0_reg;
               (`WR_REQ_DESC_4_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_1_reg;
               (`WR_REQ_DESC_4_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_2_reg;
               (`WR_REQ_DESC_4_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_3_reg;
               (`WR_REQ_DESC_4_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_4_reg;
               (`WR_REQ_DESC_4_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_5_reg;
               (`WR_REQ_DESC_4_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_6_reg;
               (`WR_REQ_DESC_4_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_7_reg;
               (`WR_REQ_DESC_4_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_8_reg;
               (`WR_REQ_DESC_4_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_9_reg;
               (`WR_REQ_DESC_4_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_10_reg;
               (`WR_REQ_DESC_4_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_11_reg;
               (`WR_REQ_DESC_4_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_12_reg;
               (`WR_REQ_DESC_4_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_13_reg;
               (`WR_REQ_DESC_4_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_14_reg;
               (`WR_REQ_DESC_4_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_4 <= wr_req_desc_4_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_4 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_5 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_5_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_txn_type_reg;
               (`WR_REQ_DESC_5_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_size_reg;
               (`WR_REQ_DESC_5_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_data_offset_reg;
               (`WR_REQ_DESC_5_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_data_host_addr_0_reg;
               (`WR_REQ_DESC_5_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_data_host_addr_1_reg;
               (`WR_REQ_DESC_5_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_data_host_addr_2_reg;
               (`WR_REQ_DESC_5_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_data_host_addr_3_reg;
               (`WR_REQ_DESC_5_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_5_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_5_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_5_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_5_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axsize_reg;
               (`WR_REQ_DESC_5_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_attr_reg;
               (`WR_REQ_DESC_5_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axaddr_0_reg;
               (`WR_REQ_DESC_5_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axaddr_1_reg;
               (`WR_REQ_DESC_5_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axaddr_2_reg;
               (`WR_REQ_DESC_5_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axaddr_3_reg;
               (`WR_REQ_DESC_5_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axid_0_reg;
               (`WR_REQ_DESC_5_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axid_1_reg;
               (`WR_REQ_DESC_5_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axid_2_reg;
               (`WR_REQ_DESC_5_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axid_3_reg;
               (`WR_REQ_DESC_5_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_0_reg;
               (`WR_REQ_DESC_5_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_1_reg;
               (`WR_REQ_DESC_5_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_2_reg;
               (`WR_REQ_DESC_5_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_3_reg;
               (`WR_REQ_DESC_5_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_4_reg;
               (`WR_REQ_DESC_5_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_5_reg;
               (`WR_REQ_DESC_5_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_6_reg;
               (`WR_REQ_DESC_5_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_7_reg;
               (`WR_REQ_DESC_5_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_8_reg;
               (`WR_REQ_DESC_5_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_9_reg;
               (`WR_REQ_DESC_5_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_10_reg;
               (`WR_REQ_DESC_5_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_11_reg;
               (`WR_REQ_DESC_5_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_12_reg;
               (`WR_REQ_DESC_5_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_13_reg;
               (`WR_REQ_DESC_5_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_14_reg;
               (`WR_REQ_DESC_5_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_axuser_15_reg;
               (`WR_REQ_DESC_5_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_0_reg;
               (`WR_REQ_DESC_5_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_1_reg;
               (`WR_REQ_DESC_5_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_2_reg;
               (`WR_REQ_DESC_5_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_3_reg;
               (`WR_REQ_DESC_5_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_4_reg;
               (`WR_REQ_DESC_5_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_5_reg;
               (`WR_REQ_DESC_5_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_6_reg;
               (`WR_REQ_DESC_5_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_7_reg;
               (`WR_REQ_DESC_5_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_8_reg;
               (`WR_REQ_DESC_5_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_9_reg;
               (`WR_REQ_DESC_5_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_10_reg;
               (`WR_REQ_DESC_5_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_11_reg;
               (`WR_REQ_DESC_5_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_12_reg;
               (`WR_REQ_DESC_5_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_13_reg;
               (`WR_REQ_DESC_5_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_14_reg;
               (`WR_REQ_DESC_5_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_5 <= wr_req_desc_5_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_5 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_6 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_6_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_txn_type_reg;
               (`WR_REQ_DESC_6_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_size_reg;
               (`WR_REQ_DESC_6_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_data_offset_reg;
               (`WR_REQ_DESC_6_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_data_host_addr_0_reg;
               (`WR_REQ_DESC_6_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_data_host_addr_1_reg;
               (`WR_REQ_DESC_6_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_data_host_addr_2_reg;
               (`WR_REQ_DESC_6_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_data_host_addr_3_reg;
               (`WR_REQ_DESC_6_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_6_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_6_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_6_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_6_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axsize_reg;
               (`WR_REQ_DESC_6_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_attr_reg;
               (`WR_REQ_DESC_6_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axaddr_0_reg;
               (`WR_REQ_DESC_6_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axaddr_1_reg;
               (`WR_REQ_DESC_6_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axaddr_2_reg;
               (`WR_REQ_DESC_6_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axaddr_3_reg;
               (`WR_REQ_DESC_6_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axid_0_reg;
               (`WR_REQ_DESC_6_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axid_1_reg;
               (`WR_REQ_DESC_6_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axid_2_reg;
               (`WR_REQ_DESC_6_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axid_3_reg;
               (`WR_REQ_DESC_6_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_0_reg;
               (`WR_REQ_DESC_6_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_1_reg;
               (`WR_REQ_DESC_6_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_2_reg;
               (`WR_REQ_DESC_6_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_3_reg;
               (`WR_REQ_DESC_6_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_4_reg;
               (`WR_REQ_DESC_6_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_5_reg;
               (`WR_REQ_DESC_6_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_6_reg;
               (`WR_REQ_DESC_6_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_7_reg;
               (`WR_REQ_DESC_6_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_8_reg;
               (`WR_REQ_DESC_6_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_9_reg;
               (`WR_REQ_DESC_6_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_10_reg;
               (`WR_REQ_DESC_6_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_11_reg;
               (`WR_REQ_DESC_6_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_12_reg;
               (`WR_REQ_DESC_6_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_13_reg;
               (`WR_REQ_DESC_6_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_14_reg;
               (`WR_REQ_DESC_6_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_axuser_15_reg;
               (`WR_REQ_DESC_6_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_0_reg;
               (`WR_REQ_DESC_6_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_1_reg;
               (`WR_REQ_DESC_6_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_2_reg;
               (`WR_REQ_DESC_6_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_3_reg;
               (`WR_REQ_DESC_6_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_4_reg;
               (`WR_REQ_DESC_6_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_5_reg;
               (`WR_REQ_DESC_6_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_6_reg;
               (`WR_REQ_DESC_6_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_7_reg;
               (`WR_REQ_DESC_6_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_8_reg;
               (`WR_REQ_DESC_6_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_9_reg;
               (`WR_REQ_DESC_6_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_10_reg;
               (`WR_REQ_DESC_6_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_11_reg;
               (`WR_REQ_DESC_6_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_12_reg;
               (`WR_REQ_DESC_6_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_13_reg;
               (`WR_REQ_DESC_6_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_14_reg;
               (`WR_REQ_DESC_6_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_6 <= wr_req_desc_6_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_6 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_7 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_7_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_txn_type_reg;
               (`WR_REQ_DESC_7_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_size_reg;
               (`WR_REQ_DESC_7_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_data_offset_reg;
               (`WR_REQ_DESC_7_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_data_host_addr_0_reg;
               (`WR_REQ_DESC_7_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_data_host_addr_1_reg;
               (`WR_REQ_DESC_7_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_data_host_addr_2_reg;
               (`WR_REQ_DESC_7_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_data_host_addr_3_reg;
               (`WR_REQ_DESC_7_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_7_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_7_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_7_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_7_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axsize_reg;
               (`WR_REQ_DESC_7_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_attr_reg;
               (`WR_REQ_DESC_7_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axaddr_0_reg;
               (`WR_REQ_DESC_7_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axaddr_1_reg;
               (`WR_REQ_DESC_7_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axaddr_2_reg;
               (`WR_REQ_DESC_7_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axaddr_3_reg;
               (`WR_REQ_DESC_7_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axid_0_reg;
               (`WR_REQ_DESC_7_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axid_1_reg;
               (`WR_REQ_DESC_7_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axid_2_reg;
               (`WR_REQ_DESC_7_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axid_3_reg;
               (`WR_REQ_DESC_7_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_0_reg;
               (`WR_REQ_DESC_7_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_1_reg;
               (`WR_REQ_DESC_7_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_2_reg;
               (`WR_REQ_DESC_7_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_3_reg;
               (`WR_REQ_DESC_7_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_4_reg;
               (`WR_REQ_DESC_7_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_5_reg;
               (`WR_REQ_DESC_7_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_6_reg;
               (`WR_REQ_DESC_7_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_7_reg;
               (`WR_REQ_DESC_7_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_8_reg;
               (`WR_REQ_DESC_7_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_9_reg;
               (`WR_REQ_DESC_7_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_10_reg;
               (`WR_REQ_DESC_7_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_11_reg;
               (`WR_REQ_DESC_7_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_12_reg;
               (`WR_REQ_DESC_7_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_13_reg;
               (`WR_REQ_DESC_7_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_14_reg;
               (`WR_REQ_DESC_7_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_axuser_15_reg;
               (`WR_REQ_DESC_7_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_0_reg;
               (`WR_REQ_DESC_7_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_1_reg;
               (`WR_REQ_DESC_7_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_2_reg;
               (`WR_REQ_DESC_7_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_3_reg;
               (`WR_REQ_DESC_7_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_4_reg;
               (`WR_REQ_DESC_7_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_5_reg;
               (`WR_REQ_DESC_7_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_6_reg;
               (`WR_REQ_DESC_7_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_7_reg;
               (`WR_REQ_DESC_7_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_8_reg;
               (`WR_REQ_DESC_7_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_9_reg;
               (`WR_REQ_DESC_7_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_10_reg;
               (`WR_REQ_DESC_7_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_11_reg;
               (`WR_REQ_DESC_7_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_12_reg;
               (`WR_REQ_DESC_7_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_13_reg;
               (`WR_REQ_DESC_7_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_14_reg;
               (`WR_REQ_DESC_7_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_7 <= wr_req_desc_7_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_7 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_8 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_8_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_txn_type_reg;
               (`WR_REQ_DESC_8_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_size_reg;
               (`WR_REQ_DESC_8_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_data_offset_reg;
               (`WR_REQ_DESC_8_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_data_host_addr_0_reg;
               (`WR_REQ_DESC_8_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_data_host_addr_1_reg;
               (`WR_REQ_DESC_8_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_data_host_addr_2_reg;
               (`WR_REQ_DESC_8_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_data_host_addr_3_reg;
               (`WR_REQ_DESC_8_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_8_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_8_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_8_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_8_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axsize_reg;
               (`WR_REQ_DESC_8_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_attr_reg;
               (`WR_REQ_DESC_8_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axaddr_0_reg;
               (`WR_REQ_DESC_8_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axaddr_1_reg;
               (`WR_REQ_DESC_8_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axaddr_2_reg;
               (`WR_REQ_DESC_8_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axaddr_3_reg;
               (`WR_REQ_DESC_8_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axid_0_reg;
               (`WR_REQ_DESC_8_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axid_1_reg;
               (`WR_REQ_DESC_8_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axid_2_reg;
               (`WR_REQ_DESC_8_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axid_3_reg;
               (`WR_REQ_DESC_8_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_0_reg;
               (`WR_REQ_DESC_8_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_1_reg;
               (`WR_REQ_DESC_8_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_2_reg;
               (`WR_REQ_DESC_8_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_3_reg;
               (`WR_REQ_DESC_8_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_4_reg;
               (`WR_REQ_DESC_8_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_5_reg;
               (`WR_REQ_DESC_8_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_6_reg;
               (`WR_REQ_DESC_8_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_7_reg;
               (`WR_REQ_DESC_8_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_8_reg;
               (`WR_REQ_DESC_8_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_9_reg;
               (`WR_REQ_DESC_8_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_10_reg;
               (`WR_REQ_DESC_8_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_11_reg;
               (`WR_REQ_DESC_8_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_12_reg;
               (`WR_REQ_DESC_8_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_13_reg;
               (`WR_REQ_DESC_8_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_14_reg;
               (`WR_REQ_DESC_8_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_axuser_15_reg;
               (`WR_REQ_DESC_8_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_0_reg;
               (`WR_REQ_DESC_8_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_1_reg;
               (`WR_REQ_DESC_8_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_2_reg;
               (`WR_REQ_DESC_8_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_3_reg;
               (`WR_REQ_DESC_8_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_4_reg;
               (`WR_REQ_DESC_8_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_5_reg;
               (`WR_REQ_DESC_8_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_6_reg;
               (`WR_REQ_DESC_8_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_7_reg;
               (`WR_REQ_DESC_8_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_8_reg;
               (`WR_REQ_DESC_8_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_9_reg;
               (`WR_REQ_DESC_8_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_10_reg;
               (`WR_REQ_DESC_8_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_11_reg;
               (`WR_REQ_DESC_8_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_12_reg;
               (`WR_REQ_DESC_8_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_13_reg;
               (`WR_REQ_DESC_8_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_14_reg;
               (`WR_REQ_DESC_8_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_8 <= wr_req_desc_8_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_8 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_9 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_9_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_txn_type_reg;
               (`WR_REQ_DESC_9_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_size_reg;
               (`WR_REQ_DESC_9_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_data_offset_reg;
               (`WR_REQ_DESC_9_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_data_host_addr_0_reg;
               (`WR_REQ_DESC_9_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_data_host_addr_1_reg;
               (`WR_REQ_DESC_9_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_data_host_addr_2_reg;
               (`WR_REQ_DESC_9_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_data_host_addr_3_reg;
               (`WR_REQ_DESC_9_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_9_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_9_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_9_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_9_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axsize_reg;
               (`WR_REQ_DESC_9_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_attr_reg;
               (`WR_REQ_DESC_9_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axaddr_0_reg;
               (`WR_REQ_DESC_9_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axaddr_1_reg;
               (`WR_REQ_DESC_9_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axaddr_2_reg;
               (`WR_REQ_DESC_9_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axaddr_3_reg;
               (`WR_REQ_DESC_9_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axid_0_reg;
               (`WR_REQ_DESC_9_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axid_1_reg;
               (`WR_REQ_DESC_9_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axid_2_reg;
               (`WR_REQ_DESC_9_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axid_3_reg;
               (`WR_REQ_DESC_9_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_0_reg;
               (`WR_REQ_DESC_9_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_1_reg;
               (`WR_REQ_DESC_9_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_2_reg;
               (`WR_REQ_DESC_9_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_3_reg;
               (`WR_REQ_DESC_9_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_4_reg;
               (`WR_REQ_DESC_9_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_5_reg;
               (`WR_REQ_DESC_9_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_6_reg;
               (`WR_REQ_DESC_9_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_7_reg;
               (`WR_REQ_DESC_9_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_8_reg;
               (`WR_REQ_DESC_9_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_9_reg;
               (`WR_REQ_DESC_9_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_10_reg;
               (`WR_REQ_DESC_9_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_11_reg;
               (`WR_REQ_DESC_9_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_12_reg;
               (`WR_REQ_DESC_9_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_13_reg;
               (`WR_REQ_DESC_9_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_14_reg;
               (`WR_REQ_DESC_9_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_axuser_15_reg;
               (`WR_REQ_DESC_9_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_0_reg;
               (`WR_REQ_DESC_9_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_1_reg;
               (`WR_REQ_DESC_9_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_2_reg;
               (`WR_REQ_DESC_9_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_3_reg;
               (`WR_REQ_DESC_9_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_4_reg;
               (`WR_REQ_DESC_9_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_5_reg;
               (`WR_REQ_DESC_9_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_6_reg;
               (`WR_REQ_DESC_9_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_7_reg;
               (`WR_REQ_DESC_9_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_8_reg;
               (`WR_REQ_DESC_9_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_9_reg;
               (`WR_REQ_DESC_9_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_10_reg;
               (`WR_REQ_DESC_9_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_11_reg;
               (`WR_REQ_DESC_9_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_12_reg;
               (`WR_REQ_DESC_9_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_13_reg;
               (`WR_REQ_DESC_9_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_14_reg;
               (`WR_REQ_DESC_9_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_9 <= wr_req_desc_9_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_9 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_a <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_A_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_txn_type_reg;
               (`WR_REQ_DESC_A_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_size_reg;
               (`WR_REQ_DESC_A_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_data_offset_reg;
               (`WR_REQ_DESC_A_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_data_host_addr_0_reg;
               (`WR_REQ_DESC_A_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_data_host_addr_1_reg;
               (`WR_REQ_DESC_A_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_data_host_addr_2_reg;
               (`WR_REQ_DESC_A_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_data_host_addr_3_reg;
               (`WR_REQ_DESC_A_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_A_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_A_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_A_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_A_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axsize_reg;
               (`WR_REQ_DESC_A_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_attr_reg;
               (`WR_REQ_DESC_A_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axaddr_0_reg;
               (`WR_REQ_DESC_A_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axaddr_1_reg;
               (`WR_REQ_DESC_A_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axaddr_2_reg;
               (`WR_REQ_DESC_A_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axaddr_3_reg;
               (`WR_REQ_DESC_A_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axid_0_reg;
               (`WR_REQ_DESC_A_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axid_1_reg;
               (`WR_REQ_DESC_A_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axid_2_reg;
               (`WR_REQ_DESC_A_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axid_3_reg;
               (`WR_REQ_DESC_A_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_0_reg;
               (`WR_REQ_DESC_A_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_1_reg;
               (`WR_REQ_DESC_A_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_2_reg;
               (`WR_REQ_DESC_A_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_3_reg;
               (`WR_REQ_DESC_A_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_4_reg;
               (`WR_REQ_DESC_A_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_5_reg;
               (`WR_REQ_DESC_A_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_6_reg;
               (`WR_REQ_DESC_A_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_7_reg;
               (`WR_REQ_DESC_A_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_8_reg;
               (`WR_REQ_DESC_A_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_9_reg;
               (`WR_REQ_DESC_A_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_10_reg;
               (`WR_REQ_DESC_A_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_11_reg;
               (`WR_REQ_DESC_A_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_12_reg;
               (`WR_REQ_DESC_A_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_13_reg;
               (`WR_REQ_DESC_A_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_14_reg;
               (`WR_REQ_DESC_A_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_axuser_15_reg;
               (`WR_REQ_DESC_A_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_0_reg;
               (`WR_REQ_DESC_A_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_1_reg;
               (`WR_REQ_DESC_A_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_2_reg;
               (`WR_REQ_DESC_A_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_3_reg;
               (`WR_REQ_DESC_A_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_4_reg;
               (`WR_REQ_DESC_A_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_5_reg;
               (`WR_REQ_DESC_A_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_6_reg;
               (`WR_REQ_DESC_A_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_7_reg;
               (`WR_REQ_DESC_A_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_8_reg;
               (`WR_REQ_DESC_A_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_9_reg;
               (`WR_REQ_DESC_A_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_10_reg;
               (`WR_REQ_DESC_A_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_11_reg;
               (`WR_REQ_DESC_A_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_12_reg;
               (`WR_REQ_DESC_A_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_13_reg;
               (`WR_REQ_DESC_A_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_14_reg;
               (`WR_REQ_DESC_A_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_a <= wr_req_desc_a_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_a <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_b <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_B_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_txn_type_reg;
               (`WR_REQ_DESC_B_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_size_reg;
               (`WR_REQ_DESC_B_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_data_offset_reg;
               (`WR_REQ_DESC_B_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_data_host_addr_0_reg;
               (`WR_REQ_DESC_B_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_data_host_addr_1_reg;
               (`WR_REQ_DESC_B_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_data_host_addr_2_reg;
               (`WR_REQ_DESC_B_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_data_host_addr_3_reg;
               (`WR_REQ_DESC_B_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_B_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_B_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_B_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_B_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axsize_reg;
               (`WR_REQ_DESC_B_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_attr_reg;
               (`WR_REQ_DESC_B_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axaddr_0_reg;
               (`WR_REQ_DESC_B_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axaddr_1_reg;
               (`WR_REQ_DESC_B_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axaddr_2_reg;
               (`WR_REQ_DESC_B_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axaddr_3_reg;
               (`WR_REQ_DESC_B_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axid_0_reg;
               (`WR_REQ_DESC_B_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axid_1_reg;
               (`WR_REQ_DESC_B_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axid_2_reg;
               (`WR_REQ_DESC_B_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axid_3_reg;
               (`WR_REQ_DESC_B_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_0_reg;
               (`WR_REQ_DESC_B_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_1_reg;
               (`WR_REQ_DESC_B_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_2_reg;
               (`WR_REQ_DESC_B_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_3_reg;
               (`WR_REQ_DESC_B_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_4_reg;
               (`WR_REQ_DESC_B_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_5_reg;
               (`WR_REQ_DESC_B_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_6_reg;
               (`WR_REQ_DESC_B_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_7_reg;
               (`WR_REQ_DESC_B_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_8_reg;
               (`WR_REQ_DESC_B_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_9_reg;
               (`WR_REQ_DESC_B_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_10_reg;
               (`WR_REQ_DESC_B_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_11_reg;
               (`WR_REQ_DESC_B_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_12_reg;
               (`WR_REQ_DESC_B_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_13_reg;
               (`WR_REQ_DESC_B_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_14_reg;
               (`WR_REQ_DESC_B_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_axuser_15_reg;
               (`WR_REQ_DESC_B_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_0_reg;
               (`WR_REQ_DESC_B_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_1_reg;
               (`WR_REQ_DESC_B_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_2_reg;
               (`WR_REQ_DESC_B_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_3_reg;
               (`WR_REQ_DESC_B_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_4_reg;
               (`WR_REQ_DESC_B_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_5_reg;
               (`WR_REQ_DESC_B_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_6_reg;
               (`WR_REQ_DESC_B_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_7_reg;
               (`WR_REQ_DESC_B_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_8_reg;
               (`WR_REQ_DESC_B_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_9_reg;
               (`WR_REQ_DESC_B_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_10_reg;
               (`WR_REQ_DESC_B_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_11_reg;
               (`WR_REQ_DESC_B_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_12_reg;
               (`WR_REQ_DESC_B_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_13_reg;
               (`WR_REQ_DESC_B_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_14_reg;
               (`WR_REQ_DESC_B_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_b <= wr_req_desc_b_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_b <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_c <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_C_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_txn_type_reg;
               (`WR_REQ_DESC_C_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_size_reg;
               (`WR_REQ_DESC_C_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_data_offset_reg;
               (`WR_REQ_DESC_C_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_data_host_addr_0_reg;
               (`WR_REQ_DESC_C_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_data_host_addr_1_reg;
               (`WR_REQ_DESC_C_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_data_host_addr_2_reg;
               (`WR_REQ_DESC_C_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_data_host_addr_3_reg;
               (`WR_REQ_DESC_C_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_C_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_C_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_C_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_C_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axsize_reg;
               (`WR_REQ_DESC_C_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_attr_reg;
               (`WR_REQ_DESC_C_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axaddr_0_reg;
               (`WR_REQ_DESC_C_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axaddr_1_reg;
               (`WR_REQ_DESC_C_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axaddr_2_reg;
               (`WR_REQ_DESC_C_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axaddr_3_reg;
               (`WR_REQ_DESC_C_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axid_0_reg;
               (`WR_REQ_DESC_C_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axid_1_reg;
               (`WR_REQ_DESC_C_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axid_2_reg;
               (`WR_REQ_DESC_C_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axid_3_reg;
               (`WR_REQ_DESC_C_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_0_reg;
               (`WR_REQ_DESC_C_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_1_reg;
               (`WR_REQ_DESC_C_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_2_reg;
               (`WR_REQ_DESC_C_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_3_reg;
               (`WR_REQ_DESC_C_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_4_reg;
               (`WR_REQ_DESC_C_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_5_reg;
               (`WR_REQ_DESC_C_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_6_reg;
               (`WR_REQ_DESC_C_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_7_reg;
               (`WR_REQ_DESC_C_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_8_reg;
               (`WR_REQ_DESC_C_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_9_reg;
               (`WR_REQ_DESC_C_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_10_reg;
               (`WR_REQ_DESC_C_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_11_reg;
               (`WR_REQ_DESC_C_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_12_reg;
               (`WR_REQ_DESC_C_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_13_reg;
               (`WR_REQ_DESC_C_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_14_reg;
               (`WR_REQ_DESC_C_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_axuser_15_reg;
               (`WR_REQ_DESC_C_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_0_reg;
               (`WR_REQ_DESC_C_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_1_reg;
               (`WR_REQ_DESC_C_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_2_reg;
               (`WR_REQ_DESC_C_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_3_reg;
               (`WR_REQ_DESC_C_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_4_reg;
               (`WR_REQ_DESC_C_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_5_reg;
               (`WR_REQ_DESC_C_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_6_reg;
               (`WR_REQ_DESC_C_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_7_reg;
               (`WR_REQ_DESC_C_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_8_reg;
               (`WR_REQ_DESC_C_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_9_reg;
               (`WR_REQ_DESC_C_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_10_reg;
               (`WR_REQ_DESC_C_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_11_reg;
               (`WR_REQ_DESC_C_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_12_reg;
               (`WR_REQ_DESC_C_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_13_reg;
               (`WR_REQ_DESC_C_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_14_reg;
               (`WR_REQ_DESC_C_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_c <= wr_req_desc_c_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_c <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_d <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_D_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_txn_type_reg;
               (`WR_REQ_DESC_D_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_size_reg;
               (`WR_REQ_DESC_D_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_data_offset_reg;
               (`WR_REQ_DESC_D_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_data_host_addr_0_reg;
               (`WR_REQ_DESC_D_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_data_host_addr_1_reg;
               (`WR_REQ_DESC_D_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_data_host_addr_2_reg;
               (`WR_REQ_DESC_D_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_data_host_addr_3_reg;
               (`WR_REQ_DESC_D_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_D_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_D_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_D_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_D_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axsize_reg;
               (`WR_REQ_DESC_D_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_attr_reg;
               (`WR_REQ_DESC_D_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axaddr_0_reg;
               (`WR_REQ_DESC_D_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axaddr_1_reg;
               (`WR_REQ_DESC_D_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axaddr_2_reg;
               (`WR_REQ_DESC_D_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axaddr_3_reg;
               (`WR_REQ_DESC_D_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axid_0_reg;
               (`WR_REQ_DESC_D_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axid_1_reg;
               (`WR_REQ_DESC_D_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axid_2_reg;
               (`WR_REQ_DESC_D_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axid_3_reg;
               (`WR_REQ_DESC_D_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_0_reg;
               (`WR_REQ_DESC_D_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_1_reg;
               (`WR_REQ_DESC_D_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_2_reg;
               (`WR_REQ_DESC_D_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_3_reg;
               (`WR_REQ_DESC_D_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_4_reg;
               (`WR_REQ_DESC_D_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_5_reg;
               (`WR_REQ_DESC_D_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_6_reg;
               (`WR_REQ_DESC_D_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_7_reg;
               (`WR_REQ_DESC_D_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_8_reg;
               (`WR_REQ_DESC_D_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_9_reg;
               (`WR_REQ_DESC_D_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_10_reg;
               (`WR_REQ_DESC_D_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_11_reg;
               (`WR_REQ_DESC_D_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_12_reg;
               (`WR_REQ_DESC_D_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_13_reg;
               (`WR_REQ_DESC_D_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_14_reg;
               (`WR_REQ_DESC_D_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_axuser_15_reg;
               (`WR_REQ_DESC_D_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_0_reg;
               (`WR_REQ_DESC_D_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_1_reg;
               (`WR_REQ_DESC_D_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_2_reg;
               (`WR_REQ_DESC_D_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_3_reg;
               (`WR_REQ_DESC_D_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_4_reg;
               (`WR_REQ_DESC_D_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_5_reg;
               (`WR_REQ_DESC_D_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_6_reg;
               (`WR_REQ_DESC_D_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_7_reg;
               (`WR_REQ_DESC_D_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_8_reg;
               (`WR_REQ_DESC_D_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_9_reg;
               (`WR_REQ_DESC_D_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_10_reg;
               (`WR_REQ_DESC_D_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_11_reg;
               (`WR_REQ_DESC_D_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_12_reg;
               (`WR_REQ_DESC_D_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_13_reg;
               (`WR_REQ_DESC_D_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_14_reg;
               (`WR_REQ_DESC_D_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_d <= wr_req_desc_d_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_d <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_e <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_E_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_txn_type_reg;
               (`WR_REQ_DESC_E_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_size_reg;
               (`WR_REQ_DESC_E_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_data_offset_reg;
               (`WR_REQ_DESC_E_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_data_host_addr_0_reg;
               (`WR_REQ_DESC_E_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_data_host_addr_1_reg;
               (`WR_REQ_DESC_E_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_data_host_addr_2_reg;
               (`WR_REQ_DESC_E_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_data_host_addr_3_reg;
               (`WR_REQ_DESC_E_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_E_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_E_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_E_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_E_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axsize_reg;
               (`WR_REQ_DESC_E_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_attr_reg;
               (`WR_REQ_DESC_E_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axaddr_0_reg;
               (`WR_REQ_DESC_E_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axaddr_1_reg;
               (`WR_REQ_DESC_E_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axaddr_2_reg;
               (`WR_REQ_DESC_E_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axaddr_3_reg;
               (`WR_REQ_DESC_E_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axid_0_reg;
               (`WR_REQ_DESC_E_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axid_1_reg;
               (`WR_REQ_DESC_E_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axid_2_reg;
               (`WR_REQ_DESC_E_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axid_3_reg;
               (`WR_REQ_DESC_E_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_0_reg;
               (`WR_REQ_DESC_E_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_1_reg;
               (`WR_REQ_DESC_E_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_2_reg;
               (`WR_REQ_DESC_E_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_3_reg;
               (`WR_REQ_DESC_E_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_4_reg;
               (`WR_REQ_DESC_E_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_5_reg;
               (`WR_REQ_DESC_E_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_6_reg;
               (`WR_REQ_DESC_E_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_7_reg;
               (`WR_REQ_DESC_E_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_8_reg;
               (`WR_REQ_DESC_E_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_9_reg;
               (`WR_REQ_DESC_E_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_10_reg;
               (`WR_REQ_DESC_E_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_11_reg;
               (`WR_REQ_DESC_E_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_12_reg;
               (`WR_REQ_DESC_E_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_13_reg;
               (`WR_REQ_DESC_E_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_14_reg;
               (`WR_REQ_DESC_E_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_axuser_15_reg;
               (`WR_REQ_DESC_E_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_0_reg;
               (`WR_REQ_DESC_E_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_1_reg;
               (`WR_REQ_DESC_E_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_2_reg;
               (`WR_REQ_DESC_E_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_3_reg;
               (`WR_REQ_DESC_E_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_4_reg;
               (`WR_REQ_DESC_E_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_5_reg;
               (`WR_REQ_DESC_E_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_6_reg;
               (`WR_REQ_DESC_E_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_7_reg;
               (`WR_REQ_DESC_E_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_8_reg;
               (`WR_REQ_DESC_E_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_9_reg;
               (`WR_REQ_DESC_E_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_10_reg;
               (`WR_REQ_DESC_E_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_11_reg;
               (`WR_REQ_DESC_E_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_12_reg;
               (`WR_REQ_DESC_E_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_13_reg;
               (`WR_REQ_DESC_E_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_14_reg;
               (`WR_REQ_DESC_E_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_e <= wr_req_desc_e_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_e <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_req_desc_f <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_REQ_DESC_F_TXN_TYPE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_txn_type_reg;
               (`WR_REQ_DESC_F_SIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_size_reg;
               (`WR_REQ_DESC_F_DATA_OFFSET_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_data_offset_reg;
               (`WR_REQ_DESC_F_DATA_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_data_host_addr_0_reg;
               (`WR_REQ_DESC_F_DATA_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_data_host_addr_1_reg;
               (`WR_REQ_DESC_F_DATA_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_data_host_addr_2_reg;
               (`WR_REQ_DESC_F_DATA_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_data_host_addr_3_reg;
               (`WR_REQ_DESC_F_WSTRB_HOST_ADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wstrb_host_addr_0_reg;
               (`WR_REQ_DESC_F_WSTRB_HOST_ADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wstrb_host_addr_1_reg;
               (`WR_REQ_DESC_F_WSTRB_HOST_ADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wstrb_host_addr_2_reg;
               (`WR_REQ_DESC_F_WSTRB_HOST_ADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wstrb_host_addr_3_reg;
               (`WR_REQ_DESC_F_AXSIZE_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axsize_reg;
               (`WR_REQ_DESC_F_ATTR_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_attr_reg;
               (`WR_REQ_DESC_F_AXADDR_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axaddr_0_reg;
               (`WR_REQ_DESC_F_AXADDR_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axaddr_1_reg;
               (`WR_REQ_DESC_F_AXADDR_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axaddr_2_reg;
               (`WR_REQ_DESC_F_AXADDR_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axaddr_3_reg;
               (`WR_REQ_DESC_F_AXID_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axid_0_reg;
               (`WR_REQ_DESC_F_AXID_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axid_1_reg;
               (`WR_REQ_DESC_F_AXID_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axid_2_reg;
               (`WR_REQ_DESC_F_AXID_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axid_3_reg;
               (`WR_REQ_DESC_F_AXUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_0_reg;
               (`WR_REQ_DESC_F_AXUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_1_reg;
               (`WR_REQ_DESC_F_AXUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_2_reg;
               (`WR_REQ_DESC_F_AXUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_3_reg;
               (`WR_REQ_DESC_F_AXUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_4_reg;
               (`WR_REQ_DESC_F_AXUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_5_reg;
               (`WR_REQ_DESC_F_AXUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_6_reg;
               (`WR_REQ_DESC_F_AXUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_7_reg;
               (`WR_REQ_DESC_F_AXUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_8_reg;
               (`WR_REQ_DESC_F_AXUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_9_reg;
               (`WR_REQ_DESC_F_AXUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_10_reg;
               (`WR_REQ_DESC_F_AXUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_11_reg;
               (`WR_REQ_DESC_F_AXUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_12_reg;
               (`WR_REQ_DESC_F_AXUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_13_reg;
               (`WR_REQ_DESC_F_AXUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_14_reg;
               (`WR_REQ_DESC_F_AXUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_axuser_15_reg;
               (`WR_REQ_DESC_F_WUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_0_reg;
               (`WR_REQ_DESC_F_WUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_1_reg;
               (`WR_REQ_DESC_F_WUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_2_reg;
               (`WR_REQ_DESC_F_WUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_3_reg;
               (`WR_REQ_DESC_F_WUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_4_reg;
               (`WR_REQ_DESC_F_WUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_5_reg;
               (`WR_REQ_DESC_F_WUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_6_reg;
               (`WR_REQ_DESC_F_WUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_7_reg;
               (`WR_REQ_DESC_F_WUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_8_reg;
               (`WR_REQ_DESC_F_WUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_9_reg;
               (`WR_REQ_DESC_F_WUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_10_reg;
               (`WR_REQ_DESC_F_WUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_11_reg;
               (`WR_REQ_DESC_F_WUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_12_reg;
               (`WR_REQ_DESC_F_WUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_13_reg;
               (`WR_REQ_DESC_F_WUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_14_reg;
               (`WR_REQ_DESC_F_WUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_req_desc_f <= wr_req_desc_f_wuser_15_reg;
               default                                  :reg_data_out_wr_req_desc_f <= 32'b0      ;        
             endcase
	  end
     end




   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_0 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_0_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_resp_reg;
               (`WR_RESP_DESC_0_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xid_0_reg;
               (`WR_RESP_DESC_0_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xid_1_reg;
               (`WR_RESP_DESC_0_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xid_2_reg;
               (`WR_RESP_DESC_0_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xid_3_reg;
               (`WR_RESP_DESC_0_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_0_reg;
               (`WR_RESP_DESC_0_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_1_reg;
               (`WR_RESP_DESC_0_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_2_reg;
               (`WR_RESP_DESC_0_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_3_reg;
               (`WR_RESP_DESC_0_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_4_reg;
               (`WR_RESP_DESC_0_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_5_reg;
               (`WR_RESP_DESC_0_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_6_reg;
               (`WR_RESP_DESC_0_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_7_reg;
               (`WR_RESP_DESC_0_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_8_reg;
               (`WR_RESP_DESC_0_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_9_reg;
               (`WR_RESP_DESC_0_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_10_reg;
               (`WR_RESP_DESC_0_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_11_reg;
               (`WR_RESP_DESC_0_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_12_reg;
               (`WR_RESP_DESC_0_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_13_reg;
               (`WR_RESP_DESC_0_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_14_reg;
               (`WR_RESP_DESC_0_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_0 <= wr_resp_desc_0_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_0 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_1 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_1_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_resp_reg;
               (`WR_RESP_DESC_1_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xid_0_reg;
               (`WR_RESP_DESC_1_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xid_1_reg;
               (`WR_RESP_DESC_1_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xid_2_reg;
               (`WR_RESP_DESC_1_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xid_3_reg;
               (`WR_RESP_DESC_1_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_0_reg;
               (`WR_RESP_DESC_1_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_1_reg;
               (`WR_RESP_DESC_1_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_2_reg;
               (`WR_RESP_DESC_1_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_3_reg;
               (`WR_RESP_DESC_1_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_4_reg;
               (`WR_RESP_DESC_1_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_5_reg;
               (`WR_RESP_DESC_1_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_6_reg;
               (`WR_RESP_DESC_1_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_7_reg;
               (`WR_RESP_DESC_1_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_8_reg;
               (`WR_RESP_DESC_1_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_9_reg;
               (`WR_RESP_DESC_1_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_10_reg;
               (`WR_RESP_DESC_1_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_11_reg;
               (`WR_RESP_DESC_1_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_12_reg;
               (`WR_RESP_DESC_1_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_13_reg;
               (`WR_RESP_DESC_1_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_14_reg;
               (`WR_RESP_DESC_1_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_1 <= wr_resp_desc_1_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_1 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_2 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_2_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_resp_reg;
               (`WR_RESP_DESC_2_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xid_0_reg;
               (`WR_RESP_DESC_2_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xid_1_reg;
               (`WR_RESP_DESC_2_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xid_2_reg;
               (`WR_RESP_DESC_2_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xid_3_reg;
               (`WR_RESP_DESC_2_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_0_reg;
               (`WR_RESP_DESC_2_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_1_reg;
               (`WR_RESP_DESC_2_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_2_reg;
               (`WR_RESP_DESC_2_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_3_reg;
               (`WR_RESP_DESC_2_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_4_reg;
               (`WR_RESP_DESC_2_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_5_reg;
               (`WR_RESP_DESC_2_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_6_reg;
               (`WR_RESP_DESC_2_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_7_reg;
               (`WR_RESP_DESC_2_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_8_reg;
               (`WR_RESP_DESC_2_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_9_reg;
               (`WR_RESP_DESC_2_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_10_reg;
               (`WR_RESP_DESC_2_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_11_reg;
               (`WR_RESP_DESC_2_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_12_reg;
               (`WR_RESP_DESC_2_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_13_reg;
               (`WR_RESP_DESC_2_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_14_reg;
               (`WR_RESP_DESC_2_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_2 <= wr_resp_desc_2_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_2 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_3 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_3_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_resp_reg;
               (`WR_RESP_DESC_3_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xid_0_reg;
               (`WR_RESP_DESC_3_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xid_1_reg;
               (`WR_RESP_DESC_3_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xid_2_reg;
               (`WR_RESP_DESC_3_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xid_3_reg;
               (`WR_RESP_DESC_3_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_0_reg;
               (`WR_RESP_DESC_3_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_1_reg;
               (`WR_RESP_DESC_3_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_2_reg;
               (`WR_RESP_DESC_3_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_3_reg;
               (`WR_RESP_DESC_3_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_4_reg;
               (`WR_RESP_DESC_3_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_5_reg;
               (`WR_RESP_DESC_3_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_6_reg;
               (`WR_RESP_DESC_3_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_7_reg;
               (`WR_RESP_DESC_3_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_8_reg;
               (`WR_RESP_DESC_3_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_9_reg;
               (`WR_RESP_DESC_3_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_10_reg;
               (`WR_RESP_DESC_3_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_11_reg;
               (`WR_RESP_DESC_3_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_12_reg;
               (`WR_RESP_DESC_3_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_13_reg;
               (`WR_RESP_DESC_3_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_14_reg;
               (`WR_RESP_DESC_3_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_3 <= wr_resp_desc_3_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_3 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_4 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_4_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_resp_reg;
               (`WR_RESP_DESC_4_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xid_0_reg;
               (`WR_RESP_DESC_4_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xid_1_reg;
               (`WR_RESP_DESC_4_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xid_2_reg;
               (`WR_RESP_DESC_4_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xid_3_reg;
               (`WR_RESP_DESC_4_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_0_reg;
               (`WR_RESP_DESC_4_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_1_reg;
               (`WR_RESP_DESC_4_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_2_reg;
               (`WR_RESP_DESC_4_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_3_reg;
               (`WR_RESP_DESC_4_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_4_reg;
               (`WR_RESP_DESC_4_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_5_reg;
               (`WR_RESP_DESC_4_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_6_reg;
               (`WR_RESP_DESC_4_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_7_reg;
               (`WR_RESP_DESC_4_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_8_reg;
               (`WR_RESP_DESC_4_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_9_reg;
               (`WR_RESP_DESC_4_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_10_reg;
               (`WR_RESP_DESC_4_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_11_reg;
               (`WR_RESP_DESC_4_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_12_reg;
               (`WR_RESP_DESC_4_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_13_reg;
               (`WR_RESP_DESC_4_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_14_reg;
               (`WR_RESP_DESC_4_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_4 <= wr_resp_desc_4_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_4 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_5 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_5_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_resp_reg;
               (`WR_RESP_DESC_5_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xid_0_reg;
               (`WR_RESP_DESC_5_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xid_1_reg;
               (`WR_RESP_DESC_5_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xid_2_reg;
               (`WR_RESP_DESC_5_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xid_3_reg;
               (`WR_RESP_DESC_5_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_0_reg;
               (`WR_RESP_DESC_5_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_1_reg;
               (`WR_RESP_DESC_5_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_2_reg;
               (`WR_RESP_DESC_5_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_3_reg;
               (`WR_RESP_DESC_5_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_4_reg;
               (`WR_RESP_DESC_5_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_5_reg;
               (`WR_RESP_DESC_5_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_6_reg;
               (`WR_RESP_DESC_5_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_7_reg;
               (`WR_RESP_DESC_5_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_8_reg;
               (`WR_RESP_DESC_5_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_9_reg;
               (`WR_RESP_DESC_5_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_10_reg;
               (`WR_RESP_DESC_5_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_11_reg;
               (`WR_RESP_DESC_5_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_12_reg;
               (`WR_RESP_DESC_5_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_13_reg;
               (`WR_RESP_DESC_5_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_14_reg;
               (`WR_RESP_DESC_5_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_5 <= wr_resp_desc_5_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_5 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_6 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_6_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_resp_reg;
               (`WR_RESP_DESC_6_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xid_0_reg;
               (`WR_RESP_DESC_6_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xid_1_reg;
               (`WR_RESP_DESC_6_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xid_2_reg;
               (`WR_RESP_DESC_6_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xid_3_reg;
               (`WR_RESP_DESC_6_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_0_reg;
               (`WR_RESP_DESC_6_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_1_reg;
               (`WR_RESP_DESC_6_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_2_reg;
               (`WR_RESP_DESC_6_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_3_reg;
               (`WR_RESP_DESC_6_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_4_reg;
               (`WR_RESP_DESC_6_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_5_reg;
               (`WR_RESP_DESC_6_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_6_reg;
               (`WR_RESP_DESC_6_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_7_reg;
               (`WR_RESP_DESC_6_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_8_reg;
               (`WR_RESP_DESC_6_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_9_reg;
               (`WR_RESP_DESC_6_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_10_reg;
               (`WR_RESP_DESC_6_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_11_reg;
               (`WR_RESP_DESC_6_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_12_reg;
               (`WR_RESP_DESC_6_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_13_reg;
               (`WR_RESP_DESC_6_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_14_reg;
               (`WR_RESP_DESC_6_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_6 <= wr_resp_desc_6_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_6 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_7 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_7_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_resp_reg;
               (`WR_RESP_DESC_7_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xid_0_reg;
               (`WR_RESP_DESC_7_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xid_1_reg;
               (`WR_RESP_DESC_7_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xid_2_reg;
               (`WR_RESP_DESC_7_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xid_3_reg;
               (`WR_RESP_DESC_7_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_0_reg;
               (`WR_RESP_DESC_7_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_1_reg;
               (`WR_RESP_DESC_7_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_2_reg;
               (`WR_RESP_DESC_7_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_3_reg;
               (`WR_RESP_DESC_7_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_4_reg;
               (`WR_RESP_DESC_7_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_5_reg;
               (`WR_RESP_DESC_7_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_6_reg;
               (`WR_RESP_DESC_7_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_7_reg;
               (`WR_RESP_DESC_7_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_8_reg;
               (`WR_RESP_DESC_7_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_9_reg;
               (`WR_RESP_DESC_7_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_10_reg;
               (`WR_RESP_DESC_7_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_11_reg;
               (`WR_RESP_DESC_7_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_12_reg;
               (`WR_RESP_DESC_7_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_13_reg;
               (`WR_RESP_DESC_7_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_14_reg;
               (`WR_RESP_DESC_7_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_7 <= wr_resp_desc_7_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_7 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_8 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_8_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_resp_reg;
               (`WR_RESP_DESC_8_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xid_0_reg;
               (`WR_RESP_DESC_8_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xid_1_reg;
               (`WR_RESP_DESC_8_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xid_2_reg;
               (`WR_RESP_DESC_8_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xid_3_reg;
               (`WR_RESP_DESC_8_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_0_reg;
               (`WR_RESP_DESC_8_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_1_reg;
               (`WR_RESP_DESC_8_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_2_reg;
               (`WR_RESP_DESC_8_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_3_reg;
               (`WR_RESP_DESC_8_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_4_reg;
               (`WR_RESP_DESC_8_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_5_reg;
               (`WR_RESP_DESC_8_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_6_reg;
               (`WR_RESP_DESC_8_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_7_reg;
               (`WR_RESP_DESC_8_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_8_reg;
               (`WR_RESP_DESC_8_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_9_reg;
               (`WR_RESP_DESC_8_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_10_reg;
               (`WR_RESP_DESC_8_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_11_reg;
               (`WR_RESP_DESC_8_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_12_reg;
               (`WR_RESP_DESC_8_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_13_reg;
               (`WR_RESP_DESC_8_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_14_reg;
               (`WR_RESP_DESC_8_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_8 <= wr_resp_desc_8_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_8 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_9 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_9_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_resp_reg;
               (`WR_RESP_DESC_9_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xid_0_reg;
               (`WR_RESP_DESC_9_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xid_1_reg;
               (`WR_RESP_DESC_9_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xid_2_reg;
               (`WR_RESP_DESC_9_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xid_3_reg;
               (`WR_RESP_DESC_9_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_0_reg;
               (`WR_RESP_DESC_9_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_1_reg;
               (`WR_RESP_DESC_9_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_2_reg;
               (`WR_RESP_DESC_9_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_3_reg;
               (`WR_RESP_DESC_9_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_4_reg;
               (`WR_RESP_DESC_9_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_5_reg;
               (`WR_RESP_DESC_9_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_6_reg;
               (`WR_RESP_DESC_9_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_7_reg;
               (`WR_RESP_DESC_9_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_8_reg;
               (`WR_RESP_DESC_9_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_9_reg;
               (`WR_RESP_DESC_9_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_10_reg;
               (`WR_RESP_DESC_9_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_11_reg;
               (`WR_RESP_DESC_9_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_12_reg;
               (`WR_RESP_DESC_9_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_13_reg;
               (`WR_RESP_DESC_9_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_14_reg;
               (`WR_RESP_DESC_9_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_9 <= wr_resp_desc_9_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_9 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_a <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_A_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_resp_reg;
               (`WR_RESP_DESC_A_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xid_0_reg;
               (`WR_RESP_DESC_A_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xid_1_reg;
               (`WR_RESP_DESC_A_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xid_2_reg;
               (`WR_RESP_DESC_A_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xid_3_reg;
               (`WR_RESP_DESC_A_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_0_reg;
               (`WR_RESP_DESC_A_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_1_reg;
               (`WR_RESP_DESC_A_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_2_reg;
               (`WR_RESP_DESC_A_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_3_reg;
               (`WR_RESP_DESC_A_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_4_reg;
               (`WR_RESP_DESC_A_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_5_reg;
               (`WR_RESP_DESC_A_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_6_reg;
               (`WR_RESP_DESC_A_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_7_reg;
               (`WR_RESP_DESC_A_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_8_reg;
               (`WR_RESP_DESC_A_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_9_reg;
               (`WR_RESP_DESC_A_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_10_reg;
               (`WR_RESP_DESC_A_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_11_reg;
               (`WR_RESP_DESC_A_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_12_reg;
               (`WR_RESP_DESC_A_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_13_reg;
               (`WR_RESP_DESC_A_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_14_reg;
               (`WR_RESP_DESC_A_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_a <= wr_resp_desc_a_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_a <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_b <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_B_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_resp_reg;
               (`WR_RESP_DESC_B_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xid_0_reg;
               (`WR_RESP_DESC_B_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xid_1_reg;
               (`WR_RESP_DESC_B_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xid_2_reg;
               (`WR_RESP_DESC_B_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xid_3_reg;
               (`WR_RESP_DESC_B_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_0_reg;
               (`WR_RESP_DESC_B_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_1_reg;
               (`WR_RESP_DESC_B_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_2_reg;
               (`WR_RESP_DESC_B_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_3_reg;
               (`WR_RESP_DESC_B_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_4_reg;
               (`WR_RESP_DESC_B_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_5_reg;
               (`WR_RESP_DESC_B_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_6_reg;
               (`WR_RESP_DESC_B_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_7_reg;
               (`WR_RESP_DESC_B_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_8_reg;
               (`WR_RESP_DESC_B_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_9_reg;
               (`WR_RESP_DESC_B_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_10_reg;
               (`WR_RESP_DESC_B_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_11_reg;
               (`WR_RESP_DESC_B_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_12_reg;
               (`WR_RESP_DESC_B_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_13_reg;
               (`WR_RESP_DESC_B_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_14_reg;
               (`WR_RESP_DESC_B_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_b <= wr_resp_desc_b_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_b <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_c <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_C_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_resp_reg;
               (`WR_RESP_DESC_C_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xid_0_reg;
               (`WR_RESP_DESC_C_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xid_1_reg;
               (`WR_RESP_DESC_C_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xid_2_reg;
               (`WR_RESP_DESC_C_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xid_3_reg;
               (`WR_RESP_DESC_C_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_0_reg;
               (`WR_RESP_DESC_C_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_1_reg;
               (`WR_RESP_DESC_C_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_2_reg;
               (`WR_RESP_DESC_C_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_3_reg;
               (`WR_RESP_DESC_C_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_4_reg;
               (`WR_RESP_DESC_C_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_5_reg;
               (`WR_RESP_DESC_C_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_6_reg;
               (`WR_RESP_DESC_C_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_7_reg;
               (`WR_RESP_DESC_C_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_8_reg;
               (`WR_RESP_DESC_C_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_9_reg;
               (`WR_RESP_DESC_C_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_10_reg;
               (`WR_RESP_DESC_C_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_11_reg;
               (`WR_RESP_DESC_C_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_12_reg;
               (`WR_RESP_DESC_C_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_13_reg;
               (`WR_RESP_DESC_C_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_14_reg;
               (`WR_RESP_DESC_C_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_c <= wr_resp_desc_c_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_c <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_d <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_D_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_resp_reg;
               (`WR_RESP_DESC_D_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xid_0_reg;
               (`WR_RESP_DESC_D_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xid_1_reg;
               (`WR_RESP_DESC_D_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xid_2_reg;
               (`WR_RESP_DESC_D_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xid_3_reg;
               (`WR_RESP_DESC_D_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_0_reg;
               (`WR_RESP_DESC_D_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_1_reg;
               (`WR_RESP_DESC_D_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_2_reg;
               (`WR_RESP_DESC_D_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_3_reg;
               (`WR_RESP_DESC_D_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_4_reg;
               (`WR_RESP_DESC_D_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_5_reg;
               (`WR_RESP_DESC_D_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_6_reg;
               (`WR_RESP_DESC_D_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_7_reg;
               (`WR_RESP_DESC_D_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_8_reg;
               (`WR_RESP_DESC_D_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_9_reg;
               (`WR_RESP_DESC_D_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_10_reg;
               (`WR_RESP_DESC_D_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_11_reg;
               (`WR_RESP_DESC_D_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_12_reg;
               (`WR_RESP_DESC_D_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_13_reg;
               (`WR_RESP_DESC_D_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_14_reg;
               (`WR_RESP_DESC_D_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_d <= wr_resp_desc_d_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_d <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_e <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_E_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_resp_reg;
               (`WR_RESP_DESC_E_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xid_0_reg;
               (`WR_RESP_DESC_E_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xid_1_reg;
               (`WR_RESP_DESC_E_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xid_2_reg;
               (`WR_RESP_DESC_E_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xid_3_reg;
               (`WR_RESP_DESC_E_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_0_reg;
               (`WR_RESP_DESC_E_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_1_reg;
               (`WR_RESP_DESC_E_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_2_reg;
               (`WR_RESP_DESC_E_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_3_reg;
               (`WR_RESP_DESC_E_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_4_reg;
               (`WR_RESP_DESC_E_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_5_reg;
               (`WR_RESP_DESC_E_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_6_reg;
               (`WR_RESP_DESC_E_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_7_reg;
               (`WR_RESP_DESC_E_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_8_reg;
               (`WR_RESP_DESC_E_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_9_reg;
               (`WR_RESP_DESC_E_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_10_reg;
               (`WR_RESP_DESC_E_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_11_reg;
               (`WR_RESP_DESC_E_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_12_reg;
               (`WR_RESP_DESC_E_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_13_reg;
               (`WR_RESP_DESC_E_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_14_reg;
               (`WR_RESP_DESC_E_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_e <= wr_resp_desc_e_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_e <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_wr_resp_desc_f <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`WR_RESP_DESC_F_RESP_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_resp_reg;
               (`WR_RESP_DESC_F_XID_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xid_0_reg;
               (`WR_RESP_DESC_F_XID_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xid_1_reg;
               (`WR_RESP_DESC_F_XID_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xid_2_reg;
               (`WR_RESP_DESC_F_XID_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xid_3_reg;
               (`WR_RESP_DESC_F_XUSER_0_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_0_reg;
               (`WR_RESP_DESC_F_XUSER_1_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_1_reg;
               (`WR_RESP_DESC_F_XUSER_2_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_2_reg;
               (`WR_RESP_DESC_F_XUSER_3_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_3_reg;
               (`WR_RESP_DESC_F_XUSER_4_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_4_reg;
               (`WR_RESP_DESC_F_XUSER_5_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_5_reg;
               (`WR_RESP_DESC_F_XUSER_6_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_6_reg;
               (`WR_RESP_DESC_F_XUSER_7_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_7_reg;
               (`WR_RESP_DESC_F_XUSER_8_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_8_reg;
               (`WR_RESP_DESC_F_XUSER_9_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_9_reg;
               (`WR_RESP_DESC_F_XUSER_10_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_10_reg;
               (`WR_RESP_DESC_F_XUSER_11_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_11_reg;
               (`WR_RESP_DESC_F_XUSER_12_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_12_reg;
               (`WR_RESP_DESC_F_XUSER_13_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_13_reg;
               (`WR_RESP_DESC_F_XUSER_14_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_14_reg;
               (`WR_RESP_DESC_F_XUSER_15_REG_ADDR&'hFF) :reg_data_out_wr_resp_desc_f <= wr_resp_desc_f_xuser_15_reg;
               default                                  :reg_data_out_wr_resp_desc_f <= 32'b0      ;        
             endcase
	  end
     end




   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_0 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_0_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_0 <= sn_req_desc_0_attr_reg;
               (`SN_REQ_DESC_0_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_0 <= sn_req_desc_0_acaddr_0_reg;
               (`SN_REQ_DESC_0_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_0 <= sn_req_desc_0_acaddr_1_reg;
               (`SN_REQ_DESC_0_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_0 <= sn_req_desc_0_acaddr_2_reg;
               (`SN_REQ_DESC_0_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_0 <= sn_req_desc_0_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_0 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_1 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_1_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_1 <= sn_req_desc_1_attr_reg;
               (`SN_REQ_DESC_1_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_1 <= sn_req_desc_1_acaddr_0_reg;
               (`SN_REQ_DESC_1_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_1 <= sn_req_desc_1_acaddr_1_reg;
               (`SN_REQ_DESC_1_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_1 <= sn_req_desc_1_acaddr_2_reg;
               (`SN_REQ_DESC_1_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_1 <= sn_req_desc_1_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_1 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_2 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_2_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_2 <= sn_req_desc_2_attr_reg;
               (`SN_REQ_DESC_2_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_2 <= sn_req_desc_2_acaddr_0_reg;
               (`SN_REQ_DESC_2_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_2 <= sn_req_desc_2_acaddr_1_reg;
               (`SN_REQ_DESC_2_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_2 <= sn_req_desc_2_acaddr_2_reg;
               (`SN_REQ_DESC_2_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_2 <= sn_req_desc_2_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_2 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_3 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_3_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_3 <= sn_req_desc_3_attr_reg;
               (`SN_REQ_DESC_3_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_3 <= sn_req_desc_3_acaddr_0_reg;
               (`SN_REQ_DESC_3_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_3 <= sn_req_desc_3_acaddr_1_reg;
               (`SN_REQ_DESC_3_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_3 <= sn_req_desc_3_acaddr_2_reg;
               (`SN_REQ_DESC_3_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_3 <= sn_req_desc_3_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_3 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_4 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_4_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_4 <= sn_req_desc_4_attr_reg;
               (`SN_REQ_DESC_4_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_4 <= sn_req_desc_4_acaddr_0_reg;
               (`SN_REQ_DESC_4_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_4 <= sn_req_desc_4_acaddr_1_reg;
               (`SN_REQ_DESC_4_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_4 <= sn_req_desc_4_acaddr_2_reg;
               (`SN_REQ_DESC_4_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_4 <= sn_req_desc_4_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_4 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_5 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_5_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_5 <= sn_req_desc_5_attr_reg;
               (`SN_REQ_DESC_5_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_5 <= sn_req_desc_5_acaddr_0_reg;
               (`SN_REQ_DESC_5_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_5 <= sn_req_desc_5_acaddr_1_reg;
               (`SN_REQ_DESC_5_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_5 <= sn_req_desc_5_acaddr_2_reg;
               (`SN_REQ_DESC_5_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_5 <= sn_req_desc_5_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_5 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_6 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_6_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_6 <= sn_req_desc_6_attr_reg;
               (`SN_REQ_DESC_6_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_6 <= sn_req_desc_6_acaddr_0_reg;
               (`SN_REQ_DESC_6_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_6 <= sn_req_desc_6_acaddr_1_reg;
               (`SN_REQ_DESC_6_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_6 <= sn_req_desc_6_acaddr_2_reg;
               (`SN_REQ_DESC_6_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_6 <= sn_req_desc_6_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_6 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_7 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_7_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_7 <= sn_req_desc_7_attr_reg;
               (`SN_REQ_DESC_7_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_7 <= sn_req_desc_7_acaddr_0_reg;
               (`SN_REQ_DESC_7_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_7 <= sn_req_desc_7_acaddr_1_reg;
               (`SN_REQ_DESC_7_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_7 <= sn_req_desc_7_acaddr_2_reg;
               (`SN_REQ_DESC_7_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_7 <= sn_req_desc_7_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_7 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_8 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_8_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_8 <= sn_req_desc_8_attr_reg;
               (`SN_REQ_DESC_8_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_8 <= sn_req_desc_8_acaddr_0_reg;
               (`SN_REQ_DESC_8_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_8 <= sn_req_desc_8_acaddr_1_reg;
               (`SN_REQ_DESC_8_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_8 <= sn_req_desc_8_acaddr_2_reg;
               (`SN_REQ_DESC_8_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_8 <= sn_req_desc_8_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_8 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_9 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_9_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_9 <= sn_req_desc_9_attr_reg;
               (`SN_REQ_DESC_9_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_9 <= sn_req_desc_9_acaddr_0_reg;
               (`SN_REQ_DESC_9_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_9 <= sn_req_desc_9_acaddr_1_reg;
               (`SN_REQ_DESC_9_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_9 <= sn_req_desc_9_acaddr_2_reg;
               (`SN_REQ_DESC_9_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_9 <= sn_req_desc_9_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_9 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_a <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_A_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_a <= sn_req_desc_a_attr_reg;
               (`SN_REQ_DESC_A_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_a <= sn_req_desc_a_acaddr_0_reg;
               (`SN_REQ_DESC_A_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_a <= sn_req_desc_a_acaddr_1_reg;
               (`SN_REQ_DESC_A_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_a <= sn_req_desc_a_acaddr_2_reg;
               (`SN_REQ_DESC_A_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_a <= sn_req_desc_a_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_a <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_b <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_B_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_b <= sn_req_desc_b_attr_reg;
               (`SN_REQ_DESC_B_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_b <= sn_req_desc_b_acaddr_0_reg;
               (`SN_REQ_DESC_B_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_b <= sn_req_desc_b_acaddr_1_reg;
               (`SN_REQ_DESC_B_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_b <= sn_req_desc_b_acaddr_2_reg;
               (`SN_REQ_DESC_B_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_b <= sn_req_desc_b_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_b <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_c <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_C_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_c <= sn_req_desc_c_attr_reg;
               (`SN_REQ_DESC_C_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_c <= sn_req_desc_c_acaddr_0_reg;
               (`SN_REQ_DESC_C_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_c <= sn_req_desc_c_acaddr_1_reg;
               (`SN_REQ_DESC_C_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_c <= sn_req_desc_c_acaddr_2_reg;
               (`SN_REQ_DESC_C_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_c <= sn_req_desc_c_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_c <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_d <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_D_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_d <= sn_req_desc_d_attr_reg;
               (`SN_REQ_DESC_D_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_d <= sn_req_desc_d_acaddr_0_reg;
               (`SN_REQ_DESC_D_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_d <= sn_req_desc_d_acaddr_1_reg;
               (`SN_REQ_DESC_D_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_d <= sn_req_desc_d_acaddr_2_reg;
               (`SN_REQ_DESC_D_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_d <= sn_req_desc_d_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_d <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_e <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_E_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_e <= sn_req_desc_e_attr_reg;
               (`SN_REQ_DESC_E_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_e <= sn_req_desc_e_acaddr_0_reg;
               (`SN_REQ_DESC_E_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_e <= sn_req_desc_e_acaddr_1_reg;
               (`SN_REQ_DESC_E_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_e <= sn_req_desc_e_acaddr_2_reg;
               (`SN_REQ_DESC_E_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_e <= sn_req_desc_e_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_e <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_req_desc_f <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_REQ_DESC_F_ATTR_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_f <= sn_req_desc_f_attr_reg;
               (`SN_REQ_DESC_F_ACADDR_0_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_f <= sn_req_desc_f_acaddr_0_reg;
               (`SN_REQ_DESC_F_ACADDR_1_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_f <= sn_req_desc_f_acaddr_1_reg;
               (`SN_REQ_DESC_F_ACADDR_2_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_f <= sn_req_desc_f_acaddr_2_reg;
               (`SN_REQ_DESC_F_ACADDR_3_REG_ADDR&'hFF) :reg_data_out_sn_req_desc_f <= sn_req_desc_f_acaddr_3_reg;
               default                                  :reg_data_out_sn_req_desc_f <= 32'b0      ;        
             endcase
	  end
     end




   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_0 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_0_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_0 <= sn_resp_desc_0_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_0 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_1 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_1_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_1 <= sn_resp_desc_1_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_1 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_2 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_2_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_2 <= sn_resp_desc_2_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_2 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_3 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_3_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_3 <= sn_resp_desc_3_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_3 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_4 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_4_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_4 <= sn_resp_desc_4_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_4 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_5 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_5_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_5 <= sn_resp_desc_5_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_5 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_6 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_6_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_6 <= sn_resp_desc_6_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_6 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_7 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_7_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_7 <= sn_resp_desc_7_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_7 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_8 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_8_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_8 <= sn_resp_desc_8_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_8 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_9 <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_9_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_9 <= sn_resp_desc_9_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_9 <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_a <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_A_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_a <= sn_resp_desc_a_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_a <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_b <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_B_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_b <= sn_resp_desc_b_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_b <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_c <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_C_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_c <= sn_resp_desc_c_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_c <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_d <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_D_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_d <= sn_resp_desc_d_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_d <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_e <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_E_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_e <= sn_resp_desc_e_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_e <= 32'b0      ;        
             endcase
	  end
     end


   always @( posedge clk )
     begin
	if (~resetn)
	  begin
             reg_data_out_sn_resp_desc_f <= 32'b0;
	  end
	else
	  begin
             case ({axi_araddr[7:0]})    


               (`SN_RESP_DESC_F_RESP_REG_ADDR&'hFF) :reg_data_out_sn_resp_desc_f <= sn_resp_desc_f_resp_reg;
               default                                  :reg_data_out_sn_resp_desc_f <= 32'b0      ;        
             endcase
	  end
     end






   

   localparam [15:0] VEC_L                                                       = 16'h0000; 

   localparam [15:0] VEC_0                                                       = 16'h0001; 
   localparam [15:0] VEC_1                                                       = 16'h0002; 
   localparam [15:0] VEC_2                                                       = 16'h0004; 
   localparam [15:0] VEC_3                                                       = 16'h0008; 
   localparam [15:0] VEC_4                                                       = 16'h0010; 
   localparam [15:0] VEC_5                                                       = 16'h0020; 
   localparam [15:0] VEC_6                                                       = 16'h0040; 
   localparam [15:0] VEC_7                                                       = 16'h0080; 
   localparam [15:0] VEC_8                                                       = 16'h0100; 
   localparam [15:0] VEC_9                                                       = 16'h0200; 
   localparam [15:0] VEC_A                                                       = 16'h0400; 
   localparam [15:0] VEC_B                                                       = 16'h0800; 
   localparam [15:0] VEC_C                                                       = 16'h1000; 
   localparam [15:0] VEC_D                                                       = 16'h2000; 
   localparam [15:0] VEC_E                                                       = 16'h4000; 
   localparam [15:0] VEC_F                                                       = 16'h8000; 


   always @(*)
     begin
        // Address decoding for reading registers
        case ({  
                 reg_block_hit_sn_resp_desc
                 ,reg_block_hit_sn_req_desc
                 ,reg_block_hit_wr_resp_desc
                 ,reg_block_hit_wr_req_desc
                 ,reg_block_hit_rd_resp_desc
                 ,reg_block_hit_rd_req_desc
                 ,reg_block_hit_1
                 ,reg_block_hit_0
                 })
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b01} : reg_data_out <= reg_data_out_0;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b10} : reg_data_out <= reg_data_out_1;
          
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_0,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_0;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_1,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_1;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_2,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_2;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_3,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_3;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_4,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_4;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_5,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_5;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_6,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_6;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_7,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_7;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_8,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_8;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_9,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_9;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_A,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_a;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_B,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_b;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_C,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_c;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_D,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_d;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_E,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_e;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,VEC_F,2'b00} : reg_data_out <= reg_data_out_rd_req_desc_f;
          
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_0,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_0;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_1,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_1;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_2,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_2;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_3,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_3;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_4,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_4;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_5,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_5;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_6,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_6;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_7,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_7;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_8,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_8;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_9,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_9;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_A,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_a;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_B,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_b;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_C,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_c;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_D,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_d;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_E,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_e;
          {VEC_L,VEC_L,VEC_L,VEC_L,VEC_F,VEC_L,2'b00} : reg_data_out <= reg_data_out_rd_resp_desc_f;

          {VEC_L,VEC_L,VEC_L,VEC_0,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_0;
          {VEC_L,VEC_L,VEC_L,VEC_1,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_1;
          {VEC_L,VEC_L,VEC_L,VEC_2,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_2;
          {VEC_L,VEC_L,VEC_L,VEC_3,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_3;
          {VEC_L,VEC_L,VEC_L,VEC_4,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_4;
          {VEC_L,VEC_L,VEC_L,VEC_5,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_5;
          {VEC_L,VEC_L,VEC_L,VEC_6,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_6;
          {VEC_L,VEC_L,VEC_L,VEC_7,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_7;
          {VEC_L,VEC_L,VEC_L,VEC_8,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_8;
          {VEC_L,VEC_L,VEC_L,VEC_9,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_9;
          {VEC_L,VEC_L,VEC_L,VEC_A,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_a;
          {VEC_L,VEC_L,VEC_L,VEC_B,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_b;
          {VEC_L,VEC_L,VEC_L,VEC_C,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_c;
          {VEC_L,VEC_L,VEC_L,VEC_D,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_d;
          {VEC_L,VEC_L,VEC_L,VEC_E,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_e;
          {VEC_L,VEC_L,VEC_L,VEC_F,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_req_desc_f;

          {VEC_L,VEC_L,VEC_0,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_0;
          {VEC_L,VEC_L,VEC_1,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_1;
          {VEC_L,VEC_L,VEC_2,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_2;
          {VEC_L,VEC_L,VEC_3,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_3;
          {VEC_L,VEC_L,VEC_4,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_4;
          {VEC_L,VEC_L,VEC_5,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_5;
          {VEC_L,VEC_L,VEC_6,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_6;
          {VEC_L,VEC_L,VEC_7,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_7;
          {VEC_L,VEC_L,VEC_8,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_8;
          {VEC_L,VEC_L,VEC_9,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_9;
          {VEC_L,VEC_L,VEC_A,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_a;
          {VEC_L,VEC_L,VEC_B,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_b;
          {VEC_L,VEC_L,VEC_C,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_c;
          {VEC_L,VEC_L,VEC_D,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_d;
          {VEC_L,VEC_L,VEC_E,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_e;
          {VEC_L,VEC_L,VEC_F,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_wr_resp_desc_f;

          {VEC_L,VEC_0,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_0;
          {VEC_L,VEC_1,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_1;
          {VEC_L,VEC_2,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_2;
          {VEC_L,VEC_3,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_3;
          {VEC_L,VEC_4,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_4;
          {VEC_L,VEC_5,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_5;
          {VEC_L,VEC_6,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_6;
          {VEC_L,VEC_7,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_7;
          {VEC_L,VEC_8,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_8;
          {VEC_L,VEC_9,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_9;
          {VEC_L,VEC_A,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_a;
          {VEC_L,VEC_B,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_b;
          {VEC_L,VEC_C,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_c;
          {VEC_L,VEC_D,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_d;
          {VEC_L,VEC_E,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_e;
          {VEC_L,VEC_F,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_req_desc_f;

          {VEC_0,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_0;
          {VEC_1,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_1;
          {VEC_2,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_2;
          {VEC_3,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_3;
          {VEC_4,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_4;
          {VEC_5,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_5;
          {VEC_6,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_6;
          {VEC_7,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_7;
          {VEC_8,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_8;
          {VEC_9,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_9;
          {VEC_A,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_a;
          {VEC_B,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_b;
          {VEC_C,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_c;
          {VEC_D,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_d;
          {VEC_E,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_e;
          {VEC_F,VEC_L,VEC_L,VEC_L,VEC_L,VEC_L,2'b00} : reg_data_out <= reg_data_out_sn_resp_desc_f;



          default : reg_data_out <= 32'b0;
        endcase 
     end // always @ (*)

   always @( posedge clk )
     begin
	if (~resetn)
          reg_data_out_pipeline <= 32'b0;
	else
          reg_data_out_pipeline <= reg_data_out;
     end


   // fifo_pop_desc registers

   always @( posedge clk )
     begin
	if (~resetn)
          begin
             rd_req_fifo_pop_desc_conn  <= 1'b0; 
             wr_req_fifo_pop_desc_conn  <= 1'b0; 
             sn_resp_fifo_pop_desc_conn <= 1'b0;
             sn_data_fifo_pop_desc_conn <= 1'b0;
          end
	else
          begin
             
             if ( (~s_axi_arready && s_axi_arvalid) && (~|s_axi_araddr[BRIDGE_MSB:10])) 
               begin

                  case (s_axi_araddr[9:0]) 
                    
                    //
                    
                    `RD_REQ_FIFO_POP_DESC_REG_ADDR : begin 
                       rd_req_fifo_pop_desc_conn  <= 1'b1; 
                       wr_req_fifo_pop_desc_conn  <= 1'b0; 
                       sn_resp_fifo_pop_desc_conn <= 1'b0;
                       sn_data_fifo_pop_desc_conn <= 1'b0;
                    end 
                    `WR_REQ_FIFO_POP_DESC_REG_ADDR : begin 
                       rd_req_fifo_pop_desc_conn  <= 1'b0; 
                       wr_req_fifo_pop_desc_conn  <= 1'b1; 
                       sn_resp_fifo_pop_desc_conn <= 1'b0;
                       sn_data_fifo_pop_desc_conn <= 1'b0;
                    end 
                    `SN_RESP_FIFO_POP_DESC_REG_ADDR : begin 
                       rd_req_fifo_pop_desc_conn  <= 1'b0; 
                       wr_req_fifo_pop_desc_conn  <= 1'b0; 
                       sn_resp_fifo_pop_desc_conn <= 1'b1;
                       sn_data_fifo_pop_desc_conn <= 1'b0;
                    end 
                    `SN_DATA_FIFO_POP_DESC_REG_ADDR : begin 
                       rd_req_fifo_pop_desc_conn  <= 1'b0; 
                       wr_req_fifo_pop_desc_conn  <= 1'b0; 
                       sn_resp_fifo_pop_desc_conn <= 1'b0;
                       sn_data_fifo_pop_desc_conn <= 1'b1;
                       
                    end 
                    default : begin 
                       rd_req_fifo_pop_desc_conn  <= 1'b0; 
                       wr_req_fifo_pop_desc_conn  <= 1'b0; 
                       sn_resp_fifo_pop_desc_conn <= 1'b0;
                       sn_data_fifo_pop_desc_conn <= 1'b0;

                    end

                  endcase
               end
             else
               begin
                  rd_req_fifo_pop_desc_conn  <= 1'b0; 
                  wr_req_fifo_pop_desc_conn  <= 1'b0; 
                  sn_resp_fifo_pop_desc_conn <= 1'b0;
                  sn_data_fifo_pop_desc_conn <= 1'b0;
               end
             //end
          end
     end



   // Updating Mecahnism of RO registers
   

   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_intr_status_0_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_intr_status_0_reg_we[i])
		c2h_intr_status_0_reg[i] <= ih2rb_c2h_intr_status_0_reg[i];
              else
		c2h_intr_status_0_reg[i] <= c2h_intr_status_0_reg[i];
           end
	end
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_intr_status_1_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_intr_status_1_reg_we[i])
		c2h_intr_status_1_reg[i] <= ih2rb_c2h_intr_status_1_reg[i];
              else
		c2h_intr_status_1_reg[i] <= c2h_intr_status_1_reg[i];
           end
	end
     end // always @ (posedge clk)




   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             intr_c2h_toggle_status_0_reg[i] <= 1'b0;
           else begin
              if (ih2rb_intr_c2h_toggle_status_0_reg_we[i])
		intr_c2h_toggle_status_0_reg[i] <= ih2rb_intr_c2h_toggle_status_0_reg[i];
              else
		intr_c2h_toggle_status_0_reg[i] <= intr_c2h_toggle_status_0_reg[i];
           end
	end
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             intr_c2h_toggle_status_1_reg[i] <= 1'b0;
           else begin
              if (ih2rb_intr_c2h_toggle_status_1_reg_we[i])
		intr_c2h_toggle_status_1_reg[i] <= ih2rb_intr_c2h_toggle_status_1_reg[i];
              else
		intr_c2h_toggle_status_1_reg[i] <= intr_c2h_toggle_status_1_reg[i];
           end
	end
     end // always @ (posedge clk)
   



   // GPIO Registers 0-7 In   
   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_0_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_0_reg_we[i])
		c2h_gpio_0_reg[i] <= ih2rb_c2h_gpio_0_reg[i];
              else
		c2h_gpio_0_reg[i] <= c2h_gpio_0_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)
   

   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_1_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_1_reg_we[i])
		c2h_gpio_1_reg[i] <= ih2rb_c2h_gpio_1_reg[i];
              else
		c2h_gpio_1_reg[i] <= c2h_gpio_1_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)



   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_2_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_2_reg_we[i])
		c2h_gpio_2_reg[i] <= ih2rb_c2h_gpio_2_reg[i];
              else
		c2h_gpio_2_reg[i] <= c2h_gpio_2_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_3_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_3_reg_we[i])
		c2h_gpio_3_reg[i] <= ih2rb_c2h_gpio_3_reg[i];
              else
		c2h_gpio_3_reg[i] <= c2h_gpio_3_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_4_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_4_reg_we[i])
		c2h_gpio_4_reg[i] <= ih2rb_c2h_gpio_4_reg[i];
              else
		c2h_gpio_4_reg[i] <= c2h_gpio_4_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_5_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_5_reg_we[i])
		c2h_gpio_5_reg[i] <= ih2rb_c2h_gpio_5_reg[i];
              else
		c2h_gpio_5_reg[i] <= c2h_gpio_5_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_6_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_6_reg_we[i])
		c2h_gpio_6_reg[i] <= ih2rb_c2h_gpio_6_reg[i];
              else
		c2h_gpio_6_reg[i] <= c2h_gpio_6_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)


   always @(posedge clk)
     begin
	for (i=0; i<32; i=i+1)begin
           if (~rst_n)
             c2h_gpio_7_reg[i] <= 1'b0;
           else begin
              if (ih2rb_c2h_gpio_7_reg_we[i])
		c2h_gpio_7_reg[i] <= ih2rb_c2h_gpio_7_reg[i];
              else
		c2h_gpio_7_reg[i] <= c2h_gpio_7_reg[i];
           end
	end // for (i=0; i<32; i=i+1)
     end // always @ (posedge clk)
   

   //GPIO From 8-15 are not implemented

   always @(posedge clk)
     begin
	c2h_gpio_8_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_9_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_10_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_11_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_12_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_13_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_14_reg <= 0;    
     end
   
   always @(posedge clk)
     begin
	c2h_gpio_15_reg <= 0;    
     end

   //Register updation from RB

   always @(*) begin
      bridge_identification_reg <= BRIDGE_IDENTIFICATION_REG;
      last_bridge_reg <= LAST_BRIDGE_REG;
      version_reg <= VERSION_REG;
      bridge_type_reg <= BRIDGE_TYPE_REG;
      bridge_config_reg <= BRIDGE_CONFIG_REG;
      bridge_rd_user_config_reg <= BRIDGE_RD_USER_CONFIG_REG;
      bridge_wr_user_config_reg <= BRIDGE_WR_USER_CONFIG_REG;
      rd_max_desc_reg <= RD_MAX_DESC_REG;
      wr_max_desc_reg <= WR_MAX_DESC_REG;
      sn_max_desc_reg <= SN_MAX_DESC_REG;
   end


   // All W1C registers will be cleared by the Reg Block.
   // Effect of All clear registers and Ownership flip register on status* and ownership register will be implemented in C block.
   // This is done so that UC block need to make multiple/local copies of these regs for its internal operations.     


   //clear intr_comp registers from Reg Block

   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_resp_intr_comp_clear_reg_clear[i] <= 1'h0;
           else 
             if (~rd_resp_intr_comp_clear_reg_clear[i])begin
		if (rd_resp_intr_comp_clear_reg[i])
                  rd_resp_intr_comp_clear_reg_clear[i] <= 1'h1;
		else
                  rd_resp_intr_comp_clear_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  rd_resp_intr_comp_clear_reg_clear[i] <= 1'h0;
                else
                  rd_resp_intr_comp_clear_reg_clear[i] <= rd_resp_intr_comp_clear_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_resp_intr_comp_clear_reg_clear[i] <= 1'h0;
           else 
             if (~wr_resp_intr_comp_clear_reg_clear[i])begin
		if (wr_resp_intr_comp_clear_reg[i])
                  wr_resp_intr_comp_clear_reg_clear[i] <= 1'h1;
		else
                  wr_resp_intr_comp_clear_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  wr_resp_intr_comp_clear_reg_clear[i] <= 1'h0;
                else
                  wr_resp_intr_comp_clear_reg_clear[i] <= wr_resp_intr_comp_clear_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_req_intr_comp_clear_reg_clear[i] <= 1'h0;
           else 
             if (~sn_req_intr_comp_clear_reg_clear[i])begin
		if (sn_req_intr_comp_clear_reg[i])
                  sn_req_intr_comp_clear_reg_clear[i] <= 1'h1;
		else
                  sn_req_intr_comp_clear_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  sn_req_intr_comp_clear_reg_clear[i] <= 1'h0;
                else
                  sn_req_intr_comp_clear_reg_clear[i] <= sn_req_intr_comp_clear_reg_clear[i] ;
             end 
        end
     end

   //clear free_desc, fifo_push_desc registers from Reg Block

   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_free_desc_reg_clear[i] <= 1'h0;
           else 
             if (~rd_req_free_desc_reg_clear[i])begin
		if (rd_req_free_desc_reg[i])
                  rd_req_free_desc_reg_clear[i] <= 1'h1;
		else
                  rd_req_free_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  rd_req_free_desc_reg_clear[i] <= 1'h0;
                else
                  rd_req_free_desc_reg_clear[i] <= rd_req_free_desc_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_resp_fifo_push_desc_reg_clear[i] <= 1'h0;
           else 
             if (~rd_resp_fifo_push_desc_reg_clear[i])begin
		if (rd_resp_fifo_push_desc_reg[i])
                  rd_resp_fifo_push_desc_reg_clear[i] <= 1'h1;
		else
                  rd_resp_fifo_push_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  rd_resp_fifo_push_desc_reg_clear[i] <= 1'h0;
                else
                  rd_resp_fifo_push_desc_reg_clear[i] <= rd_resp_fifo_push_desc_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_free_desc_reg_clear[i] <= 1'h0;
           else 
             if (~wr_req_free_desc_reg_clear[i])begin
		if (wr_req_free_desc_reg[i])
                  wr_req_free_desc_reg_clear[i] <= 1'h1;
		else
                  wr_req_free_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  wr_req_free_desc_reg_clear[i] <= 1'h0;
                else
                  wr_req_free_desc_reg_clear[i] <= wr_req_free_desc_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_resp_fifo_push_desc_reg_clear[i] <= 1'h0;
           else 
             if (~wr_resp_fifo_push_desc_reg_clear[i])begin
		if (wr_resp_fifo_push_desc_reg[i])
                  wr_resp_fifo_push_desc_reg_clear[i] <= 1'h1;
		else
                  wr_resp_fifo_push_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  wr_resp_fifo_push_desc_reg_clear[i] <= 1'h0;
                else
                  wr_resp_fifo_push_desc_reg_clear[i] <= wr_resp_fifo_push_desc_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_req_fifo_push_desc_reg_clear[i] <= 1'h0;
           else 
             if (~sn_req_fifo_push_desc_reg_clear[i])begin
		if (sn_req_fifo_push_desc_reg[i])
                  sn_req_fifo_push_desc_reg_clear[i] <= 1'h1;
		else
                  sn_req_fifo_push_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  sn_req_fifo_push_desc_reg_clear[i] <= 1'h0;
                else
                  sn_req_fifo_push_desc_reg_clear[i] <= sn_req_fifo_push_desc_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_free_desc_reg_clear[i] <= 1'h0;
           else 
             if (~sn_resp_free_desc_reg_clear[i])begin
		if (sn_resp_free_desc_reg[i])
                  sn_resp_free_desc_reg_clear[i] <= 1'h1;
		else
                  sn_resp_free_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  sn_resp_free_desc_reg_clear[i] <= 1'h0;
                else
                  sn_resp_free_desc_reg_clear[i] <= sn_resp_free_desc_reg_clear[i] ;
             end 
        end
     end
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_data_free_desc_reg_clear[i] <= 1'h0;
           else 
             if (~sn_data_free_desc_reg_clear[i])begin
		if (sn_data_free_desc_reg[i])
                  sn_data_free_desc_reg_clear[i] <= 1'h1;
		else
                  sn_data_free_desc_reg_clear[i] <= 1'h0;
             end
             else begin
                if (~reg_wr_en)
                  sn_data_free_desc_reg_clear[i] <= 1'h0;
                else
                  sn_data_free_desc_reg_clear[i] <= sn_data_free_desc_reg_clear[i] ;
             end 
        end
     end

   
   always @( posedge clk )
     begin
        if (~rst_n)
          intr_error_status_reg[0] <= 1'b0;
        else begin
           if (uc2rb_intr_error_status_reg_we[0])
             intr_error_status_reg[0] <= uc2rb_intr_error_status_reg[0];
           else
             intr_error_status_reg[0] <= intr_error_status_reg[0];
        end
     end // always @ ( posedge clk )
   
   always @( posedge clk )
     begin
        if (~rst_n)
          intr_error_status_reg[1] <= 1'b0;
        else begin
           if (hm2rb_intr_error_status_reg_we[1])
             intr_error_status_reg[1] <= hm2rb_intr_error_status_reg[0];
           else
             intr_error_status_reg[1] <= intr_error_status_reg[1];
        end
     end // always @ ( posedge clk )
   
   

   // Tying of unused bits to 0

   always @(posedge clk)
     begin
        intr_error_status_reg[31:2] <= 30'h0;
     end
   


   always @( posedge clk )
     begin
        if (~rst_n)
          intr_error_clear_reg_clear[0] <= 1'b0;
        else begin 
           if (~intr_error_clear_reg_clear[0])begin
              if (intr_error_status_reg[0] && intr_error_clear_reg[0]) 
		intr_error_clear_reg_clear[0] <= 1'b1;
              else
		intr_error_clear_reg_clear[0] <= 1'b0;
           end
           else begin
              if (~reg_wr_en)
		intr_error_clear_reg_clear[0] <= 1'b0;
              else
		intr_error_clear_reg_clear[0] <= intr_error_clear_reg_clear[0];
           end // else: !if(~intr_error_clear_reg_clear[0])
        end // else: !if(~rst_n)
     end // always @ ( posedge clk )
   
   always @( posedge clk )
     begin
        if (~rst_n)
          intr_error_clear_reg_clear[1] <= 1'b0;
        else begin 
           if (~intr_error_clear_reg_clear[1])begin
              if (intr_error_status_reg[1] && intr_error_clear_reg[1]) 
		intr_error_clear_reg_clear[1] <= 1'b1;
              else
		intr_error_clear_reg_clear[1] <= 1'b0;
           end
           else begin
              if (~reg_wr_en)
		intr_error_clear_reg_clear[1] <= 1'b0;
              else
		intr_error_clear_reg_clear[1] <= intr_error_clear_reg_clear[1];
           end // else: !if(~intr_error_clear_reg_clear[0])
        end // else: !if(~rst_n)
     end // always @ ( posedge clk )

   always @( posedge clk )
     begin
        if (~rst_n)
          intr_error_clear_reg_clear[2] <= 1'b0;
        else begin 
           if (~intr_error_clear_reg_clear[2])begin
              if (intr_error_status_reg[2] && intr_error_clear_reg[2]) 
		intr_error_clear_reg_clear[2] <= 1'b1;
              else
		intr_error_clear_reg_clear[2] <= 1'b0;
           end
           else begin
              if (~reg_wr_en)
		intr_error_clear_reg_clear[2] <= 1'b0;
              else
		intr_error_clear_reg_clear[2] <= intr_error_clear_reg_clear[2];
           end // else: !if(~intr_error_clear_reg_clear[0])
        end // else: !if(~rst_n)
     end // always @ ( posedge clk )
   
   always @( posedge clk )
     begin
        for (i = 3; i < 32 ; i = i + 1) begin
           intr_error_clear_reg_clear[i] <= 1'b0;
        end
     end // always @ ( posedge clk )




   // INTR_C2H_TOGGLE_CLEAR_0_REG
   always @( posedge clk )
     begin
	for(i = 0; i < 32; i = i + 1 )
	  begin
	     if (~rst_n)
	       intr_c2h_toggle_clear_0_reg_clear[i] <= 1'b0;
	     else begin 
		if (~intr_c2h_toggle_clear_0_reg_clear[i])begin
		   if (intr_c2h_toggle_clear_0_reg[i]) 
		     intr_c2h_toggle_clear_0_reg_clear[i] <= 1'b1;
		   else
		     intr_c2h_toggle_clear_0_reg_clear[i] <= 1'b0;
		end
		else begin
		   if (~reg_wr_en)
		     intr_c2h_toggle_clear_0_reg_clear[i] <= 1'b0;
		   else
		     intr_c2h_toggle_clear_0_reg_clear[i] <= intr_c2h_toggle_clear_0_reg_clear[i];
		end // else: !if(~intr_c2h_toggle_clear_0_reg_clear[i])
	     end // else: !if(~rst_n)
	  end // always @ ( posedge clk )
     end // always @ ( posedge clk )
   


   // INTR_C2H_TOGGLE_CLEAR_1_REG
   always @( posedge clk )
     begin
	for(i = 0; i < 32; i = i + 1 )
	  begin
	     if (~rst_n)
	       intr_c2h_toggle_clear_1_reg_clear[i] <= 1'b0;
	     else begin 
		if (~intr_c2h_toggle_clear_1_reg_clear[i])begin
		   if (intr_c2h_toggle_clear_1_reg[i]) 
		     intr_c2h_toggle_clear_1_reg_clear[i] <= 1'b1;
		   else
		     intr_c2h_toggle_clear_1_reg_clear[i] <= 1'b0;
		end
		else begin
		   if (~reg_wr_en)
		     intr_c2h_toggle_clear_1_reg_clear[i] <= 1'b0;
		   else
		     intr_c2h_toggle_clear_1_reg_clear[i] <= intr_c2h_toggle_clear_1_reg_clear[i];
		end // else: !if(~intr_c2h_toggle_clear_0_reg_clear[i])
	     end // else: !if(~rst_n)
	  end // always @ ( posedge clk )
     end // always @ ( posedge clk )



   


   //INTR_STATUS_REG
   always @( posedge clk )
     begin
        if (~rst_n)
          intr_status_reg <= 32'b0;
        else
          intr_status_reg <= { 21'b0, |(sn_data_fifo_fill_level_reg), |(sn_resp_fifo_fill_level_reg), |(sn_req_intr_comp_status_reg), |(wr_resp_intr_comp_status_reg), |(wr_req_fifo_fill_level_reg), |(rd_resp_intr_comp_status_reg), |(rd_req_fifo_fill_level_reg), 1'b0, |({ intr_c2h_toggle_status_0_reg , intr_c2h_toggle_status_1_reg }), |(intr_error_status_reg), 1'b0 };
     end

   //Register updation from UC

   //RD_REQ_FIFO_POP_DESC_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_fifo_pop_desc_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_fifo_pop_desc_reg_we[i])
               rd_req_fifo_pop_desc_reg[i] <= uc2rb_rd_req_fifo_pop_desc_reg[i];
             else 
               rd_req_fifo_pop_desc_reg[i] <= rd_req_fifo_pop_desc_reg[i];
        end
     end
   //RD_REQ_FIFO_FILL_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_fifo_fill_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_fifo_fill_level_reg_we[i])
               rd_req_fifo_fill_level_reg[i] <= uc2rb_rd_req_fifo_fill_level_reg[i];
             else 
               rd_req_fifo_fill_level_reg[i] <= rd_req_fifo_fill_level_reg[i];
        end
     end
   //RD_RESP_FIFO_FREE_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_resp_fifo_free_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_resp_fifo_free_level_reg_we[i])
               rd_resp_fifo_free_level_reg[i] <= uc2rb_rd_resp_fifo_free_level_reg[i];
             else 
               rd_resp_fifo_free_level_reg[i] <= rd_resp_fifo_free_level_reg[i];
        end
     end
   //RD_RESP_INTR_COMP_STATUS_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_resp_intr_comp_status_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_resp_intr_comp_status_reg_we[i])
               rd_resp_intr_comp_status_reg[i] <= uc2rb_rd_resp_intr_comp_status_reg[i];
             else 
               rd_resp_intr_comp_status_reg[i] <= rd_resp_intr_comp_status_reg[i];
        end
     end
   //WR_REQ_FIFO_POP_DESC_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_fifo_pop_desc_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_fifo_pop_desc_reg_we[i])
               wr_req_fifo_pop_desc_reg[i] <= uc2rb_wr_req_fifo_pop_desc_reg[i];
             else 
               wr_req_fifo_pop_desc_reg[i] <= wr_req_fifo_pop_desc_reg[i];
        end
     end
   //WR_REQ_FIFO_FILL_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_fifo_fill_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_fifo_fill_level_reg_we[i])
               wr_req_fifo_fill_level_reg[i] <= uc2rb_wr_req_fifo_fill_level_reg[i];
             else 
               wr_req_fifo_fill_level_reg[i] <= wr_req_fifo_fill_level_reg[i];
        end
     end
   //WR_RESP_FIFO_FREE_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_resp_fifo_free_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_resp_fifo_free_level_reg_we[i])
               wr_resp_fifo_free_level_reg[i] <= uc2rb_wr_resp_fifo_free_level_reg[i];
             else 
               wr_resp_fifo_free_level_reg[i] <= wr_resp_fifo_free_level_reg[i];
        end
     end
   //WR_RESP_INTR_COMP_STATUS_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_resp_intr_comp_status_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_resp_intr_comp_status_reg_we[i])
               wr_resp_intr_comp_status_reg[i] <= uc2rb_wr_resp_intr_comp_status_reg[i];
             else 
               wr_resp_intr_comp_status_reg[i] <= wr_resp_intr_comp_status_reg[i];
        end
     end
   //SN_REQ_FIFO_FREE_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_req_fifo_free_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_req_fifo_free_level_reg_we[i])
               sn_req_fifo_free_level_reg[i] <= uc2rb_sn_req_fifo_free_level_reg[i];
             else 
               sn_req_fifo_free_level_reg[i] <= sn_req_fifo_free_level_reg[i];
        end
     end
   //SN_REQ_INTR_COMP_STATUS_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_req_intr_comp_status_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_req_intr_comp_status_reg_we[i])
               sn_req_intr_comp_status_reg[i] <= uc2rb_sn_req_intr_comp_status_reg[i];
             else 
               sn_req_intr_comp_status_reg[i] <= sn_req_intr_comp_status_reg[i];
        end
     end
   //SN_RESP_FIFO_POP_DESC_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_fifo_pop_desc_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_fifo_pop_desc_reg_we[i])
               sn_resp_fifo_pop_desc_reg[i] <= uc2rb_sn_resp_fifo_pop_desc_reg[i];
             else 
               sn_resp_fifo_pop_desc_reg[i] <= sn_resp_fifo_pop_desc_reg[i];
        end
     end
   //SN_RESP_FIFO_FILL_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_fifo_fill_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_fifo_fill_level_reg_we[i])
               sn_resp_fifo_fill_level_reg[i] <= uc2rb_sn_resp_fifo_fill_level_reg[i];
             else 
               sn_resp_fifo_fill_level_reg[i] <= sn_resp_fifo_fill_level_reg[i];
        end
     end
   //SN_DATA_FIFO_POP_DESC_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_data_fifo_pop_desc_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_data_fifo_pop_desc_reg_we[i])
               sn_data_fifo_pop_desc_reg[i] <= uc2rb_sn_data_fifo_pop_desc_reg[i];
             else 
               sn_data_fifo_pop_desc_reg[i] <= sn_data_fifo_pop_desc_reg[i];
        end
     end
   //SN_DATA_FIFO_FILL_LEVEL_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_data_fifo_fill_level_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_data_fifo_fill_level_reg_we[i])
               sn_data_fifo_fill_level_reg[i] <= uc2rb_sn_data_fifo_fill_level_reg[i];
             else 
               sn_data_fifo_fill_level_reg[i] <= sn_data_fifo_fill_level_reg[i];
        end
     end
   //RD_REQ_DESC_0_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_txn_type_reg_we[i])
               rd_req_desc_0_txn_type_reg[i] <= uc2rb_rd_req_desc_0_txn_type_reg[i];
             else 
               rd_req_desc_0_txn_type_reg[i] <= rd_req_desc_0_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_0_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_size_reg_we[i])
               rd_req_desc_0_size_reg[i] <= uc2rb_rd_req_desc_0_size_reg[i];
             else 
               rd_req_desc_0_size_reg[i] <= rd_req_desc_0_size_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axsize_reg_we[i])
               rd_req_desc_0_axsize_reg[i] <= uc2rb_rd_req_desc_0_axsize_reg[i];
             else 
               rd_req_desc_0_axsize_reg[i] <= rd_req_desc_0_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_0_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_attr_reg_we[i])
               rd_req_desc_0_attr_reg[i] <= uc2rb_rd_req_desc_0_attr_reg[i];
             else 
               rd_req_desc_0_attr_reg[i] <= rd_req_desc_0_attr_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axaddr_0_reg_we[i])
               rd_req_desc_0_axaddr_0_reg[i] <= uc2rb_rd_req_desc_0_axaddr_0_reg[i];
             else 
               rd_req_desc_0_axaddr_0_reg[i] <= rd_req_desc_0_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axaddr_1_reg_we[i])
               rd_req_desc_0_axaddr_1_reg[i] <= uc2rb_rd_req_desc_0_axaddr_1_reg[i];
             else 
               rd_req_desc_0_axaddr_1_reg[i] <= rd_req_desc_0_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axaddr_2_reg_we[i])
               rd_req_desc_0_axaddr_2_reg[i] <= uc2rb_rd_req_desc_0_axaddr_2_reg[i];
             else 
               rd_req_desc_0_axaddr_2_reg[i] <= rd_req_desc_0_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axaddr_3_reg_we[i])
               rd_req_desc_0_axaddr_3_reg[i] <= uc2rb_rd_req_desc_0_axaddr_3_reg[i];
             else 
               rd_req_desc_0_axaddr_3_reg[i] <= rd_req_desc_0_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axid_0_reg_we[i])
               rd_req_desc_0_axid_0_reg[i] <= uc2rb_rd_req_desc_0_axid_0_reg[i];
             else 
               rd_req_desc_0_axid_0_reg[i] <= rd_req_desc_0_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axid_1_reg_we[i])
               rd_req_desc_0_axid_1_reg[i] <= uc2rb_rd_req_desc_0_axid_1_reg[i];
             else 
               rd_req_desc_0_axid_1_reg[i] <= rd_req_desc_0_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axid_2_reg_we[i])
               rd_req_desc_0_axid_2_reg[i] <= uc2rb_rd_req_desc_0_axid_2_reg[i];
             else 
               rd_req_desc_0_axid_2_reg[i] <= rd_req_desc_0_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axid_3_reg_we[i])
               rd_req_desc_0_axid_3_reg[i] <= uc2rb_rd_req_desc_0_axid_3_reg[i];
             else 
               rd_req_desc_0_axid_3_reg[i] <= rd_req_desc_0_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_0_reg_we[i])
               rd_req_desc_0_axuser_0_reg[i] <= uc2rb_rd_req_desc_0_axuser_0_reg[i];
             else 
               rd_req_desc_0_axuser_0_reg[i] <= rd_req_desc_0_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_1_reg_we[i])
               rd_req_desc_0_axuser_1_reg[i] <= uc2rb_rd_req_desc_0_axuser_1_reg[i];
             else 
               rd_req_desc_0_axuser_1_reg[i] <= rd_req_desc_0_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_2_reg_we[i])
               rd_req_desc_0_axuser_2_reg[i] <= uc2rb_rd_req_desc_0_axuser_2_reg[i];
             else 
               rd_req_desc_0_axuser_2_reg[i] <= rd_req_desc_0_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_3_reg_we[i])
               rd_req_desc_0_axuser_3_reg[i] <= uc2rb_rd_req_desc_0_axuser_3_reg[i];
             else 
               rd_req_desc_0_axuser_3_reg[i] <= rd_req_desc_0_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_4_reg_we[i])
               rd_req_desc_0_axuser_4_reg[i] <= uc2rb_rd_req_desc_0_axuser_4_reg[i];
             else 
               rd_req_desc_0_axuser_4_reg[i] <= rd_req_desc_0_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_5_reg_we[i])
               rd_req_desc_0_axuser_5_reg[i] <= uc2rb_rd_req_desc_0_axuser_5_reg[i];
             else 
               rd_req_desc_0_axuser_5_reg[i] <= rd_req_desc_0_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_6_reg_we[i])
               rd_req_desc_0_axuser_6_reg[i] <= uc2rb_rd_req_desc_0_axuser_6_reg[i];
             else 
               rd_req_desc_0_axuser_6_reg[i] <= rd_req_desc_0_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_7_reg_we[i])
               rd_req_desc_0_axuser_7_reg[i] <= uc2rb_rd_req_desc_0_axuser_7_reg[i];
             else 
               rd_req_desc_0_axuser_7_reg[i] <= rd_req_desc_0_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_8_reg_we[i])
               rd_req_desc_0_axuser_8_reg[i] <= uc2rb_rd_req_desc_0_axuser_8_reg[i];
             else 
               rd_req_desc_0_axuser_8_reg[i] <= rd_req_desc_0_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_9_reg_we[i])
               rd_req_desc_0_axuser_9_reg[i] <= uc2rb_rd_req_desc_0_axuser_9_reg[i];
             else 
               rd_req_desc_0_axuser_9_reg[i] <= rd_req_desc_0_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_10_reg_we[i])
               rd_req_desc_0_axuser_10_reg[i] <= uc2rb_rd_req_desc_0_axuser_10_reg[i];
             else 
               rd_req_desc_0_axuser_10_reg[i] <= rd_req_desc_0_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_11_reg_we[i])
               rd_req_desc_0_axuser_11_reg[i] <= uc2rb_rd_req_desc_0_axuser_11_reg[i];
             else 
               rd_req_desc_0_axuser_11_reg[i] <= rd_req_desc_0_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_12_reg_we[i])
               rd_req_desc_0_axuser_12_reg[i] <= uc2rb_rd_req_desc_0_axuser_12_reg[i];
             else 
               rd_req_desc_0_axuser_12_reg[i] <= rd_req_desc_0_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_13_reg_we[i])
               rd_req_desc_0_axuser_13_reg[i] <= uc2rb_rd_req_desc_0_axuser_13_reg[i];
             else 
               rd_req_desc_0_axuser_13_reg[i] <= rd_req_desc_0_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_14_reg_we[i])
               rd_req_desc_0_axuser_14_reg[i] <= uc2rb_rd_req_desc_0_axuser_14_reg[i];
             else 
               rd_req_desc_0_axuser_14_reg[i] <= rd_req_desc_0_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_0_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_0_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_0_axuser_15_reg_we[i])
               rd_req_desc_0_axuser_15_reg[i] <= uc2rb_rd_req_desc_0_axuser_15_reg[i];
             else 
               rd_req_desc_0_axuser_15_reg[i] <= rd_req_desc_0_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_0_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_txn_type_reg_we[i])
               wr_req_desc_0_txn_type_reg[i] <= uc2rb_wr_req_desc_0_txn_type_reg[i];
             else 
               wr_req_desc_0_txn_type_reg[i] <= wr_req_desc_0_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_0_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_size_reg_we[i])
               wr_req_desc_0_size_reg[i] <= uc2rb_wr_req_desc_0_size_reg[i];
             else 
               wr_req_desc_0_size_reg[i] <= wr_req_desc_0_size_reg[i];
        end
     end
   //WR_REQ_DESC_0_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_data_offset_reg_we[i])
               wr_req_desc_0_data_offset_reg[i] <= uc2rb_wr_req_desc_0_data_offset_reg[i];
             else 
               wr_req_desc_0_data_offset_reg[i] <= wr_req_desc_0_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axsize_reg_we[i])
               wr_req_desc_0_axsize_reg[i] <= uc2rb_wr_req_desc_0_axsize_reg[i];
             else 
               wr_req_desc_0_axsize_reg[i] <= wr_req_desc_0_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_0_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_attr_reg_we[i])
               wr_req_desc_0_attr_reg[i] <= uc2rb_wr_req_desc_0_attr_reg[i];
             else 
               wr_req_desc_0_attr_reg[i] <= wr_req_desc_0_attr_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axaddr_0_reg_we[i])
               wr_req_desc_0_axaddr_0_reg[i] <= uc2rb_wr_req_desc_0_axaddr_0_reg[i];
             else 
               wr_req_desc_0_axaddr_0_reg[i] <= wr_req_desc_0_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axaddr_1_reg_we[i])
               wr_req_desc_0_axaddr_1_reg[i] <= uc2rb_wr_req_desc_0_axaddr_1_reg[i];
             else 
               wr_req_desc_0_axaddr_1_reg[i] <= wr_req_desc_0_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axaddr_2_reg_we[i])
               wr_req_desc_0_axaddr_2_reg[i] <= uc2rb_wr_req_desc_0_axaddr_2_reg[i];
             else 
               wr_req_desc_0_axaddr_2_reg[i] <= wr_req_desc_0_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axaddr_3_reg_we[i])
               wr_req_desc_0_axaddr_3_reg[i] <= uc2rb_wr_req_desc_0_axaddr_3_reg[i];
             else 
               wr_req_desc_0_axaddr_3_reg[i] <= wr_req_desc_0_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axid_0_reg_we[i])
               wr_req_desc_0_axid_0_reg[i] <= uc2rb_wr_req_desc_0_axid_0_reg[i];
             else 
               wr_req_desc_0_axid_0_reg[i] <= wr_req_desc_0_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axid_1_reg_we[i])
               wr_req_desc_0_axid_1_reg[i] <= uc2rb_wr_req_desc_0_axid_1_reg[i];
             else 
               wr_req_desc_0_axid_1_reg[i] <= wr_req_desc_0_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axid_2_reg_we[i])
               wr_req_desc_0_axid_2_reg[i] <= uc2rb_wr_req_desc_0_axid_2_reg[i];
             else 
               wr_req_desc_0_axid_2_reg[i] <= wr_req_desc_0_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axid_3_reg_we[i])
               wr_req_desc_0_axid_3_reg[i] <= uc2rb_wr_req_desc_0_axid_3_reg[i];
             else 
               wr_req_desc_0_axid_3_reg[i] <= wr_req_desc_0_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_0_reg_we[i])
               wr_req_desc_0_axuser_0_reg[i] <= uc2rb_wr_req_desc_0_axuser_0_reg[i];
             else 
               wr_req_desc_0_axuser_0_reg[i] <= wr_req_desc_0_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_1_reg_we[i])
               wr_req_desc_0_axuser_1_reg[i] <= uc2rb_wr_req_desc_0_axuser_1_reg[i];
             else 
               wr_req_desc_0_axuser_1_reg[i] <= wr_req_desc_0_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_2_reg_we[i])
               wr_req_desc_0_axuser_2_reg[i] <= uc2rb_wr_req_desc_0_axuser_2_reg[i];
             else 
               wr_req_desc_0_axuser_2_reg[i] <= wr_req_desc_0_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_3_reg_we[i])
               wr_req_desc_0_axuser_3_reg[i] <= uc2rb_wr_req_desc_0_axuser_3_reg[i];
             else 
               wr_req_desc_0_axuser_3_reg[i] <= wr_req_desc_0_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_4_reg_we[i])
               wr_req_desc_0_axuser_4_reg[i] <= uc2rb_wr_req_desc_0_axuser_4_reg[i];
             else 
               wr_req_desc_0_axuser_4_reg[i] <= wr_req_desc_0_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_5_reg_we[i])
               wr_req_desc_0_axuser_5_reg[i] <= uc2rb_wr_req_desc_0_axuser_5_reg[i];
             else 
               wr_req_desc_0_axuser_5_reg[i] <= wr_req_desc_0_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_6_reg_we[i])
               wr_req_desc_0_axuser_6_reg[i] <= uc2rb_wr_req_desc_0_axuser_6_reg[i];
             else 
               wr_req_desc_0_axuser_6_reg[i] <= wr_req_desc_0_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_7_reg_we[i])
               wr_req_desc_0_axuser_7_reg[i] <= uc2rb_wr_req_desc_0_axuser_7_reg[i];
             else 
               wr_req_desc_0_axuser_7_reg[i] <= wr_req_desc_0_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_8_reg_we[i])
               wr_req_desc_0_axuser_8_reg[i] <= uc2rb_wr_req_desc_0_axuser_8_reg[i];
             else 
               wr_req_desc_0_axuser_8_reg[i] <= wr_req_desc_0_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_9_reg_we[i])
               wr_req_desc_0_axuser_9_reg[i] <= uc2rb_wr_req_desc_0_axuser_9_reg[i];
             else 
               wr_req_desc_0_axuser_9_reg[i] <= wr_req_desc_0_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_10_reg_we[i])
               wr_req_desc_0_axuser_10_reg[i] <= uc2rb_wr_req_desc_0_axuser_10_reg[i];
             else 
               wr_req_desc_0_axuser_10_reg[i] <= wr_req_desc_0_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_11_reg_we[i])
               wr_req_desc_0_axuser_11_reg[i] <= uc2rb_wr_req_desc_0_axuser_11_reg[i];
             else 
               wr_req_desc_0_axuser_11_reg[i] <= wr_req_desc_0_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_12_reg_we[i])
               wr_req_desc_0_axuser_12_reg[i] <= uc2rb_wr_req_desc_0_axuser_12_reg[i];
             else 
               wr_req_desc_0_axuser_12_reg[i] <= wr_req_desc_0_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_13_reg_we[i])
               wr_req_desc_0_axuser_13_reg[i] <= uc2rb_wr_req_desc_0_axuser_13_reg[i];
             else 
               wr_req_desc_0_axuser_13_reg[i] <= wr_req_desc_0_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_14_reg_we[i])
               wr_req_desc_0_axuser_14_reg[i] <= uc2rb_wr_req_desc_0_axuser_14_reg[i];
             else 
               wr_req_desc_0_axuser_14_reg[i] <= wr_req_desc_0_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_0_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_axuser_15_reg_we[i])
               wr_req_desc_0_axuser_15_reg[i] <= uc2rb_wr_req_desc_0_axuser_15_reg[i];
             else 
               wr_req_desc_0_axuser_15_reg[i] <= wr_req_desc_0_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_0_reg_we[i])
               wr_req_desc_0_wuser_0_reg[i] <= uc2rb_wr_req_desc_0_wuser_0_reg[i];
             else 
               wr_req_desc_0_wuser_0_reg[i] <= wr_req_desc_0_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_1_reg_we[i])
               wr_req_desc_0_wuser_1_reg[i] <= uc2rb_wr_req_desc_0_wuser_1_reg[i];
             else 
               wr_req_desc_0_wuser_1_reg[i] <= wr_req_desc_0_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_2_reg_we[i])
               wr_req_desc_0_wuser_2_reg[i] <= uc2rb_wr_req_desc_0_wuser_2_reg[i];
             else 
               wr_req_desc_0_wuser_2_reg[i] <= wr_req_desc_0_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_3_reg_we[i])
               wr_req_desc_0_wuser_3_reg[i] <= uc2rb_wr_req_desc_0_wuser_3_reg[i];
             else 
               wr_req_desc_0_wuser_3_reg[i] <= wr_req_desc_0_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_4_reg_we[i])
               wr_req_desc_0_wuser_4_reg[i] <= uc2rb_wr_req_desc_0_wuser_4_reg[i];
             else 
               wr_req_desc_0_wuser_4_reg[i] <= wr_req_desc_0_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_5_reg_we[i])
               wr_req_desc_0_wuser_5_reg[i] <= uc2rb_wr_req_desc_0_wuser_5_reg[i];
             else 
               wr_req_desc_0_wuser_5_reg[i] <= wr_req_desc_0_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_6_reg_we[i])
               wr_req_desc_0_wuser_6_reg[i] <= uc2rb_wr_req_desc_0_wuser_6_reg[i];
             else 
               wr_req_desc_0_wuser_6_reg[i] <= wr_req_desc_0_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_7_reg_we[i])
               wr_req_desc_0_wuser_7_reg[i] <= uc2rb_wr_req_desc_0_wuser_7_reg[i];
             else 
               wr_req_desc_0_wuser_7_reg[i] <= wr_req_desc_0_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_8_reg_we[i])
               wr_req_desc_0_wuser_8_reg[i] <= uc2rb_wr_req_desc_0_wuser_8_reg[i];
             else 
               wr_req_desc_0_wuser_8_reg[i] <= wr_req_desc_0_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_9_reg_we[i])
               wr_req_desc_0_wuser_9_reg[i] <= uc2rb_wr_req_desc_0_wuser_9_reg[i];
             else 
               wr_req_desc_0_wuser_9_reg[i] <= wr_req_desc_0_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_10_reg_we[i])
               wr_req_desc_0_wuser_10_reg[i] <= uc2rb_wr_req_desc_0_wuser_10_reg[i];
             else 
               wr_req_desc_0_wuser_10_reg[i] <= wr_req_desc_0_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_11_reg_we[i])
               wr_req_desc_0_wuser_11_reg[i] <= uc2rb_wr_req_desc_0_wuser_11_reg[i];
             else 
               wr_req_desc_0_wuser_11_reg[i] <= wr_req_desc_0_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_12_reg_we[i])
               wr_req_desc_0_wuser_12_reg[i] <= uc2rb_wr_req_desc_0_wuser_12_reg[i];
             else 
               wr_req_desc_0_wuser_12_reg[i] <= wr_req_desc_0_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_13_reg_we[i])
               wr_req_desc_0_wuser_13_reg[i] <= uc2rb_wr_req_desc_0_wuser_13_reg[i];
             else 
               wr_req_desc_0_wuser_13_reg[i] <= wr_req_desc_0_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_14_reg_we[i])
               wr_req_desc_0_wuser_14_reg[i] <= uc2rb_wr_req_desc_0_wuser_14_reg[i];
             else 
               wr_req_desc_0_wuser_14_reg[i] <= wr_req_desc_0_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_0_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_0_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_0_wuser_15_reg_we[i])
               wr_req_desc_0_wuser_15_reg[i] <= uc2rb_wr_req_desc_0_wuser_15_reg[i];
             else 
               wr_req_desc_0_wuser_15_reg[i] <= wr_req_desc_0_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_0_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_0_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_0_resp_reg_we[i])
               sn_resp_desc_0_resp_reg[i] <= uc2rb_sn_resp_desc_0_resp_reg[i];
             else 
               sn_resp_desc_0_resp_reg[i] <= sn_resp_desc_0_resp_reg[i];
        end
     end
   //RD_REQ_DESC_1_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_txn_type_reg_we[i])
               rd_req_desc_1_txn_type_reg[i] <= uc2rb_rd_req_desc_1_txn_type_reg[i];
             else 
               rd_req_desc_1_txn_type_reg[i] <= rd_req_desc_1_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_1_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_size_reg_we[i])
               rd_req_desc_1_size_reg[i] <= uc2rb_rd_req_desc_1_size_reg[i];
             else 
               rd_req_desc_1_size_reg[i] <= rd_req_desc_1_size_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axsize_reg_we[i])
               rd_req_desc_1_axsize_reg[i] <= uc2rb_rd_req_desc_1_axsize_reg[i];
             else 
               rd_req_desc_1_axsize_reg[i] <= rd_req_desc_1_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_1_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_attr_reg_we[i])
               rd_req_desc_1_attr_reg[i] <= uc2rb_rd_req_desc_1_attr_reg[i];
             else 
               rd_req_desc_1_attr_reg[i] <= rd_req_desc_1_attr_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axaddr_0_reg_we[i])
               rd_req_desc_1_axaddr_0_reg[i] <= uc2rb_rd_req_desc_1_axaddr_0_reg[i];
             else 
               rd_req_desc_1_axaddr_0_reg[i] <= rd_req_desc_1_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axaddr_1_reg_we[i])
               rd_req_desc_1_axaddr_1_reg[i] <= uc2rb_rd_req_desc_1_axaddr_1_reg[i];
             else 
               rd_req_desc_1_axaddr_1_reg[i] <= rd_req_desc_1_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axaddr_2_reg_we[i])
               rd_req_desc_1_axaddr_2_reg[i] <= uc2rb_rd_req_desc_1_axaddr_2_reg[i];
             else 
               rd_req_desc_1_axaddr_2_reg[i] <= rd_req_desc_1_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axaddr_3_reg_we[i])
               rd_req_desc_1_axaddr_3_reg[i] <= uc2rb_rd_req_desc_1_axaddr_3_reg[i];
             else 
               rd_req_desc_1_axaddr_3_reg[i] <= rd_req_desc_1_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axid_0_reg_we[i])
               rd_req_desc_1_axid_0_reg[i] <= uc2rb_rd_req_desc_1_axid_0_reg[i];
             else 
               rd_req_desc_1_axid_0_reg[i] <= rd_req_desc_1_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axid_1_reg_we[i])
               rd_req_desc_1_axid_1_reg[i] <= uc2rb_rd_req_desc_1_axid_1_reg[i];
             else 
               rd_req_desc_1_axid_1_reg[i] <= rd_req_desc_1_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axid_2_reg_we[i])
               rd_req_desc_1_axid_2_reg[i] <= uc2rb_rd_req_desc_1_axid_2_reg[i];
             else 
               rd_req_desc_1_axid_2_reg[i] <= rd_req_desc_1_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axid_3_reg_we[i])
               rd_req_desc_1_axid_3_reg[i] <= uc2rb_rd_req_desc_1_axid_3_reg[i];
             else 
               rd_req_desc_1_axid_3_reg[i] <= rd_req_desc_1_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_0_reg_we[i])
               rd_req_desc_1_axuser_0_reg[i] <= uc2rb_rd_req_desc_1_axuser_0_reg[i];
             else 
               rd_req_desc_1_axuser_0_reg[i] <= rd_req_desc_1_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_1_reg_we[i])
               rd_req_desc_1_axuser_1_reg[i] <= uc2rb_rd_req_desc_1_axuser_1_reg[i];
             else 
               rd_req_desc_1_axuser_1_reg[i] <= rd_req_desc_1_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_2_reg_we[i])
               rd_req_desc_1_axuser_2_reg[i] <= uc2rb_rd_req_desc_1_axuser_2_reg[i];
             else 
               rd_req_desc_1_axuser_2_reg[i] <= rd_req_desc_1_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_3_reg_we[i])
               rd_req_desc_1_axuser_3_reg[i] <= uc2rb_rd_req_desc_1_axuser_3_reg[i];
             else 
               rd_req_desc_1_axuser_3_reg[i] <= rd_req_desc_1_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_4_reg_we[i])
               rd_req_desc_1_axuser_4_reg[i] <= uc2rb_rd_req_desc_1_axuser_4_reg[i];
             else 
               rd_req_desc_1_axuser_4_reg[i] <= rd_req_desc_1_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_5_reg_we[i])
               rd_req_desc_1_axuser_5_reg[i] <= uc2rb_rd_req_desc_1_axuser_5_reg[i];
             else 
               rd_req_desc_1_axuser_5_reg[i] <= rd_req_desc_1_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_6_reg_we[i])
               rd_req_desc_1_axuser_6_reg[i] <= uc2rb_rd_req_desc_1_axuser_6_reg[i];
             else 
               rd_req_desc_1_axuser_6_reg[i] <= rd_req_desc_1_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_7_reg_we[i])
               rd_req_desc_1_axuser_7_reg[i] <= uc2rb_rd_req_desc_1_axuser_7_reg[i];
             else 
               rd_req_desc_1_axuser_7_reg[i] <= rd_req_desc_1_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_8_reg_we[i])
               rd_req_desc_1_axuser_8_reg[i] <= uc2rb_rd_req_desc_1_axuser_8_reg[i];
             else 
               rd_req_desc_1_axuser_8_reg[i] <= rd_req_desc_1_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_9_reg_we[i])
               rd_req_desc_1_axuser_9_reg[i] <= uc2rb_rd_req_desc_1_axuser_9_reg[i];
             else 
               rd_req_desc_1_axuser_9_reg[i] <= rd_req_desc_1_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_10_reg_we[i])
               rd_req_desc_1_axuser_10_reg[i] <= uc2rb_rd_req_desc_1_axuser_10_reg[i];
             else 
               rd_req_desc_1_axuser_10_reg[i] <= rd_req_desc_1_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_11_reg_we[i])
               rd_req_desc_1_axuser_11_reg[i] <= uc2rb_rd_req_desc_1_axuser_11_reg[i];
             else 
               rd_req_desc_1_axuser_11_reg[i] <= rd_req_desc_1_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_12_reg_we[i])
               rd_req_desc_1_axuser_12_reg[i] <= uc2rb_rd_req_desc_1_axuser_12_reg[i];
             else 
               rd_req_desc_1_axuser_12_reg[i] <= rd_req_desc_1_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_13_reg_we[i])
               rd_req_desc_1_axuser_13_reg[i] <= uc2rb_rd_req_desc_1_axuser_13_reg[i];
             else 
               rd_req_desc_1_axuser_13_reg[i] <= rd_req_desc_1_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_14_reg_we[i])
               rd_req_desc_1_axuser_14_reg[i] <= uc2rb_rd_req_desc_1_axuser_14_reg[i];
             else 
               rd_req_desc_1_axuser_14_reg[i] <= rd_req_desc_1_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_1_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_1_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_1_axuser_15_reg_we[i])
               rd_req_desc_1_axuser_15_reg[i] <= uc2rb_rd_req_desc_1_axuser_15_reg[i];
             else 
               rd_req_desc_1_axuser_15_reg[i] <= rd_req_desc_1_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_1_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_txn_type_reg_we[i])
               wr_req_desc_1_txn_type_reg[i] <= uc2rb_wr_req_desc_1_txn_type_reg[i];
             else 
               wr_req_desc_1_txn_type_reg[i] <= wr_req_desc_1_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_1_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_size_reg_we[i])
               wr_req_desc_1_size_reg[i] <= uc2rb_wr_req_desc_1_size_reg[i];
             else 
               wr_req_desc_1_size_reg[i] <= wr_req_desc_1_size_reg[i];
        end
     end
   //WR_REQ_DESC_1_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_data_offset_reg_we[i])
               wr_req_desc_1_data_offset_reg[i] <= uc2rb_wr_req_desc_1_data_offset_reg[i];
             else 
               wr_req_desc_1_data_offset_reg[i] <= wr_req_desc_1_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axsize_reg_we[i])
               wr_req_desc_1_axsize_reg[i] <= uc2rb_wr_req_desc_1_axsize_reg[i];
             else 
               wr_req_desc_1_axsize_reg[i] <= wr_req_desc_1_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_1_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_attr_reg_we[i])
               wr_req_desc_1_attr_reg[i] <= uc2rb_wr_req_desc_1_attr_reg[i];
             else 
               wr_req_desc_1_attr_reg[i] <= wr_req_desc_1_attr_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axaddr_0_reg_we[i])
               wr_req_desc_1_axaddr_0_reg[i] <= uc2rb_wr_req_desc_1_axaddr_0_reg[i];
             else 
               wr_req_desc_1_axaddr_0_reg[i] <= wr_req_desc_1_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axaddr_1_reg_we[i])
               wr_req_desc_1_axaddr_1_reg[i] <= uc2rb_wr_req_desc_1_axaddr_1_reg[i];
             else 
               wr_req_desc_1_axaddr_1_reg[i] <= wr_req_desc_1_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axaddr_2_reg_we[i])
               wr_req_desc_1_axaddr_2_reg[i] <= uc2rb_wr_req_desc_1_axaddr_2_reg[i];
             else 
               wr_req_desc_1_axaddr_2_reg[i] <= wr_req_desc_1_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axaddr_3_reg_we[i])
               wr_req_desc_1_axaddr_3_reg[i] <= uc2rb_wr_req_desc_1_axaddr_3_reg[i];
             else 
               wr_req_desc_1_axaddr_3_reg[i] <= wr_req_desc_1_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axid_0_reg_we[i])
               wr_req_desc_1_axid_0_reg[i] <= uc2rb_wr_req_desc_1_axid_0_reg[i];
             else 
               wr_req_desc_1_axid_0_reg[i] <= wr_req_desc_1_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axid_1_reg_we[i])
               wr_req_desc_1_axid_1_reg[i] <= uc2rb_wr_req_desc_1_axid_1_reg[i];
             else 
               wr_req_desc_1_axid_1_reg[i] <= wr_req_desc_1_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axid_2_reg_we[i])
               wr_req_desc_1_axid_2_reg[i] <= uc2rb_wr_req_desc_1_axid_2_reg[i];
             else 
               wr_req_desc_1_axid_2_reg[i] <= wr_req_desc_1_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axid_3_reg_we[i])
               wr_req_desc_1_axid_3_reg[i] <= uc2rb_wr_req_desc_1_axid_3_reg[i];
             else 
               wr_req_desc_1_axid_3_reg[i] <= wr_req_desc_1_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_0_reg_we[i])
               wr_req_desc_1_axuser_0_reg[i] <= uc2rb_wr_req_desc_1_axuser_0_reg[i];
             else 
               wr_req_desc_1_axuser_0_reg[i] <= wr_req_desc_1_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_1_reg_we[i])
               wr_req_desc_1_axuser_1_reg[i] <= uc2rb_wr_req_desc_1_axuser_1_reg[i];
             else 
               wr_req_desc_1_axuser_1_reg[i] <= wr_req_desc_1_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_2_reg_we[i])
               wr_req_desc_1_axuser_2_reg[i] <= uc2rb_wr_req_desc_1_axuser_2_reg[i];
             else 
               wr_req_desc_1_axuser_2_reg[i] <= wr_req_desc_1_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_3_reg_we[i])
               wr_req_desc_1_axuser_3_reg[i] <= uc2rb_wr_req_desc_1_axuser_3_reg[i];
             else 
               wr_req_desc_1_axuser_3_reg[i] <= wr_req_desc_1_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_4_reg_we[i])
               wr_req_desc_1_axuser_4_reg[i] <= uc2rb_wr_req_desc_1_axuser_4_reg[i];
             else 
               wr_req_desc_1_axuser_4_reg[i] <= wr_req_desc_1_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_5_reg_we[i])
               wr_req_desc_1_axuser_5_reg[i] <= uc2rb_wr_req_desc_1_axuser_5_reg[i];
             else 
               wr_req_desc_1_axuser_5_reg[i] <= wr_req_desc_1_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_6_reg_we[i])
               wr_req_desc_1_axuser_6_reg[i] <= uc2rb_wr_req_desc_1_axuser_6_reg[i];
             else 
               wr_req_desc_1_axuser_6_reg[i] <= wr_req_desc_1_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_7_reg_we[i])
               wr_req_desc_1_axuser_7_reg[i] <= uc2rb_wr_req_desc_1_axuser_7_reg[i];
             else 
               wr_req_desc_1_axuser_7_reg[i] <= wr_req_desc_1_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_8_reg_we[i])
               wr_req_desc_1_axuser_8_reg[i] <= uc2rb_wr_req_desc_1_axuser_8_reg[i];
             else 
               wr_req_desc_1_axuser_8_reg[i] <= wr_req_desc_1_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_9_reg_we[i])
               wr_req_desc_1_axuser_9_reg[i] <= uc2rb_wr_req_desc_1_axuser_9_reg[i];
             else 
               wr_req_desc_1_axuser_9_reg[i] <= wr_req_desc_1_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_10_reg_we[i])
               wr_req_desc_1_axuser_10_reg[i] <= uc2rb_wr_req_desc_1_axuser_10_reg[i];
             else 
               wr_req_desc_1_axuser_10_reg[i] <= wr_req_desc_1_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_11_reg_we[i])
               wr_req_desc_1_axuser_11_reg[i] <= uc2rb_wr_req_desc_1_axuser_11_reg[i];
             else 
               wr_req_desc_1_axuser_11_reg[i] <= wr_req_desc_1_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_12_reg_we[i])
               wr_req_desc_1_axuser_12_reg[i] <= uc2rb_wr_req_desc_1_axuser_12_reg[i];
             else 
               wr_req_desc_1_axuser_12_reg[i] <= wr_req_desc_1_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_13_reg_we[i])
               wr_req_desc_1_axuser_13_reg[i] <= uc2rb_wr_req_desc_1_axuser_13_reg[i];
             else 
               wr_req_desc_1_axuser_13_reg[i] <= wr_req_desc_1_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_14_reg_we[i])
               wr_req_desc_1_axuser_14_reg[i] <= uc2rb_wr_req_desc_1_axuser_14_reg[i];
             else 
               wr_req_desc_1_axuser_14_reg[i] <= wr_req_desc_1_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_1_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_axuser_15_reg_we[i])
               wr_req_desc_1_axuser_15_reg[i] <= uc2rb_wr_req_desc_1_axuser_15_reg[i];
             else 
               wr_req_desc_1_axuser_15_reg[i] <= wr_req_desc_1_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_0_reg_we[i])
               wr_req_desc_1_wuser_0_reg[i] <= uc2rb_wr_req_desc_1_wuser_0_reg[i];
             else 
               wr_req_desc_1_wuser_0_reg[i] <= wr_req_desc_1_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_1_reg_we[i])
               wr_req_desc_1_wuser_1_reg[i] <= uc2rb_wr_req_desc_1_wuser_1_reg[i];
             else 
               wr_req_desc_1_wuser_1_reg[i] <= wr_req_desc_1_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_2_reg_we[i])
               wr_req_desc_1_wuser_2_reg[i] <= uc2rb_wr_req_desc_1_wuser_2_reg[i];
             else 
               wr_req_desc_1_wuser_2_reg[i] <= wr_req_desc_1_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_3_reg_we[i])
               wr_req_desc_1_wuser_3_reg[i] <= uc2rb_wr_req_desc_1_wuser_3_reg[i];
             else 
               wr_req_desc_1_wuser_3_reg[i] <= wr_req_desc_1_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_4_reg_we[i])
               wr_req_desc_1_wuser_4_reg[i] <= uc2rb_wr_req_desc_1_wuser_4_reg[i];
             else 
               wr_req_desc_1_wuser_4_reg[i] <= wr_req_desc_1_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_5_reg_we[i])
               wr_req_desc_1_wuser_5_reg[i] <= uc2rb_wr_req_desc_1_wuser_5_reg[i];
             else 
               wr_req_desc_1_wuser_5_reg[i] <= wr_req_desc_1_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_6_reg_we[i])
               wr_req_desc_1_wuser_6_reg[i] <= uc2rb_wr_req_desc_1_wuser_6_reg[i];
             else 
               wr_req_desc_1_wuser_6_reg[i] <= wr_req_desc_1_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_7_reg_we[i])
               wr_req_desc_1_wuser_7_reg[i] <= uc2rb_wr_req_desc_1_wuser_7_reg[i];
             else 
               wr_req_desc_1_wuser_7_reg[i] <= wr_req_desc_1_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_8_reg_we[i])
               wr_req_desc_1_wuser_8_reg[i] <= uc2rb_wr_req_desc_1_wuser_8_reg[i];
             else 
               wr_req_desc_1_wuser_8_reg[i] <= wr_req_desc_1_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_9_reg_we[i])
               wr_req_desc_1_wuser_9_reg[i] <= uc2rb_wr_req_desc_1_wuser_9_reg[i];
             else 
               wr_req_desc_1_wuser_9_reg[i] <= wr_req_desc_1_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_10_reg_we[i])
               wr_req_desc_1_wuser_10_reg[i] <= uc2rb_wr_req_desc_1_wuser_10_reg[i];
             else 
               wr_req_desc_1_wuser_10_reg[i] <= wr_req_desc_1_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_11_reg_we[i])
               wr_req_desc_1_wuser_11_reg[i] <= uc2rb_wr_req_desc_1_wuser_11_reg[i];
             else 
               wr_req_desc_1_wuser_11_reg[i] <= wr_req_desc_1_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_12_reg_we[i])
               wr_req_desc_1_wuser_12_reg[i] <= uc2rb_wr_req_desc_1_wuser_12_reg[i];
             else 
               wr_req_desc_1_wuser_12_reg[i] <= wr_req_desc_1_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_13_reg_we[i])
               wr_req_desc_1_wuser_13_reg[i] <= uc2rb_wr_req_desc_1_wuser_13_reg[i];
             else 
               wr_req_desc_1_wuser_13_reg[i] <= wr_req_desc_1_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_14_reg_we[i])
               wr_req_desc_1_wuser_14_reg[i] <= uc2rb_wr_req_desc_1_wuser_14_reg[i];
             else 
               wr_req_desc_1_wuser_14_reg[i] <= wr_req_desc_1_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_1_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_1_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_1_wuser_15_reg_we[i])
               wr_req_desc_1_wuser_15_reg[i] <= uc2rb_wr_req_desc_1_wuser_15_reg[i];
             else 
               wr_req_desc_1_wuser_15_reg[i] <= wr_req_desc_1_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_1_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_1_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_1_resp_reg_we[i])
               sn_resp_desc_1_resp_reg[i] <= uc2rb_sn_resp_desc_1_resp_reg[i];
             else 
               sn_resp_desc_1_resp_reg[i] <= sn_resp_desc_1_resp_reg[i];
        end
     end
   //RD_REQ_DESC_2_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_txn_type_reg_we[i])
               rd_req_desc_2_txn_type_reg[i] <= uc2rb_rd_req_desc_2_txn_type_reg[i];
             else 
               rd_req_desc_2_txn_type_reg[i] <= rd_req_desc_2_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_2_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_size_reg_we[i])
               rd_req_desc_2_size_reg[i] <= uc2rb_rd_req_desc_2_size_reg[i];
             else 
               rd_req_desc_2_size_reg[i] <= rd_req_desc_2_size_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axsize_reg_we[i])
               rd_req_desc_2_axsize_reg[i] <= uc2rb_rd_req_desc_2_axsize_reg[i];
             else 
               rd_req_desc_2_axsize_reg[i] <= rd_req_desc_2_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_2_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_attr_reg_we[i])
               rd_req_desc_2_attr_reg[i] <= uc2rb_rd_req_desc_2_attr_reg[i];
             else 
               rd_req_desc_2_attr_reg[i] <= rd_req_desc_2_attr_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axaddr_0_reg_we[i])
               rd_req_desc_2_axaddr_0_reg[i] <= uc2rb_rd_req_desc_2_axaddr_0_reg[i];
             else 
               rd_req_desc_2_axaddr_0_reg[i] <= rd_req_desc_2_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axaddr_1_reg_we[i])
               rd_req_desc_2_axaddr_1_reg[i] <= uc2rb_rd_req_desc_2_axaddr_1_reg[i];
             else 
               rd_req_desc_2_axaddr_1_reg[i] <= rd_req_desc_2_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axaddr_2_reg_we[i])
               rd_req_desc_2_axaddr_2_reg[i] <= uc2rb_rd_req_desc_2_axaddr_2_reg[i];
             else 
               rd_req_desc_2_axaddr_2_reg[i] <= rd_req_desc_2_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axaddr_3_reg_we[i])
               rd_req_desc_2_axaddr_3_reg[i] <= uc2rb_rd_req_desc_2_axaddr_3_reg[i];
             else 
               rd_req_desc_2_axaddr_3_reg[i] <= rd_req_desc_2_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axid_0_reg_we[i])
               rd_req_desc_2_axid_0_reg[i] <= uc2rb_rd_req_desc_2_axid_0_reg[i];
             else 
               rd_req_desc_2_axid_0_reg[i] <= rd_req_desc_2_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axid_1_reg_we[i])
               rd_req_desc_2_axid_1_reg[i] <= uc2rb_rd_req_desc_2_axid_1_reg[i];
             else 
               rd_req_desc_2_axid_1_reg[i] <= rd_req_desc_2_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axid_2_reg_we[i])
               rd_req_desc_2_axid_2_reg[i] <= uc2rb_rd_req_desc_2_axid_2_reg[i];
             else 
               rd_req_desc_2_axid_2_reg[i] <= rd_req_desc_2_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axid_3_reg_we[i])
               rd_req_desc_2_axid_3_reg[i] <= uc2rb_rd_req_desc_2_axid_3_reg[i];
             else 
               rd_req_desc_2_axid_3_reg[i] <= rd_req_desc_2_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_0_reg_we[i])
               rd_req_desc_2_axuser_0_reg[i] <= uc2rb_rd_req_desc_2_axuser_0_reg[i];
             else 
               rd_req_desc_2_axuser_0_reg[i] <= rd_req_desc_2_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_1_reg_we[i])
               rd_req_desc_2_axuser_1_reg[i] <= uc2rb_rd_req_desc_2_axuser_1_reg[i];
             else 
               rd_req_desc_2_axuser_1_reg[i] <= rd_req_desc_2_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_2_reg_we[i])
               rd_req_desc_2_axuser_2_reg[i] <= uc2rb_rd_req_desc_2_axuser_2_reg[i];
             else 
               rd_req_desc_2_axuser_2_reg[i] <= rd_req_desc_2_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_3_reg_we[i])
               rd_req_desc_2_axuser_3_reg[i] <= uc2rb_rd_req_desc_2_axuser_3_reg[i];
             else 
               rd_req_desc_2_axuser_3_reg[i] <= rd_req_desc_2_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_4_reg_we[i])
               rd_req_desc_2_axuser_4_reg[i] <= uc2rb_rd_req_desc_2_axuser_4_reg[i];
             else 
               rd_req_desc_2_axuser_4_reg[i] <= rd_req_desc_2_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_5_reg_we[i])
               rd_req_desc_2_axuser_5_reg[i] <= uc2rb_rd_req_desc_2_axuser_5_reg[i];
             else 
               rd_req_desc_2_axuser_5_reg[i] <= rd_req_desc_2_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_6_reg_we[i])
               rd_req_desc_2_axuser_6_reg[i] <= uc2rb_rd_req_desc_2_axuser_6_reg[i];
             else 
               rd_req_desc_2_axuser_6_reg[i] <= rd_req_desc_2_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_7_reg_we[i])
               rd_req_desc_2_axuser_7_reg[i] <= uc2rb_rd_req_desc_2_axuser_7_reg[i];
             else 
               rd_req_desc_2_axuser_7_reg[i] <= rd_req_desc_2_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_8_reg_we[i])
               rd_req_desc_2_axuser_8_reg[i] <= uc2rb_rd_req_desc_2_axuser_8_reg[i];
             else 
               rd_req_desc_2_axuser_8_reg[i] <= rd_req_desc_2_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_9_reg_we[i])
               rd_req_desc_2_axuser_9_reg[i] <= uc2rb_rd_req_desc_2_axuser_9_reg[i];
             else 
               rd_req_desc_2_axuser_9_reg[i] <= rd_req_desc_2_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_10_reg_we[i])
               rd_req_desc_2_axuser_10_reg[i] <= uc2rb_rd_req_desc_2_axuser_10_reg[i];
             else 
               rd_req_desc_2_axuser_10_reg[i] <= rd_req_desc_2_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_11_reg_we[i])
               rd_req_desc_2_axuser_11_reg[i] <= uc2rb_rd_req_desc_2_axuser_11_reg[i];
             else 
               rd_req_desc_2_axuser_11_reg[i] <= rd_req_desc_2_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_12_reg_we[i])
               rd_req_desc_2_axuser_12_reg[i] <= uc2rb_rd_req_desc_2_axuser_12_reg[i];
             else 
               rd_req_desc_2_axuser_12_reg[i] <= rd_req_desc_2_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_13_reg_we[i])
               rd_req_desc_2_axuser_13_reg[i] <= uc2rb_rd_req_desc_2_axuser_13_reg[i];
             else 
               rd_req_desc_2_axuser_13_reg[i] <= rd_req_desc_2_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_14_reg_we[i])
               rd_req_desc_2_axuser_14_reg[i] <= uc2rb_rd_req_desc_2_axuser_14_reg[i];
             else 
               rd_req_desc_2_axuser_14_reg[i] <= rd_req_desc_2_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_2_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_2_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_2_axuser_15_reg_we[i])
               rd_req_desc_2_axuser_15_reg[i] <= uc2rb_rd_req_desc_2_axuser_15_reg[i];
             else 
               rd_req_desc_2_axuser_15_reg[i] <= rd_req_desc_2_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_2_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_txn_type_reg_we[i])
               wr_req_desc_2_txn_type_reg[i] <= uc2rb_wr_req_desc_2_txn_type_reg[i];
             else 
               wr_req_desc_2_txn_type_reg[i] <= wr_req_desc_2_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_2_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_size_reg_we[i])
               wr_req_desc_2_size_reg[i] <= uc2rb_wr_req_desc_2_size_reg[i];
             else 
               wr_req_desc_2_size_reg[i] <= wr_req_desc_2_size_reg[i];
        end
     end
   //WR_REQ_DESC_2_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_data_offset_reg_we[i])
               wr_req_desc_2_data_offset_reg[i] <= uc2rb_wr_req_desc_2_data_offset_reg[i];
             else 
               wr_req_desc_2_data_offset_reg[i] <= wr_req_desc_2_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axsize_reg_we[i])
               wr_req_desc_2_axsize_reg[i] <= uc2rb_wr_req_desc_2_axsize_reg[i];
             else 
               wr_req_desc_2_axsize_reg[i] <= wr_req_desc_2_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_2_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_attr_reg_we[i])
               wr_req_desc_2_attr_reg[i] <= uc2rb_wr_req_desc_2_attr_reg[i];
             else 
               wr_req_desc_2_attr_reg[i] <= wr_req_desc_2_attr_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axaddr_0_reg_we[i])
               wr_req_desc_2_axaddr_0_reg[i] <= uc2rb_wr_req_desc_2_axaddr_0_reg[i];
             else 
               wr_req_desc_2_axaddr_0_reg[i] <= wr_req_desc_2_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axaddr_1_reg_we[i])
               wr_req_desc_2_axaddr_1_reg[i] <= uc2rb_wr_req_desc_2_axaddr_1_reg[i];
             else 
               wr_req_desc_2_axaddr_1_reg[i] <= wr_req_desc_2_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axaddr_2_reg_we[i])
               wr_req_desc_2_axaddr_2_reg[i] <= uc2rb_wr_req_desc_2_axaddr_2_reg[i];
             else 
               wr_req_desc_2_axaddr_2_reg[i] <= wr_req_desc_2_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axaddr_3_reg_we[i])
               wr_req_desc_2_axaddr_3_reg[i] <= uc2rb_wr_req_desc_2_axaddr_3_reg[i];
             else 
               wr_req_desc_2_axaddr_3_reg[i] <= wr_req_desc_2_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axid_0_reg_we[i])
               wr_req_desc_2_axid_0_reg[i] <= uc2rb_wr_req_desc_2_axid_0_reg[i];
             else 
               wr_req_desc_2_axid_0_reg[i] <= wr_req_desc_2_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axid_1_reg_we[i])
               wr_req_desc_2_axid_1_reg[i] <= uc2rb_wr_req_desc_2_axid_1_reg[i];
             else 
               wr_req_desc_2_axid_1_reg[i] <= wr_req_desc_2_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axid_2_reg_we[i])
               wr_req_desc_2_axid_2_reg[i] <= uc2rb_wr_req_desc_2_axid_2_reg[i];
             else 
               wr_req_desc_2_axid_2_reg[i] <= wr_req_desc_2_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axid_3_reg_we[i])
               wr_req_desc_2_axid_3_reg[i] <= uc2rb_wr_req_desc_2_axid_3_reg[i];
             else 
               wr_req_desc_2_axid_3_reg[i] <= wr_req_desc_2_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_0_reg_we[i])
               wr_req_desc_2_axuser_0_reg[i] <= uc2rb_wr_req_desc_2_axuser_0_reg[i];
             else 
               wr_req_desc_2_axuser_0_reg[i] <= wr_req_desc_2_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_1_reg_we[i])
               wr_req_desc_2_axuser_1_reg[i] <= uc2rb_wr_req_desc_2_axuser_1_reg[i];
             else 
               wr_req_desc_2_axuser_1_reg[i] <= wr_req_desc_2_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_2_reg_we[i])
               wr_req_desc_2_axuser_2_reg[i] <= uc2rb_wr_req_desc_2_axuser_2_reg[i];
             else 
               wr_req_desc_2_axuser_2_reg[i] <= wr_req_desc_2_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_3_reg_we[i])
               wr_req_desc_2_axuser_3_reg[i] <= uc2rb_wr_req_desc_2_axuser_3_reg[i];
             else 
               wr_req_desc_2_axuser_3_reg[i] <= wr_req_desc_2_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_4_reg_we[i])
               wr_req_desc_2_axuser_4_reg[i] <= uc2rb_wr_req_desc_2_axuser_4_reg[i];
             else 
               wr_req_desc_2_axuser_4_reg[i] <= wr_req_desc_2_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_5_reg_we[i])
               wr_req_desc_2_axuser_5_reg[i] <= uc2rb_wr_req_desc_2_axuser_5_reg[i];
             else 
               wr_req_desc_2_axuser_5_reg[i] <= wr_req_desc_2_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_6_reg_we[i])
               wr_req_desc_2_axuser_6_reg[i] <= uc2rb_wr_req_desc_2_axuser_6_reg[i];
             else 
               wr_req_desc_2_axuser_6_reg[i] <= wr_req_desc_2_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_7_reg_we[i])
               wr_req_desc_2_axuser_7_reg[i] <= uc2rb_wr_req_desc_2_axuser_7_reg[i];
             else 
               wr_req_desc_2_axuser_7_reg[i] <= wr_req_desc_2_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_8_reg_we[i])
               wr_req_desc_2_axuser_8_reg[i] <= uc2rb_wr_req_desc_2_axuser_8_reg[i];
             else 
               wr_req_desc_2_axuser_8_reg[i] <= wr_req_desc_2_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_9_reg_we[i])
               wr_req_desc_2_axuser_9_reg[i] <= uc2rb_wr_req_desc_2_axuser_9_reg[i];
             else 
               wr_req_desc_2_axuser_9_reg[i] <= wr_req_desc_2_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_10_reg_we[i])
               wr_req_desc_2_axuser_10_reg[i] <= uc2rb_wr_req_desc_2_axuser_10_reg[i];
             else 
               wr_req_desc_2_axuser_10_reg[i] <= wr_req_desc_2_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_11_reg_we[i])
               wr_req_desc_2_axuser_11_reg[i] <= uc2rb_wr_req_desc_2_axuser_11_reg[i];
             else 
               wr_req_desc_2_axuser_11_reg[i] <= wr_req_desc_2_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_12_reg_we[i])
               wr_req_desc_2_axuser_12_reg[i] <= uc2rb_wr_req_desc_2_axuser_12_reg[i];
             else 
               wr_req_desc_2_axuser_12_reg[i] <= wr_req_desc_2_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_13_reg_we[i])
               wr_req_desc_2_axuser_13_reg[i] <= uc2rb_wr_req_desc_2_axuser_13_reg[i];
             else 
               wr_req_desc_2_axuser_13_reg[i] <= wr_req_desc_2_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_14_reg_we[i])
               wr_req_desc_2_axuser_14_reg[i] <= uc2rb_wr_req_desc_2_axuser_14_reg[i];
             else 
               wr_req_desc_2_axuser_14_reg[i] <= wr_req_desc_2_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_2_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_axuser_15_reg_we[i])
               wr_req_desc_2_axuser_15_reg[i] <= uc2rb_wr_req_desc_2_axuser_15_reg[i];
             else 
               wr_req_desc_2_axuser_15_reg[i] <= wr_req_desc_2_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_0_reg_we[i])
               wr_req_desc_2_wuser_0_reg[i] <= uc2rb_wr_req_desc_2_wuser_0_reg[i];
             else 
               wr_req_desc_2_wuser_0_reg[i] <= wr_req_desc_2_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_1_reg_we[i])
               wr_req_desc_2_wuser_1_reg[i] <= uc2rb_wr_req_desc_2_wuser_1_reg[i];
             else 
               wr_req_desc_2_wuser_1_reg[i] <= wr_req_desc_2_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_2_reg_we[i])
               wr_req_desc_2_wuser_2_reg[i] <= uc2rb_wr_req_desc_2_wuser_2_reg[i];
             else 
               wr_req_desc_2_wuser_2_reg[i] <= wr_req_desc_2_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_3_reg_we[i])
               wr_req_desc_2_wuser_3_reg[i] <= uc2rb_wr_req_desc_2_wuser_3_reg[i];
             else 
               wr_req_desc_2_wuser_3_reg[i] <= wr_req_desc_2_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_4_reg_we[i])
               wr_req_desc_2_wuser_4_reg[i] <= uc2rb_wr_req_desc_2_wuser_4_reg[i];
             else 
               wr_req_desc_2_wuser_4_reg[i] <= wr_req_desc_2_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_5_reg_we[i])
               wr_req_desc_2_wuser_5_reg[i] <= uc2rb_wr_req_desc_2_wuser_5_reg[i];
             else 
               wr_req_desc_2_wuser_5_reg[i] <= wr_req_desc_2_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_6_reg_we[i])
               wr_req_desc_2_wuser_6_reg[i] <= uc2rb_wr_req_desc_2_wuser_6_reg[i];
             else 
               wr_req_desc_2_wuser_6_reg[i] <= wr_req_desc_2_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_7_reg_we[i])
               wr_req_desc_2_wuser_7_reg[i] <= uc2rb_wr_req_desc_2_wuser_7_reg[i];
             else 
               wr_req_desc_2_wuser_7_reg[i] <= wr_req_desc_2_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_8_reg_we[i])
               wr_req_desc_2_wuser_8_reg[i] <= uc2rb_wr_req_desc_2_wuser_8_reg[i];
             else 
               wr_req_desc_2_wuser_8_reg[i] <= wr_req_desc_2_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_9_reg_we[i])
               wr_req_desc_2_wuser_9_reg[i] <= uc2rb_wr_req_desc_2_wuser_9_reg[i];
             else 
               wr_req_desc_2_wuser_9_reg[i] <= wr_req_desc_2_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_10_reg_we[i])
               wr_req_desc_2_wuser_10_reg[i] <= uc2rb_wr_req_desc_2_wuser_10_reg[i];
             else 
               wr_req_desc_2_wuser_10_reg[i] <= wr_req_desc_2_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_11_reg_we[i])
               wr_req_desc_2_wuser_11_reg[i] <= uc2rb_wr_req_desc_2_wuser_11_reg[i];
             else 
               wr_req_desc_2_wuser_11_reg[i] <= wr_req_desc_2_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_12_reg_we[i])
               wr_req_desc_2_wuser_12_reg[i] <= uc2rb_wr_req_desc_2_wuser_12_reg[i];
             else 
               wr_req_desc_2_wuser_12_reg[i] <= wr_req_desc_2_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_13_reg_we[i])
               wr_req_desc_2_wuser_13_reg[i] <= uc2rb_wr_req_desc_2_wuser_13_reg[i];
             else 
               wr_req_desc_2_wuser_13_reg[i] <= wr_req_desc_2_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_14_reg_we[i])
               wr_req_desc_2_wuser_14_reg[i] <= uc2rb_wr_req_desc_2_wuser_14_reg[i];
             else 
               wr_req_desc_2_wuser_14_reg[i] <= wr_req_desc_2_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_2_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_2_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_2_wuser_15_reg_we[i])
               wr_req_desc_2_wuser_15_reg[i] <= uc2rb_wr_req_desc_2_wuser_15_reg[i];
             else 
               wr_req_desc_2_wuser_15_reg[i] <= wr_req_desc_2_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_2_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_2_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_2_resp_reg_we[i])
               sn_resp_desc_2_resp_reg[i] <= uc2rb_sn_resp_desc_2_resp_reg[i];
             else 
               sn_resp_desc_2_resp_reg[i] <= sn_resp_desc_2_resp_reg[i];
        end
     end
   //RD_REQ_DESC_3_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_txn_type_reg_we[i])
               rd_req_desc_3_txn_type_reg[i] <= uc2rb_rd_req_desc_3_txn_type_reg[i];
             else 
               rd_req_desc_3_txn_type_reg[i] <= rd_req_desc_3_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_3_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_size_reg_we[i])
               rd_req_desc_3_size_reg[i] <= uc2rb_rd_req_desc_3_size_reg[i];
             else 
               rd_req_desc_3_size_reg[i] <= rd_req_desc_3_size_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axsize_reg_we[i])
               rd_req_desc_3_axsize_reg[i] <= uc2rb_rd_req_desc_3_axsize_reg[i];
             else 
               rd_req_desc_3_axsize_reg[i] <= rd_req_desc_3_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_3_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_attr_reg_we[i])
               rd_req_desc_3_attr_reg[i] <= uc2rb_rd_req_desc_3_attr_reg[i];
             else 
               rd_req_desc_3_attr_reg[i] <= rd_req_desc_3_attr_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axaddr_0_reg_we[i])
               rd_req_desc_3_axaddr_0_reg[i] <= uc2rb_rd_req_desc_3_axaddr_0_reg[i];
             else 
               rd_req_desc_3_axaddr_0_reg[i] <= rd_req_desc_3_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axaddr_1_reg_we[i])
               rd_req_desc_3_axaddr_1_reg[i] <= uc2rb_rd_req_desc_3_axaddr_1_reg[i];
             else 
               rd_req_desc_3_axaddr_1_reg[i] <= rd_req_desc_3_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axaddr_2_reg_we[i])
               rd_req_desc_3_axaddr_2_reg[i] <= uc2rb_rd_req_desc_3_axaddr_2_reg[i];
             else 
               rd_req_desc_3_axaddr_2_reg[i] <= rd_req_desc_3_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axaddr_3_reg_we[i])
               rd_req_desc_3_axaddr_3_reg[i] <= uc2rb_rd_req_desc_3_axaddr_3_reg[i];
             else 
               rd_req_desc_3_axaddr_3_reg[i] <= rd_req_desc_3_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axid_0_reg_we[i])
               rd_req_desc_3_axid_0_reg[i] <= uc2rb_rd_req_desc_3_axid_0_reg[i];
             else 
               rd_req_desc_3_axid_0_reg[i] <= rd_req_desc_3_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axid_1_reg_we[i])
               rd_req_desc_3_axid_1_reg[i] <= uc2rb_rd_req_desc_3_axid_1_reg[i];
             else 
               rd_req_desc_3_axid_1_reg[i] <= rd_req_desc_3_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axid_2_reg_we[i])
               rd_req_desc_3_axid_2_reg[i] <= uc2rb_rd_req_desc_3_axid_2_reg[i];
             else 
               rd_req_desc_3_axid_2_reg[i] <= rd_req_desc_3_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axid_3_reg_we[i])
               rd_req_desc_3_axid_3_reg[i] <= uc2rb_rd_req_desc_3_axid_3_reg[i];
             else 
               rd_req_desc_3_axid_3_reg[i] <= rd_req_desc_3_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_0_reg_we[i])
               rd_req_desc_3_axuser_0_reg[i] <= uc2rb_rd_req_desc_3_axuser_0_reg[i];
             else 
               rd_req_desc_3_axuser_0_reg[i] <= rd_req_desc_3_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_1_reg_we[i])
               rd_req_desc_3_axuser_1_reg[i] <= uc2rb_rd_req_desc_3_axuser_1_reg[i];
             else 
               rd_req_desc_3_axuser_1_reg[i] <= rd_req_desc_3_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_2_reg_we[i])
               rd_req_desc_3_axuser_2_reg[i] <= uc2rb_rd_req_desc_3_axuser_2_reg[i];
             else 
               rd_req_desc_3_axuser_2_reg[i] <= rd_req_desc_3_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_3_reg_we[i])
               rd_req_desc_3_axuser_3_reg[i] <= uc2rb_rd_req_desc_3_axuser_3_reg[i];
             else 
               rd_req_desc_3_axuser_3_reg[i] <= rd_req_desc_3_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_4_reg_we[i])
               rd_req_desc_3_axuser_4_reg[i] <= uc2rb_rd_req_desc_3_axuser_4_reg[i];
             else 
               rd_req_desc_3_axuser_4_reg[i] <= rd_req_desc_3_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_5_reg_we[i])
               rd_req_desc_3_axuser_5_reg[i] <= uc2rb_rd_req_desc_3_axuser_5_reg[i];
             else 
               rd_req_desc_3_axuser_5_reg[i] <= rd_req_desc_3_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_6_reg_we[i])
               rd_req_desc_3_axuser_6_reg[i] <= uc2rb_rd_req_desc_3_axuser_6_reg[i];
             else 
               rd_req_desc_3_axuser_6_reg[i] <= rd_req_desc_3_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_7_reg_we[i])
               rd_req_desc_3_axuser_7_reg[i] <= uc2rb_rd_req_desc_3_axuser_7_reg[i];
             else 
               rd_req_desc_3_axuser_7_reg[i] <= rd_req_desc_3_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_8_reg_we[i])
               rd_req_desc_3_axuser_8_reg[i] <= uc2rb_rd_req_desc_3_axuser_8_reg[i];
             else 
               rd_req_desc_3_axuser_8_reg[i] <= rd_req_desc_3_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_9_reg_we[i])
               rd_req_desc_3_axuser_9_reg[i] <= uc2rb_rd_req_desc_3_axuser_9_reg[i];
             else 
               rd_req_desc_3_axuser_9_reg[i] <= rd_req_desc_3_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_10_reg_we[i])
               rd_req_desc_3_axuser_10_reg[i] <= uc2rb_rd_req_desc_3_axuser_10_reg[i];
             else 
               rd_req_desc_3_axuser_10_reg[i] <= rd_req_desc_3_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_11_reg_we[i])
               rd_req_desc_3_axuser_11_reg[i] <= uc2rb_rd_req_desc_3_axuser_11_reg[i];
             else 
               rd_req_desc_3_axuser_11_reg[i] <= rd_req_desc_3_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_12_reg_we[i])
               rd_req_desc_3_axuser_12_reg[i] <= uc2rb_rd_req_desc_3_axuser_12_reg[i];
             else 
               rd_req_desc_3_axuser_12_reg[i] <= rd_req_desc_3_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_13_reg_we[i])
               rd_req_desc_3_axuser_13_reg[i] <= uc2rb_rd_req_desc_3_axuser_13_reg[i];
             else 
               rd_req_desc_3_axuser_13_reg[i] <= rd_req_desc_3_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_14_reg_we[i])
               rd_req_desc_3_axuser_14_reg[i] <= uc2rb_rd_req_desc_3_axuser_14_reg[i];
             else 
               rd_req_desc_3_axuser_14_reg[i] <= rd_req_desc_3_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_3_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_3_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_3_axuser_15_reg_we[i])
               rd_req_desc_3_axuser_15_reg[i] <= uc2rb_rd_req_desc_3_axuser_15_reg[i];
             else 
               rd_req_desc_3_axuser_15_reg[i] <= rd_req_desc_3_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_3_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_txn_type_reg_we[i])
               wr_req_desc_3_txn_type_reg[i] <= uc2rb_wr_req_desc_3_txn_type_reg[i];
             else 
               wr_req_desc_3_txn_type_reg[i] <= wr_req_desc_3_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_3_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_size_reg_we[i])
               wr_req_desc_3_size_reg[i] <= uc2rb_wr_req_desc_3_size_reg[i];
             else 
               wr_req_desc_3_size_reg[i] <= wr_req_desc_3_size_reg[i];
        end
     end
   //WR_REQ_DESC_3_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_data_offset_reg_we[i])
               wr_req_desc_3_data_offset_reg[i] <= uc2rb_wr_req_desc_3_data_offset_reg[i];
             else 
               wr_req_desc_3_data_offset_reg[i] <= wr_req_desc_3_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axsize_reg_we[i])
               wr_req_desc_3_axsize_reg[i] <= uc2rb_wr_req_desc_3_axsize_reg[i];
             else 
               wr_req_desc_3_axsize_reg[i] <= wr_req_desc_3_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_3_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_attr_reg_we[i])
               wr_req_desc_3_attr_reg[i] <= uc2rb_wr_req_desc_3_attr_reg[i];
             else 
               wr_req_desc_3_attr_reg[i] <= wr_req_desc_3_attr_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axaddr_0_reg_we[i])
               wr_req_desc_3_axaddr_0_reg[i] <= uc2rb_wr_req_desc_3_axaddr_0_reg[i];
             else 
               wr_req_desc_3_axaddr_0_reg[i] <= wr_req_desc_3_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axaddr_1_reg_we[i])
               wr_req_desc_3_axaddr_1_reg[i] <= uc2rb_wr_req_desc_3_axaddr_1_reg[i];
             else 
               wr_req_desc_3_axaddr_1_reg[i] <= wr_req_desc_3_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axaddr_2_reg_we[i])
               wr_req_desc_3_axaddr_2_reg[i] <= uc2rb_wr_req_desc_3_axaddr_2_reg[i];
             else 
               wr_req_desc_3_axaddr_2_reg[i] <= wr_req_desc_3_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axaddr_3_reg_we[i])
               wr_req_desc_3_axaddr_3_reg[i] <= uc2rb_wr_req_desc_3_axaddr_3_reg[i];
             else 
               wr_req_desc_3_axaddr_3_reg[i] <= wr_req_desc_3_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axid_0_reg_we[i])
               wr_req_desc_3_axid_0_reg[i] <= uc2rb_wr_req_desc_3_axid_0_reg[i];
             else 
               wr_req_desc_3_axid_0_reg[i] <= wr_req_desc_3_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axid_1_reg_we[i])
               wr_req_desc_3_axid_1_reg[i] <= uc2rb_wr_req_desc_3_axid_1_reg[i];
             else 
               wr_req_desc_3_axid_1_reg[i] <= wr_req_desc_3_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axid_2_reg_we[i])
               wr_req_desc_3_axid_2_reg[i] <= uc2rb_wr_req_desc_3_axid_2_reg[i];
             else 
               wr_req_desc_3_axid_2_reg[i] <= wr_req_desc_3_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axid_3_reg_we[i])
               wr_req_desc_3_axid_3_reg[i] <= uc2rb_wr_req_desc_3_axid_3_reg[i];
             else 
               wr_req_desc_3_axid_3_reg[i] <= wr_req_desc_3_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_0_reg_we[i])
               wr_req_desc_3_axuser_0_reg[i] <= uc2rb_wr_req_desc_3_axuser_0_reg[i];
             else 
               wr_req_desc_3_axuser_0_reg[i] <= wr_req_desc_3_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_1_reg_we[i])
               wr_req_desc_3_axuser_1_reg[i] <= uc2rb_wr_req_desc_3_axuser_1_reg[i];
             else 
               wr_req_desc_3_axuser_1_reg[i] <= wr_req_desc_3_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_2_reg_we[i])
               wr_req_desc_3_axuser_2_reg[i] <= uc2rb_wr_req_desc_3_axuser_2_reg[i];
             else 
               wr_req_desc_3_axuser_2_reg[i] <= wr_req_desc_3_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_3_reg_we[i])
               wr_req_desc_3_axuser_3_reg[i] <= uc2rb_wr_req_desc_3_axuser_3_reg[i];
             else 
               wr_req_desc_3_axuser_3_reg[i] <= wr_req_desc_3_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_4_reg_we[i])
               wr_req_desc_3_axuser_4_reg[i] <= uc2rb_wr_req_desc_3_axuser_4_reg[i];
             else 
               wr_req_desc_3_axuser_4_reg[i] <= wr_req_desc_3_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_5_reg_we[i])
               wr_req_desc_3_axuser_5_reg[i] <= uc2rb_wr_req_desc_3_axuser_5_reg[i];
             else 
               wr_req_desc_3_axuser_5_reg[i] <= wr_req_desc_3_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_6_reg_we[i])
               wr_req_desc_3_axuser_6_reg[i] <= uc2rb_wr_req_desc_3_axuser_6_reg[i];
             else 
               wr_req_desc_3_axuser_6_reg[i] <= wr_req_desc_3_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_7_reg_we[i])
               wr_req_desc_3_axuser_7_reg[i] <= uc2rb_wr_req_desc_3_axuser_7_reg[i];
             else 
               wr_req_desc_3_axuser_7_reg[i] <= wr_req_desc_3_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_8_reg_we[i])
               wr_req_desc_3_axuser_8_reg[i] <= uc2rb_wr_req_desc_3_axuser_8_reg[i];
             else 
               wr_req_desc_3_axuser_8_reg[i] <= wr_req_desc_3_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_9_reg_we[i])
               wr_req_desc_3_axuser_9_reg[i] <= uc2rb_wr_req_desc_3_axuser_9_reg[i];
             else 
               wr_req_desc_3_axuser_9_reg[i] <= wr_req_desc_3_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_10_reg_we[i])
               wr_req_desc_3_axuser_10_reg[i] <= uc2rb_wr_req_desc_3_axuser_10_reg[i];
             else 
               wr_req_desc_3_axuser_10_reg[i] <= wr_req_desc_3_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_11_reg_we[i])
               wr_req_desc_3_axuser_11_reg[i] <= uc2rb_wr_req_desc_3_axuser_11_reg[i];
             else 
               wr_req_desc_3_axuser_11_reg[i] <= wr_req_desc_3_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_12_reg_we[i])
               wr_req_desc_3_axuser_12_reg[i] <= uc2rb_wr_req_desc_3_axuser_12_reg[i];
             else 
               wr_req_desc_3_axuser_12_reg[i] <= wr_req_desc_3_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_13_reg_we[i])
               wr_req_desc_3_axuser_13_reg[i] <= uc2rb_wr_req_desc_3_axuser_13_reg[i];
             else 
               wr_req_desc_3_axuser_13_reg[i] <= wr_req_desc_3_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_14_reg_we[i])
               wr_req_desc_3_axuser_14_reg[i] <= uc2rb_wr_req_desc_3_axuser_14_reg[i];
             else 
               wr_req_desc_3_axuser_14_reg[i] <= wr_req_desc_3_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_3_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_axuser_15_reg_we[i])
               wr_req_desc_3_axuser_15_reg[i] <= uc2rb_wr_req_desc_3_axuser_15_reg[i];
             else 
               wr_req_desc_3_axuser_15_reg[i] <= wr_req_desc_3_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_0_reg_we[i])
               wr_req_desc_3_wuser_0_reg[i] <= uc2rb_wr_req_desc_3_wuser_0_reg[i];
             else 
               wr_req_desc_3_wuser_0_reg[i] <= wr_req_desc_3_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_1_reg_we[i])
               wr_req_desc_3_wuser_1_reg[i] <= uc2rb_wr_req_desc_3_wuser_1_reg[i];
             else 
               wr_req_desc_3_wuser_1_reg[i] <= wr_req_desc_3_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_2_reg_we[i])
               wr_req_desc_3_wuser_2_reg[i] <= uc2rb_wr_req_desc_3_wuser_2_reg[i];
             else 
               wr_req_desc_3_wuser_2_reg[i] <= wr_req_desc_3_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_3_reg_we[i])
               wr_req_desc_3_wuser_3_reg[i] <= uc2rb_wr_req_desc_3_wuser_3_reg[i];
             else 
               wr_req_desc_3_wuser_3_reg[i] <= wr_req_desc_3_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_4_reg_we[i])
               wr_req_desc_3_wuser_4_reg[i] <= uc2rb_wr_req_desc_3_wuser_4_reg[i];
             else 
               wr_req_desc_3_wuser_4_reg[i] <= wr_req_desc_3_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_5_reg_we[i])
               wr_req_desc_3_wuser_5_reg[i] <= uc2rb_wr_req_desc_3_wuser_5_reg[i];
             else 
               wr_req_desc_3_wuser_5_reg[i] <= wr_req_desc_3_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_6_reg_we[i])
               wr_req_desc_3_wuser_6_reg[i] <= uc2rb_wr_req_desc_3_wuser_6_reg[i];
             else 
               wr_req_desc_3_wuser_6_reg[i] <= wr_req_desc_3_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_7_reg_we[i])
               wr_req_desc_3_wuser_7_reg[i] <= uc2rb_wr_req_desc_3_wuser_7_reg[i];
             else 
               wr_req_desc_3_wuser_7_reg[i] <= wr_req_desc_3_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_8_reg_we[i])
               wr_req_desc_3_wuser_8_reg[i] <= uc2rb_wr_req_desc_3_wuser_8_reg[i];
             else 
               wr_req_desc_3_wuser_8_reg[i] <= wr_req_desc_3_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_9_reg_we[i])
               wr_req_desc_3_wuser_9_reg[i] <= uc2rb_wr_req_desc_3_wuser_9_reg[i];
             else 
               wr_req_desc_3_wuser_9_reg[i] <= wr_req_desc_3_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_10_reg_we[i])
               wr_req_desc_3_wuser_10_reg[i] <= uc2rb_wr_req_desc_3_wuser_10_reg[i];
             else 
               wr_req_desc_3_wuser_10_reg[i] <= wr_req_desc_3_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_11_reg_we[i])
               wr_req_desc_3_wuser_11_reg[i] <= uc2rb_wr_req_desc_3_wuser_11_reg[i];
             else 
               wr_req_desc_3_wuser_11_reg[i] <= wr_req_desc_3_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_12_reg_we[i])
               wr_req_desc_3_wuser_12_reg[i] <= uc2rb_wr_req_desc_3_wuser_12_reg[i];
             else 
               wr_req_desc_3_wuser_12_reg[i] <= wr_req_desc_3_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_13_reg_we[i])
               wr_req_desc_3_wuser_13_reg[i] <= uc2rb_wr_req_desc_3_wuser_13_reg[i];
             else 
               wr_req_desc_3_wuser_13_reg[i] <= wr_req_desc_3_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_14_reg_we[i])
               wr_req_desc_3_wuser_14_reg[i] <= uc2rb_wr_req_desc_3_wuser_14_reg[i];
             else 
               wr_req_desc_3_wuser_14_reg[i] <= wr_req_desc_3_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_3_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_3_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_3_wuser_15_reg_we[i])
               wr_req_desc_3_wuser_15_reg[i] <= uc2rb_wr_req_desc_3_wuser_15_reg[i];
             else 
               wr_req_desc_3_wuser_15_reg[i] <= wr_req_desc_3_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_3_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_3_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_3_resp_reg_we[i])
               sn_resp_desc_3_resp_reg[i] <= uc2rb_sn_resp_desc_3_resp_reg[i];
             else 
               sn_resp_desc_3_resp_reg[i] <= sn_resp_desc_3_resp_reg[i];
        end
     end
   //RD_REQ_DESC_4_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_txn_type_reg_we[i])
               rd_req_desc_4_txn_type_reg[i] <= uc2rb_rd_req_desc_4_txn_type_reg[i];
             else 
               rd_req_desc_4_txn_type_reg[i] <= rd_req_desc_4_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_4_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_size_reg_we[i])
               rd_req_desc_4_size_reg[i] <= uc2rb_rd_req_desc_4_size_reg[i];
             else 
               rd_req_desc_4_size_reg[i] <= rd_req_desc_4_size_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axsize_reg_we[i])
               rd_req_desc_4_axsize_reg[i] <= uc2rb_rd_req_desc_4_axsize_reg[i];
             else 
               rd_req_desc_4_axsize_reg[i] <= rd_req_desc_4_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_4_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_attr_reg_we[i])
               rd_req_desc_4_attr_reg[i] <= uc2rb_rd_req_desc_4_attr_reg[i];
             else 
               rd_req_desc_4_attr_reg[i] <= rd_req_desc_4_attr_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axaddr_0_reg_we[i])
               rd_req_desc_4_axaddr_0_reg[i] <= uc2rb_rd_req_desc_4_axaddr_0_reg[i];
             else 
               rd_req_desc_4_axaddr_0_reg[i] <= rd_req_desc_4_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axaddr_1_reg_we[i])
               rd_req_desc_4_axaddr_1_reg[i] <= uc2rb_rd_req_desc_4_axaddr_1_reg[i];
             else 
               rd_req_desc_4_axaddr_1_reg[i] <= rd_req_desc_4_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axaddr_2_reg_we[i])
               rd_req_desc_4_axaddr_2_reg[i] <= uc2rb_rd_req_desc_4_axaddr_2_reg[i];
             else 
               rd_req_desc_4_axaddr_2_reg[i] <= rd_req_desc_4_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axaddr_3_reg_we[i])
               rd_req_desc_4_axaddr_3_reg[i] <= uc2rb_rd_req_desc_4_axaddr_3_reg[i];
             else 
               rd_req_desc_4_axaddr_3_reg[i] <= rd_req_desc_4_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axid_0_reg_we[i])
               rd_req_desc_4_axid_0_reg[i] <= uc2rb_rd_req_desc_4_axid_0_reg[i];
             else 
               rd_req_desc_4_axid_0_reg[i] <= rd_req_desc_4_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axid_1_reg_we[i])
               rd_req_desc_4_axid_1_reg[i] <= uc2rb_rd_req_desc_4_axid_1_reg[i];
             else 
               rd_req_desc_4_axid_1_reg[i] <= rd_req_desc_4_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axid_2_reg_we[i])
               rd_req_desc_4_axid_2_reg[i] <= uc2rb_rd_req_desc_4_axid_2_reg[i];
             else 
               rd_req_desc_4_axid_2_reg[i] <= rd_req_desc_4_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axid_3_reg_we[i])
               rd_req_desc_4_axid_3_reg[i] <= uc2rb_rd_req_desc_4_axid_3_reg[i];
             else 
               rd_req_desc_4_axid_3_reg[i] <= rd_req_desc_4_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_0_reg_we[i])
               rd_req_desc_4_axuser_0_reg[i] <= uc2rb_rd_req_desc_4_axuser_0_reg[i];
             else 
               rd_req_desc_4_axuser_0_reg[i] <= rd_req_desc_4_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_1_reg_we[i])
               rd_req_desc_4_axuser_1_reg[i] <= uc2rb_rd_req_desc_4_axuser_1_reg[i];
             else 
               rd_req_desc_4_axuser_1_reg[i] <= rd_req_desc_4_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_2_reg_we[i])
               rd_req_desc_4_axuser_2_reg[i] <= uc2rb_rd_req_desc_4_axuser_2_reg[i];
             else 
               rd_req_desc_4_axuser_2_reg[i] <= rd_req_desc_4_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_3_reg_we[i])
               rd_req_desc_4_axuser_3_reg[i] <= uc2rb_rd_req_desc_4_axuser_3_reg[i];
             else 
               rd_req_desc_4_axuser_3_reg[i] <= rd_req_desc_4_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_4_reg_we[i])
               rd_req_desc_4_axuser_4_reg[i] <= uc2rb_rd_req_desc_4_axuser_4_reg[i];
             else 
               rd_req_desc_4_axuser_4_reg[i] <= rd_req_desc_4_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_5_reg_we[i])
               rd_req_desc_4_axuser_5_reg[i] <= uc2rb_rd_req_desc_4_axuser_5_reg[i];
             else 
               rd_req_desc_4_axuser_5_reg[i] <= rd_req_desc_4_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_6_reg_we[i])
               rd_req_desc_4_axuser_6_reg[i] <= uc2rb_rd_req_desc_4_axuser_6_reg[i];
             else 
               rd_req_desc_4_axuser_6_reg[i] <= rd_req_desc_4_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_7_reg_we[i])
               rd_req_desc_4_axuser_7_reg[i] <= uc2rb_rd_req_desc_4_axuser_7_reg[i];
             else 
               rd_req_desc_4_axuser_7_reg[i] <= rd_req_desc_4_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_8_reg_we[i])
               rd_req_desc_4_axuser_8_reg[i] <= uc2rb_rd_req_desc_4_axuser_8_reg[i];
             else 
               rd_req_desc_4_axuser_8_reg[i] <= rd_req_desc_4_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_9_reg_we[i])
               rd_req_desc_4_axuser_9_reg[i] <= uc2rb_rd_req_desc_4_axuser_9_reg[i];
             else 
               rd_req_desc_4_axuser_9_reg[i] <= rd_req_desc_4_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_10_reg_we[i])
               rd_req_desc_4_axuser_10_reg[i] <= uc2rb_rd_req_desc_4_axuser_10_reg[i];
             else 
               rd_req_desc_4_axuser_10_reg[i] <= rd_req_desc_4_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_11_reg_we[i])
               rd_req_desc_4_axuser_11_reg[i] <= uc2rb_rd_req_desc_4_axuser_11_reg[i];
             else 
               rd_req_desc_4_axuser_11_reg[i] <= rd_req_desc_4_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_12_reg_we[i])
               rd_req_desc_4_axuser_12_reg[i] <= uc2rb_rd_req_desc_4_axuser_12_reg[i];
             else 
               rd_req_desc_4_axuser_12_reg[i] <= rd_req_desc_4_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_13_reg_we[i])
               rd_req_desc_4_axuser_13_reg[i] <= uc2rb_rd_req_desc_4_axuser_13_reg[i];
             else 
               rd_req_desc_4_axuser_13_reg[i] <= rd_req_desc_4_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_14_reg_we[i])
               rd_req_desc_4_axuser_14_reg[i] <= uc2rb_rd_req_desc_4_axuser_14_reg[i];
             else 
               rd_req_desc_4_axuser_14_reg[i] <= rd_req_desc_4_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_4_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_4_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_4_axuser_15_reg_we[i])
               rd_req_desc_4_axuser_15_reg[i] <= uc2rb_rd_req_desc_4_axuser_15_reg[i];
             else 
               rd_req_desc_4_axuser_15_reg[i] <= rd_req_desc_4_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_4_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_txn_type_reg_we[i])
               wr_req_desc_4_txn_type_reg[i] <= uc2rb_wr_req_desc_4_txn_type_reg[i];
             else 
               wr_req_desc_4_txn_type_reg[i] <= wr_req_desc_4_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_4_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_size_reg_we[i])
               wr_req_desc_4_size_reg[i] <= uc2rb_wr_req_desc_4_size_reg[i];
             else 
               wr_req_desc_4_size_reg[i] <= wr_req_desc_4_size_reg[i];
        end
     end
   //WR_REQ_DESC_4_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_data_offset_reg_we[i])
               wr_req_desc_4_data_offset_reg[i] <= uc2rb_wr_req_desc_4_data_offset_reg[i];
             else 
               wr_req_desc_4_data_offset_reg[i] <= wr_req_desc_4_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axsize_reg_we[i])
               wr_req_desc_4_axsize_reg[i] <= uc2rb_wr_req_desc_4_axsize_reg[i];
             else 
               wr_req_desc_4_axsize_reg[i] <= wr_req_desc_4_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_4_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_attr_reg_we[i])
               wr_req_desc_4_attr_reg[i] <= uc2rb_wr_req_desc_4_attr_reg[i];
             else 
               wr_req_desc_4_attr_reg[i] <= wr_req_desc_4_attr_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axaddr_0_reg_we[i])
               wr_req_desc_4_axaddr_0_reg[i] <= uc2rb_wr_req_desc_4_axaddr_0_reg[i];
             else 
               wr_req_desc_4_axaddr_0_reg[i] <= wr_req_desc_4_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axaddr_1_reg_we[i])
               wr_req_desc_4_axaddr_1_reg[i] <= uc2rb_wr_req_desc_4_axaddr_1_reg[i];
             else 
               wr_req_desc_4_axaddr_1_reg[i] <= wr_req_desc_4_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axaddr_2_reg_we[i])
               wr_req_desc_4_axaddr_2_reg[i] <= uc2rb_wr_req_desc_4_axaddr_2_reg[i];
             else 
               wr_req_desc_4_axaddr_2_reg[i] <= wr_req_desc_4_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axaddr_3_reg_we[i])
               wr_req_desc_4_axaddr_3_reg[i] <= uc2rb_wr_req_desc_4_axaddr_3_reg[i];
             else 
               wr_req_desc_4_axaddr_3_reg[i] <= wr_req_desc_4_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axid_0_reg_we[i])
               wr_req_desc_4_axid_0_reg[i] <= uc2rb_wr_req_desc_4_axid_0_reg[i];
             else 
               wr_req_desc_4_axid_0_reg[i] <= wr_req_desc_4_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axid_1_reg_we[i])
               wr_req_desc_4_axid_1_reg[i] <= uc2rb_wr_req_desc_4_axid_1_reg[i];
             else 
               wr_req_desc_4_axid_1_reg[i] <= wr_req_desc_4_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axid_2_reg_we[i])
               wr_req_desc_4_axid_2_reg[i] <= uc2rb_wr_req_desc_4_axid_2_reg[i];
             else 
               wr_req_desc_4_axid_2_reg[i] <= wr_req_desc_4_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axid_3_reg_we[i])
               wr_req_desc_4_axid_3_reg[i] <= uc2rb_wr_req_desc_4_axid_3_reg[i];
             else 
               wr_req_desc_4_axid_3_reg[i] <= wr_req_desc_4_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_0_reg_we[i])
               wr_req_desc_4_axuser_0_reg[i] <= uc2rb_wr_req_desc_4_axuser_0_reg[i];
             else 
               wr_req_desc_4_axuser_0_reg[i] <= wr_req_desc_4_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_1_reg_we[i])
               wr_req_desc_4_axuser_1_reg[i] <= uc2rb_wr_req_desc_4_axuser_1_reg[i];
             else 
               wr_req_desc_4_axuser_1_reg[i] <= wr_req_desc_4_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_2_reg_we[i])
               wr_req_desc_4_axuser_2_reg[i] <= uc2rb_wr_req_desc_4_axuser_2_reg[i];
             else 
               wr_req_desc_4_axuser_2_reg[i] <= wr_req_desc_4_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_3_reg_we[i])
               wr_req_desc_4_axuser_3_reg[i] <= uc2rb_wr_req_desc_4_axuser_3_reg[i];
             else 
               wr_req_desc_4_axuser_3_reg[i] <= wr_req_desc_4_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_4_reg_we[i])
               wr_req_desc_4_axuser_4_reg[i] <= uc2rb_wr_req_desc_4_axuser_4_reg[i];
             else 
               wr_req_desc_4_axuser_4_reg[i] <= wr_req_desc_4_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_5_reg_we[i])
               wr_req_desc_4_axuser_5_reg[i] <= uc2rb_wr_req_desc_4_axuser_5_reg[i];
             else 
               wr_req_desc_4_axuser_5_reg[i] <= wr_req_desc_4_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_6_reg_we[i])
               wr_req_desc_4_axuser_6_reg[i] <= uc2rb_wr_req_desc_4_axuser_6_reg[i];
             else 
               wr_req_desc_4_axuser_6_reg[i] <= wr_req_desc_4_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_7_reg_we[i])
               wr_req_desc_4_axuser_7_reg[i] <= uc2rb_wr_req_desc_4_axuser_7_reg[i];
             else 
               wr_req_desc_4_axuser_7_reg[i] <= wr_req_desc_4_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_8_reg_we[i])
               wr_req_desc_4_axuser_8_reg[i] <= uc2rb_wr_req_desc_4_axuser_8_reg[i];
             else 
               wr_req_desc_4_axuser_8_reg[i] <= wr_req_desc_4_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_9_reg_we[i])
               wr_req_desc_4_axuser_9_reg[i] <= uc2rb_wr_req_desc_4_axuser_9_reg[i];
             else 
               wr_req_desc_4_axuser_9_reg[i] <= wr_req_desc_4_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_10_reg_we[i])
               wr_req_desc_4_axuser_10_reg[i] <= uc2rb_wr_req_desc_4_axuser_10_reg[i];
             else 
               wr_req_desc_4_axuser_10_reg[i] <= wr_req_desc_4_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_11_reg_we[i])
               wr_req_desc_4_axuser_11_reg[i] <= uc2rb_wr_req_desc_4_axuser_11_reg[i];
             else 
               wr_req_desc_4_axuser_11_reg[i] <= wr_req_desc_4_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_12_reg_we[i])
               wr_req_desc_4_axuser_12_reg[i] <= uc2rb_wr_req_desc_4_axuser_12_reg[i];
             else 
               wr_req_desc_4_axuser_12_reg[i] <= wr_req_desc_4_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_13_reg_we[i])
               wr_req_desc_4_axuser_13_reg[i] <= uc2rb_wr_req_desc_4_axuser_13_reg[i];
             else 
               wr_req_desc_4_axuser_13_reg[i] <= wr_req_desc_4_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_14_reg_we[i])
               wr_req_desc_4_axuser_14_reg[i] <= uc2rb_wr_req_desc_4_axuser_14_reg[i];
             else 
               wr_req_desc_4_axuser_14_reg[i] <= wr_req_desc_4_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_4_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_axuser_15_reg_we[i])
               wr_req_desc_4_axuser_15_reg[i] <= uc2rb_wr_req_desc_4_axuser_15_reg[i];
             else 
               wr_req_desc_4_axuser_15_reg[i] <= wr_req_desc_4_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_0_reg_we[i])
               wr_req_desc_4_wuser_0_reg[i] <= uc2rb_wr_req_desc_4_wuser_0_reg[i];
             else 
               wr_req_desc_4_wuser_0_reg[i] <= wr_req_desc_4_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_1_reg_we[i])
               wr_req_desc_4_wuser_1_reg[i] <= uc2rb_wr_req_desc_4_wuser_1_reg[i];
             else 
               wr_req_desc_4_wuser_1_reg[i] <= wr_req_desc_4_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_2_reg_we[i])
               wr_req_desc_4_wuser_2_reg[i] <= uc2rb_wr_req_desc_4_wuser_2_reg[i];
             else 
               wr_req_desc_4_wuser_2_reg[i] <= wr_req_desc_4_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_3_reg_we[i])
               wr_req_desc_4_wuser_3_reg[i] <= uc2rb_wr_req_desc_4_wuser_3_reg[i];
             else 
               wr_req_desc_4_wuser_3_reg[i] <= wr_req_desc_4_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_4_reg_we[i])
               wr_req_desc_4_wuser_4_reg[i] <= uc2rb_wr_req_desc_4_wuser_4_reg[i];
             else 
               wr_req_desc_4_wuser_4_reg[i] <= wr_req_desc_4_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_5_reg_we[i])
               wr_req_desc_4_wuser_5_reg[i] <= uc2rb_wr_req_desc_4_wuser_5_reg[i];
             else 
               wr_req_desc_4_wuser_5_reg[i] <= wr_req_desc_4_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_6_reg_we[i])
               wr_req_desc_4_wuser_6_reg[i] <= uc2rb_wr_req_desc_4_wuser_6_reg[i];
             else 
               wr_req_desc_4_wuser_6_reg[i] <= wr_req_desc_4_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_7_reg_we[i])
               wr_req_desc_4_wuser_7_reg[i] <= uc2rb_wr_req_desc_4_wuser_7_reg[i];
             else 
               wr_req_desc_4_wuser_7_reg[i] <= wr_req_desc_4_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_8_reg_we[i])
               wr_req_desc_4_wuser_8_reg[i] <= uc2rb_wr_req_desc_4_wuser_8_reg[i];
             else 
               wr_req_desc_4_wuser_8_reg[i] <= wr_req_desc_4_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_9_reg_we[i])
               wr_req_desc_4_wuser_9_reg[i] <= uc2rb_wr_req_desc_4_wuser_9_reg[i];
             else 
               wr_req_desc_4_wuser_9_reg[i] <= wr_req_desc_4_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_10_reg_we[i])
               wr_req_desc_4_wuser_10_reg[i] <= uc2rb_wr_req_desc_4_wuser_10_reg[i];
             else 
               wr_req_desc_4_wuser_10_reg[i] <= wr_req_desc_4_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_11_reg_we[i])
               wr_req_desc_4_wuser_11_reg[i] <= uc2rb_wr_req_desc_4_wuser_11_reg[i];
             else 
               wr_req_desc_4_wuser_11_reg[i] <= wr_req_desc_4_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_12_reg_we[i])
               wr_req_desc_4_wuser_12_reg[i] <= uc2rb_wr_req_desc_4_wuser_12_reg[i];
             else 
               wr_req_desc_4_wuser_12_reg[i] <= wr_req_desc_4_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_13_reg_we[i])
               wr_req_desc_4_wuser_13_reg[i] <= uc2rb_wr_req_desc_4_wuser_13_reg[i];
             else 
               wr_req_desc_4_wuser_13_reg[i] <= wr_req_desc_4_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_14_reg_we[i])
               wr_req_desc_4_wuser_14_reg[i] <= uc2rb_wr_req_desc_4_wuser_14_reg[i];
             else 
               wr_req_desc_4_wuser_14_reg[i] <= wr_req_desc_4_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_4_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_4_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_4_wuser_15_reg_we[i])
               wr_req_desc_4_wuser_15_reg[i] <= uc2rb_wr_req_desc_4_wuser_15_reg[i];
             else 
               wr_req_desc_4_wuser_15_reg[i] <= wr_req_desc_4_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_4_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_4_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_4_resp_reg_we[i])
               sn_resp_desc_4_resp_reg[i] <= uc2rb_sn_resp_desc_4_resp_reg[i];
             else 
               sn_resp_desc_4_resp_reg[i] <= sn_resp_desc_4_resp_reg[i];
        end
     end
   //RD_REQ_DESC_5_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_txn_type_reg_we[i])
               rd_req_desc_5_txn_type_reg[i] <= uc2rb_rd_req_desc_5_txn_type_reg[i];
             else 
               rd_req_desc_5_txn_type_reg[i] <= rd_req_desc_5_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_5_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_size_reg_we[i])
               rd_req_desc_5_size_reg[i] <= uc2rb_rd_req_desc_5_size_reg[i];
             else 
               rd_req_desc_5_size_reg[i] <= rd_req_desc_5_size_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axsize_reg_we[i])
               rd_req_desc_5_axsize_reg[i] <= uc2rb_rd_req_desc_5_axsize_reg[i];
             else 
               rd_req_desc_5_axsize_reg[i] <= rd_req_desc_5_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_5_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_attr_reg_we[i])
               rd_req_desc_5_attr_reg[i] <= uc2rb_rd_req_desc_5_attr_reg[i];
             else 
               rd_req_desc_5_attr_reg[i] <= rd_req_desc_5_attr_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axaddr_0_reg_we[i])
               rd_req_desc_5_axaddr_0_reg[i] <= uc2rb_rd_req_desc_5_axaddr_0_reg[i];
             else 
               rd_req_desc_5_axaddr_0_reg[i] <= rd_req_desc_5_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axaddr_1_reg_we[i])
               rd_req_desc_5_axaddr_1_reg[i] <= uc2rb_rd_req_desc_5_axaddr_1_reg[i];
             else 
               rd_req_desc_5_axaddr_1_reg[i] <= rd_req_desc_5_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axaddr_2_reg_we[i])
               rd_req_desc_5_axaddr_2_reg[i] <= uc2rb_rd_req_desc_5_axaddr_2_reg[i];
             else 
               rd_req_desc_5_axaddr_2_reg[i] <= rd_req_desc_5_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axaddr_3_reg_we[i])
               rd_req_desc_5_axaddr_3_reg[i] <= uc2rb_rd_req_desc_5_axaddr_3_reg[i];
             else 
               rd_req_desc_5_axaddr_3_reg[i] <= rd_req_desc_5_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axid_0_reg_we[i])
               rd_req_desc_5_axid_0_reg[i] <= uc2rb_rd_req_desc_5_axid_0_reg[i];
             else 
               rd_req_desc_5_axid_0_reg[i] <= rd_req_desc_5_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axid_1_reg_we[i])
               rd_req_desc_5_axid_1_reg[i] <= uc2rb_rd_req_desc_5_axid_1_reg[i];
             else 
               rd_req_desc_5_axid_1_reg[i] <= rd_req_desc_5_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axid_2_reg_we[i])
               rd_req_desc_5_axid_2_reg[i] <= uc2rb_rd_req_desc_5_axid_2_reg[i];
             else 
               rd_req_desc_5_axid_2_reg[i] <= rd_req_desc_5_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axid_3_reg_we[i])
               rd_req_desc_5_axid_3_reg[i] <= uc2rb_rd_req_desc_5_axid_3_reg[i];
             else 
               rd_req_desc_5_axid_3_reg[i] <= rd_req_desc_5_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_0_reg_we[i])
               rd_req_desc_5_axuser_0_reg[i] <= uc2rb_rd_req_desc_5_axuser_0_reg[i];
             else 
               rd_req_desc_5_axuser_0_reg[i] <= rd_req_desc_5_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_1_reg_we[i])
               rd_req_desc_5_axuser_1_reg[i] <= uc2rb_rd_req_desc_5_axuser_1_reg[i];
             else 
               rd_req_desc_5_axuser_1_reg[i] <= rd_req_desc_5_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_2_reg_we[i])
               rd_req_desc_5_axuser_2_reg[i] <= uc2rb_rd_req_desc_5_axuser_2_reg[i];
             else 
               rd_req_desc_5_axuser_2_reg[i] <= rd_req_desc_5_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_3_reg_we[i])
               rd_req_desc_5_axuser_3_reg[i] <= uc2rb_rd_req_desc_5_axuser_3_reg[i];
             else 
               rd_req_desc_5_axuser_3_reg[i] <= rd_req_desc_5_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_4_reg_we[i])
               rd_req_desc_5_axuser_4_reg[i] <= uc2rb_rd_req_desc_5_axuser_4_reg[i];
             else 
               rd_req_desc_5_axuser_4_reg[i] <= rd_req_desc_5_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_5_reg_we[i])
               rd_req_desc_5_axuser_5_reg[i] <= uc2rb_rd_req_desc_5_axuser_5_reg[i];
             else 
               rd_req_desc_5_axuser_5_reg[i] <= rd_req_desc_5_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_6_reg_we[i])
               rd_req_desc_5_axuser_6_reg[i] <= uc2rb_rd_req_desc_5_axuser_6_reg[i];
             else 
               rd_req_desc_5_axuser_6_reg[i] <= rd_req_desc_5_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_7_reg_we[i])
               rd_req_desc_5_axuser_7_reg[i] <= uc2rb_rd_req_desc_5_axuser_7_reg[i];
             else 
               rd_req_desc_5_axuser_7_reg[i] <= rd_req_desc_5_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_8_reg_we[i])
               rd_req_desc_5_axuser_8_reg[i] <= uc2rb_rd_req_desc_5_axuser_8_reg[i];
             else 
               rd_req_desc_5_axuser_8_reg[i] <= rd_req_desc_5_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_9_reg_we[i])
               rd_req_desc_5_axuser_9_reg[i] <= uc2rb_rd_req_desc_5_axuser_9_reg[i];
             else 
               rd_req_desc_5_axuser_9_reg[i] <= rd_req_desc_5_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_10_reg_we[i])
               rd_req_desc_5_axuser_10_reg[i] <= uc2rb_rd_req_desc_5_axuser_10_reg[i];
             else 
               rd_req_desc_5_axuser_10_reg[i] <= rd_req_desc_5_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_11_reg_we[i])
               rd_req_desc_5_axuser_11_reg[i] <= uc2rb_rd_req_desc_5_axuser_11_reg[i];
             else 
               rd_req_desc_5_axuser_11_reg[i] <= rd_req_desc_5_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_12_reg_we[i])
               rd_req_desc_5_axuser_12_reg[i] <= uc2rb_rd_req_desc_5_axuser_12_reg[i];
             else 
               rd_req_desc_5_axuser_12_reg[i] <= rd_req_desc_5_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_13_reg_we[i])
               rd_req_desc_5_axuser_13_reg[i] <= uc2rb_rd_req_desc_5_axuser_13_reg[i];
             else 
               rd_req_desc_5_axuser_13_reg[i] <= rd_req_desc_5_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_14_reg_we[i])
               rd_req_desc_5_axuser_14_reg[i] <= uc2rb_rd_req_desc_5_axuser_14_reg[i];
             else 
               rd_req_desc_5_axuser_14_reg[i] <= rd_req_desc_5_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_5_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_5_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_5_axuser_15_reg_we[i])
               rd_req_desc_5_axuser_15_reg[i] <= uc2rb_rd_req_desc_5_axuser_15_reg[i];
             else 
               rd_req_desc_5_axuser_15_reg[i] <= rd_req_desc_5_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_5_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_txn_type_reg_we[i])
               wr_req_desc_5_txn_type_reg[i] <= uc2rb_wr_req_desc_5_txn_type_reg[i];
             else 
               wr_req_desc_5_txn_type_reg[i] <= wr_req_desc_5_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_5_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_size_reg_we[i])
               wr_req_desc_5_size_reg[i] <= uc2rb_wr_req_desc_5_size_reg[i];
             else 
               wr_req_desc_5_size_reg[i] <= wr_req_desc_5_size_reg[i];
        end
     end
   //WR_REQ_DESC_5_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_data_offset_reg_we[i])
               wr_req_desc_5_data_offset_reg[i] <= uc2rb_wr_req_desc_5_data_offset_reg[i];
             else 
               wr_req_desc_5_data_offset_reg[i] <= wr_req_desc_5_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axsize_reg_we[i])
               wr_req_desc_5_axsize_reg[i] <= uc2rb_wr_req_desc_5_axsize_reg[i];
             else 
               wr_req_desc_5_axsize_reg[i] <= wr_req_desc_5_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_5_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_attr_reg_we[i])
               wr_req_desc_5_attr_reg[i] <= uc2rb_wr_req_desc_5_attr_reg[i];
             else 
               wr_req_desc_5_attr_reg[i] <= wr_req_desc_5_attr_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axaddr_0_reg_we[i])
               wr_req_desc_5_axaddr_0_reg[i] <= uc2rb_wr_req_desc_5_axaddr_0_reg[i];
             else 
               wr_req_desc_5_axaddr_0_reg[i] <= wr_req_desc_5_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axaddr_1_reg_we[i])
               wr_req_desc_5_axaddr_1_reg[i] <= uc2rb_wr_req_desc_5_axaddr_1_reg[i];
             else 
               wr_req_desc_5_axaddr_1_reg[i] <= wr_req_desc_5_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axaddr_2_reg_we[i])
               wr_req_desc_5_axaddr_2_reg[i] <= uc2rb_wr_req_desc_5_axaddr_2_reg[i];
             else 
               wr_req_desc_5_axaddr_2_reg[i] <= wr_req_desc_5_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axaddr_3_reg_we[i])
               wr_req_desc_5_axaddr_3_reg[i] <= uc2rb_wr_req_desc_5_axaddr_3_reg[i];
             else 
               wr_req_desc_5_axaddr_3_reg[i] <= wr_req_desc_5_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axid_0_reg_we[i])
               wr_req_desc_5_axid_0_reg[i] <= uc2rb_wr_req_desc_5_axid_0_reg[i];
             else 
               wr_req_desc_5_axid_0_reg[i] <= wr_req_desc_5_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axid_1_reg_we[i])
               wr_req_desc_5_axid_1_reg[i] <= uc2rb_wr_req_desc_5_axid_1_reg[i];
             else 
               wr_req_desc_5_axid_1_reg[i] <= wr_req_desc_5_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axid_2_reg_we[i])
               wr_req_desc_5_axid_2_reg[i] <= uc2rb_wr_req_desc_5_axid_2_reg[i];
             else 
               wr_req_desc_5_axid_2_reg[i] <= wr_req_desc_5_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axid_3_reg_we[i])
               wr_req_desc_5_axid_3_reg[i] <= uc2rb_wr_req_desc_5_axid_3_reg[i];
             else 
               wr_req_desc_5_axid_3_reg[i] <= wr_req_desc_5_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_0_reg_we[i])
               wr_req_desc_5_axuser_0_reg[i] <= uc2rb_wr_req_desc_5_axuser_0_reg[i];
             else 
               wr_req_desc_5_axuser_0_reg[i] <= wr_req_desc_5_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_1_reg_we[i])
               wr_req_desc_5_axuser_1_reg[i] <= uc2rb_wr_req_desc_5_axuser_1_reg[i];
             else 
               wr_req_desc_5_axuser_1_reg[i] <= wr_req_desc_5_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_2_reg_we[i])
               wr_req_desc_5_axuser_2_reg[i] <= uc2rb_wr_req_desc_5_axuser_2_reg[i];
             else 
               wr_req_desc_5_axuser_2_reg[i] <= wr_req_desc_5_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_3_reg_we[i])
               wr_req_desc_5_axuser_3_reg[i] <= uc2rb_wr_req_desc_5_axuser_3_reg[i];
             else 
               wr_req_desc_5_axuser_3_reg[i] <= wr_req_desc_5_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_4_reg_we[i])
               wr_req_desc_5_axuser_4_reg[i] <= uc2rb_wr_req_desc_5_axuser_4_reg[i];
             else 
               wr_req_desc_5_axuser_4_reg[i] <= wr_req_desc_5_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_5_reg_we[i])
               wr_req_desc_5_axuser_5_reg[i] <= uc2rb_wr_req_desc_5_axuser_5_reg[i];
             else 
               wr_req_desc_5_axuser_5_reg[i] <= wr_req_desc_5_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_6_reg_we[i])
               wr_req_desc_5_axuser_6_reg[i] <= uc2rb_wr_req_desc_5_axuser_6_reg[i];
             else 
               wr_req_desc_5_axuser_6_reg[i] <= wr_req_desc_5_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_7_reg_we[i])
               wr_req_desc_5_axuser_7_reg[i] <= uc2rb_wr_req_desc_5_axuser_7_reg[i];
             else 
               wr_req_desc_5_axuser_7_reg[i] <= wr_req_desc_5_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_8_reg_we[i])
               wr_req_desc_5_axuser_8_reg[i] <= uc2rb_wr_req_desc_5_axuser_8_reg[i];
             else 
               wr_req_desc_5_axuser_8_reg[i] <= wr_req_desc_5_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_9_reg_we[i])
               wr_req_desc_5_axuser_9_reg[i] <= uc2rb_wr_req_desc_5_axuser_9_reg[i];
             else 
               wr_req_desc_5_axuser_9_reg[i] <= wr_req_desc_5_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_10_reg_we[i])
               wr_req_desc_5_axuser_10_reg[i] <= uc2rb_wr_req_desc_5_axuser_10_reg[i];
             else 
               wr_req_desc_5_axuser_10_reg[i] <= wr_req_desc_5_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_11_reg_we[i])
               wr_req_desc_5_axuser_11_reg[i] <= uc2rb_wr_req_desc_5_axuser_11_reg[i];
             else 
               wr_req_desc_5_axuser_11_reg[i] <= wr_req_desc_5_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_12_reg_we[i])
               wr_req_desc_5_axuser_12_reg[i] <= uc2rb_wr_req_desc_5_axuser_12_reg[i];
             else 
               wr_req_desc_5_axuser_12_reg[i] <= wr_req_desc_5_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_13_reg_we[i])
               wr_req_desc_5_axuser_13_reg[i] <= uc2rb_wr_req_desc_5_axuser_13_reg[i];
             else 
               wr_req_desc_5_axuser_13_reg[i] <= wr_req_desc_5_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_14_reg_we[i])
               wr_req_desc_5_axuser_14_reg[i] <= uc2rb_wr_req_desc_5_axuser_14_reg[i];
             else 
               wr_req_desc_5_axuser_14_reg[i] <= wr_req_desc_5_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_5_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_axuser_15_reg_we[i])
               wr_req_desc_5_axuser_15_reg[i] <= uc2rb_wr_req_desc_5_axuser_15_reg[i];
             else 
               wr_req_desc_5_axuser_15_reg[i] <= wr_req_desc_5_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_0_reg_we[i])
               wr_req_desc_5_wuser_0_reg[i] <= uc2rb_wr_req_desc_5_wuser_0_reg[i];
             else 
               wr_req_desc_5_wuser_0_reg[i] <= wr_req_desc_5_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_1_reg_we[i])
               wr_req_desc_5_wuser_1_reg[i] <= uc2rb_wr_req_desc_5_wuser_1_reg[i];
             else 
               wr_req_desc_5_wuser_1_reg[i] <= wr_req_desc_5_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_2_reg_we[i])
               wr_req_desc_5_wuser_2_reg[i] <= uc2rb_wr_req_desc_5_wuser_2_reg[i];
             else 
               wr_req_desc_5_wuser_2_reg[i] <= wr_req_desc_5_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_3_reg_we[i])
               wr_req_desc_5_wuser_3_reg[i] <= uc2rb_wr_req_desc_5_wuser_3_reg[i];
             else 
               wr_req_desc_5_wuser_3_reg[i] <= wr_req_desc_5_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_4_reg_we[i])
               wr_req_desc_5_wuser_4_reg[i] <= uc2rb_wr_req_desc_5_wuser_4_reg[i];
             else 
               wr_req_desc_5_wuser_4_reg[i] <= wr_req_desc_5_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_5_reg_we[i])
               wr_req_desc_5_wuser_5_reg[i] <= uc2rb_wr_req_desc_5_wuser_5_reg[i];
             else 
               wr_req_desc_5_wuser_5_reg[i] <= wr_req_desc_5_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_6_reg_we[i])
               wr_req_desc_5_wuser_6_reg[i] <= uc2rb_wr_req_desc_5_wuser_6_reg[i];
             else 
               wr_req_desc_5_wuser_6_reg[i] <= wr_req_desc_5_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_7_reg_we[i])
               wr_req_desc_5_wuser_7_reg[i] <= uc2rb_wr_req_desc_5_wuser_7_reg[i];
             else 
               wr_req_desc_5_wuser_7_reg[i] <= wr_req_desc_5_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_8_reg_we[i])
               wr_req_desc_5_wuser_8_reg[i] <= uc2rb_wr_req_desc_5_wuser_8_reg[i];
             else 
               wr_req_desc_5_wuser_8_reg[i] <= wr_req_desc_5_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_9_reg_we[i])
               wr_req_desc_5_wuser_9_reg[i] <= uc2rb_wr_req_desc_5_wuser_9_reg[i];
             else 
               wr_req_desc_5_wuser_9_reg[i] <= wr_req_desc_5_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_10_reg_we[i])
               wr_req_desc_5_wuser_10_reg[i] <= uc2rb_wr_req_desc_5_wuser_10_reg[i];
             else 
               wr_req_desc_5_wuser_10_reg[i] <= wr_req_desc_5_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_11_reg_we[i])
               wr_req_desc_5_wuser_11_reg[i] <= uc2rb_wr_req_desc_5_wuser_11_reg[i];
             else 
               wr_req_desc_5_wuser_11_reg[i] <= wr_req_desc_5_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_12_reg_we[i])
               wr_req_desc_5_wuser_12_reg[i] <= uc2rb_wr_req_desc_5_wuser_12_reg[i];
             else 
               wr_req_desc_5_wuser_12_reg[i] <= wr_req_desc_5_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_13_reg_we[i])
               wr_req_desc_5_wuser_13_reg[i] <= uc2rb_wr_req_desc_5_wuser_13_reg[i];
             else 
               wr_req_desc_5_wuser_13_reg[i] <= wr_req_desc_5_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_14_reg_we[i])
               wr_req_desc_5_wuser_14_reg[i] <= uc2rb_wr_req_desc_5_wuser_14_reg[i];
             else 
               wr_req_desc_5_wuser_14_reg[i] <= wr_req_desc_5_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_5_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_5_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_5_wuser_15_reg_we[i])
               wr_req_desc_5_wuser_15_reg[i] <= uc2rb_wr_req_desc_5_wuser_15_reg[i];
             else 
               wr_req_desc_5_wuser_15_reg[i] <= wr_req_desc_5_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_5_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_5_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_5_resp_reg_we[i])
               sn_resp_desc_5_resp_reg[i] <= uc2rb_sn_resp_desc_5_resp_reg[i];
             else 
               sn_resp_desc_5_resp_reg[i] <= sn_resp_desc_5_resp_reg[i];
        end
     end
   //RD_REQ_DESC_6_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_txn_type_reg_we[i])
               rd_req_desc_6_txn_type_reg[i] <= uc2rb_rd_req_desc_6_txn_type_reg[i];
             else 
               rd_req_desc_6_txn_type_reg[i] <= rd_req_desc_6_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_6_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_size_reg_we[i])
               rd_req_desc_6_size_reg[i] <= uc2rb_rd_req_desc_6_size_reg[i];
             else 
               rd_req_desc_6_size_reg[i] <= rd_req_desc_6_size_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axsize_reg_we[i])
               rd_req_desc_6_axsize_reg[i] <= uc2rb_rd_req_desc_6_axsize_reg[i];
             else 
               rd_req_desc_6_axsize_reg[i] <= rd_req_desc_6_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_6_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_attr_reg_we[i])
               rd_req_desc_6_attr_reg[i] <= uc2rb_rd_req_desc_6_attr_reg[i];
             else 
               rd_req_desc_6_attr_reg[i] <= rd_req_desc_6_attr_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axaddr_0_reg_we[i])
               rd_req_desc_6_axaddr_0_reg[i] <= uc2rb_rd_req_desc_6_axaddr_0_reg[i];
             else 
               rd_req_desc_6_axaddr_0_reg[i] <= rd_req_desc_6_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axaddr_1_reg_we[i])
               rd_req_desc_6_axaddr_1_reg[i] <= uc2rb_rd_req_desc_6_axaddr_1_reg[i];
             else 
               rd_req_desc_6_axaddr_1_reg[i] <= rd_req_desc_6_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axaddr_2_reg_we[i])
               rd_req_desc_6_axaddr_2_reg[i] <= uc2rb_rd_req_desc_6_axaddr_2_reg[i];
             else 
               rd_req_desc_6_axaddr_2_reg[i] <= rd_req_desc_6_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axaddr_3_reg_we[i])
               rd_req_desc_6_axaddr_3_reg[i] <= uc2rb_rd_req_desc_6_axaddr_3_reg[i];
             else 
               rd_req_desc_6_axaddr_3_reg[i] <= rd_req_desc_6_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axid_0_reg_we[i])
               rd_req_desc_6_axid_0_reg[i] <= uc2rb_rd_req_desc_6_axid_0_reg[i];
             else 
               rd_req_desc_6_axid_0_reg[i] <= rd_req_desc_6_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axid_1_reg_we[i])
               rd_req_desc_6_axid_1_reg[i] <= uc2rb_rd_req_desc_6_axid_1_reg[i];
             else 
               rd_req_desc_6_axid_1_reg[i] <= rd_req_desc_6_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axid_2_reg_we[i])
               rd_req_desc_6_axid_2_reg[i] <= uc2rb_rd_req_desc_6_axid_2_reg[i];
             else 
               rd_req_desc_6_axid_2_reg[i] <= rd_req_desc_6_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axid_3_reg_we[i])
               rd_req_desc_6_axid_3_reg[i] <= uc2rb_rd_req_desc_6_axid_3_reg[i];
             else 
               rd_req_desc_6_axid_3_reg[i] <= rd_req_desc_6_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_0_reg_we[i])
               rd_req_desc_6_axuser_0_reg[i] <= uc2rb_rd_req_desc_6_axuser_0_reg[i];
             else 
               rd_req_desc_6_axuser_0_reg[i] <= rd_req_desc_6_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_1_reg_we[i])
               rd_req_desc_6_axuser_1_reg[i] <= uc2rb_rd_req_desc_6_axuser_1_reg[i];
             else 
               rd_req_desc_6_axuser_1_reg[i] <= rd_req_desc_6_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_2_reg_we[i])
               rd_req_desc_6_axuser_2_reg[i] <= uc2rb_rd_req_desc_6_axuser_2_reg[i];
             else 
               rd_req_desc_6_axuser_2_reg[i] <= rd_req_desc_6_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_3_reg_we[i])
               rd_req_desc_6_axuser_3_reg[i] <= uc2rb_rd_req_desc_6_axuser_3_reg[i];
             else 
               rd_req_desc_6_axuser_3_reg[i] <= rd_req_desc_6_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_4_reg_we[i])
               rd_req_desc_6_axuser_4_reg[i] <= uc2rb_rd_req_desc_6_axuser_4_reg[i];
             else 
               rd_req_desc_6_axuser_4_reg[i] <= rd_req_desc_6_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_5_reg_we[i])
               rd_req_desc_6_axuser_5_reg[i] <= uc2rb_rd_req_desc_6_axuser_5_reg[i];
             else 
               rd_req_desc_6_axuser_5_reg[i] <= rd_req_desc_6_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_6_reg_we[i])
               rd_req_desc_6_axuser_6_reg[i] <= uc2rb_rd_req_desc_6_axuser_6_reg[i];
             else 
               rd_req_desc_6_axuser_6_reg[i] <= rd_req_desc_6_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_7_reg_we[i])
               rd_req_desc_6_axuser_7_reg[i] <= uc2rb_rd_req_desc_6_axuser_7_reg[i];
             else 
               rd_req_desc_6_axuser_7_reg[i] <= rd_req_desc_6_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_8_reg_we[i])
               rd_req_desc_6_axuser_8_reg[i] <= uc2rb_rd_req_desc_6_axuser_8_reg[i];
             else 
               rd_req_desc_6_axuser_8_reg[i] <= rd_req_desc_6_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_9_reg_we[i])
               rd_req_desc_6_axuser_9_reg[i] <= uc2rb_rd_req_desc_6_axuser_9_reg[i];
             else 
               rd_req_desc_6_axuser_9_reg[i] <= rd_req_desc_6_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_10_reg_we[i])
               rd_req_desc_6_axuser_10_reg[i] <= uc2rb_rd_req_desc_6_axuser_10_reg[i];
             else 
               rd_req_desc_6_axuser_10_reg[i] <= rd_req_desc_6_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_11_reg_we[i])
               rd_req_desc_6_axuser_11_reg[i] <= uc2rb_rd_req_desc_6_axuser_11_reg[i];
             else 
               rd_req_desc_6_axuser_11_reg[i] <= rd_req_desc_6_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_12_reg_we[i])
               rd_req_desc_6_axuser_12_reg[i] <= uc2rb_rd_req_desc_6_axuser_12_reg[i];
             else 
               rd_req_desc_6_axuser_12_reg[i] <= rd_req_desc_6_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_13_reg_we[i])
               rd_req_desc_6_axuser_13_reg[i] <= uc2rb_rd_req_desc_6_axuser_13_reg[i];
             else 
               rd_req_desc_6_axuser_13_reg[i] <= rd_req_desc_6_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_14_reg_we[i])
               rd_req_desc_6_axuser_14_reg[i] <= uc2rb_rd_req_desc_6_axuser_14_reg[i];
             else 
               rd_req_desc_6_axuser_14_reg[i] <= rd_req_desc_6_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_6_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_6_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_6_axuser_15_reg_we[i])
               rd_req_desc_6_axuser_15_reg[i] <= uc2rb_rd_req_desc_6_axuser_15_reg[i];
             else 
               rd_req_desc_6_axuser_15_reg[i] <= rd_req_desc_6_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_6_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_txn_type_reg_we[i])
               wr_req_desc_6_txn_type_reg[i] <= uc2rb_wr_req_desc_6_txn_type_reg[i];
             else 
               wr_req_desc_6_txn_type_reg[i] <= wr_req_desc_6_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_6_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_size_reg_we[i])
               wr_req_desc_6_size_reg[i] <= uc2rb_wr_req_desc_6_size_reg[i];
             else 
               wr_req_desc_6_size_reg[i] <= wr_req_desc_6_size_reg[i];
        end
     end
   //WR_REQ_DESC_6_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_data_offset_reg_we[i])
               wr_req_desc_6_data_offset_reg[i] <= uc2rb_wr_req_desc_6_data_offset_reg[i];
             else 
               wr_req_desc_6_data_offset_reg[i] <= wr_req_desc_6_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axsize_reg_we[i])
               wr_req_desc_6_axsize_reg[i] <= uc2rb_wr_req_desc_6_axsize_reg[i];
             else 
               wr_req_desc_6_axsize_reg[i] <= wr_req_desc_6_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_6_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_attr_reg_we[i])
               wr_req_desc_6_attr_reg[i] <= uc2rb_wr_req_desc_6_attr_reg[i];
             else 
               wr_req_desc_6_attr_reg[i] <= wr_req_desc_6_attr_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axaddr_0_reg_we[i])
               wr_req_desc_6_axaddr_0_reg[i] <= uc2rb_wr_req_desc_6_axaddr_0_reg[i];
             else 
               wr_req_desc_6_axaddr_0_reg[i] <= wr_req_desc_6_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axaddr_1_reg_we[i])
               wr_req_desc_6_axaddr_1_reg[i] <= uc2rb_wr_req_desc_6_axaddr_1_reg[i];
             else 
               wr_req_desc_6_axaddr_1_reg[i] <= wr_req_desc_6_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axaddr_2_reg_we[i])
               wr_req_desc_6_axaddr_2_reg[i] <= uc2rb_wr_req_desc_6_axaddr_2_reg[i];
             else 
               wr_req_desc_6_axaddr_2_reg[i] <= wr_req_desc_6_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axaddr_3_reg_we[i])
               wr_req_desc_6_axaddr_3_reg[i] <= uc2rb_wr_req_desc_6_axaddr_3_reg[i];
             else 
               wr_req_desc_6_axaddr_3_reg[i] <= wr_req_desc_6_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axid_0_reg_we[i])
               wr_req_desc_6_axid_0_reg[i] <= uc2rb_wr_req_desc_6_axid_0_reg[i];
             else 
               wr_req_desc_6_axid_0_reg[i] <= wr_req_desc_6_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axid_1_reg_we[i])
               wr_req_desc_6_axid_1_reg[i] <= uc2rb_wr_req_desc_6_axid_1_reg[i];
             else 
               wr_req_desc_6_axid_1_reg[i] <= wr_req_desc_6_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axid_2_reg_we[i])
               wr_req_desc_6_axid_2_reg[i] <= uc2rb_wr_req_desc_6_axid_2_reg[i];
             else 
               wr_req_desc_6_axid_2_reg[i] <= wr_req_desc_6_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axid_3_reg_we[i])
               wr_req_desc_6_axid_3_reg[i] <= uc2rb_wr_req_desc_6_axid_3_reg[i];
             else 
               wr_req_desc_6_axid_3_reg[i] <= wr_req_desc_6_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_0_reg_we[i])
               wr_req_desc_6_axuser_0_reg[i] <= uc2rb_wr_req_desc_6_axuser_0_reg[i];
             else 
               wr_req_desc_6_axuser_0_reg[i] <= wr_req_desc_6_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_1_reg_we[i])
               wr_req_desc_6_axuser_1_reg[i] <= uc2rb_wr_req_desc_6_axuser_1_reg[i];
             else 
               wr_req_desc_6_axuser_1_reg[i] <= wr_req_desc_6_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_2_reg_we[i])
               wr_req_desc_6_axuser_2_reg[i] <= uc2rb_wr_req_desc_6_axuser_2_reg[i];
             else 
               wr_req_desc_6_axuser_2_reg[i] <= wr_req_desc_6_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_3_reg_we[i])
               wr_req_desc_6_axuser_3_reg[i] <= uc2rb_wr_req_desc_6_axuser_3_reg[i];
             else 
               wr_req_desc_6_axuser_3_reg[i] <= wr_req_desc_6_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_4_reg_we[i])
               wr_req_desc_6_axuser_4_reg[i] <= uc2rb_wr_req_desc_6_axuser_4_reg[i];
             else 
               wr_req_desc_6_axuser_4_reg[i] <= wr_req_desc_6_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_5_reg_we[i])
               wr_req_desc_6_axuser_5_reg[i] <= uc2rb_wr_req_desc_6_axuser_5_reg[i];
             else 
               wr_req_desc_6_axuser_5_reg[i] <= wr_req_desc_6_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_6_reg_we[i])
               wr_req_desc_6_axuser_6_reg[i] <= uc2rb_wr_req_desc_6_axuser_6_reg[i];
             else 
               wr_req_desc_6_axuser_6_reg[i] <= wr_req_desc_6_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_7_reg_we[i])
               wr_req_desc_6_axuser_7_reg[i] <= uc2rb_wr_req_desc_6_axuser_7_reg[i];
             else 
               wr_req_desc_6_axuser_7_reg[i] <= wr_req_desc_6_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_8_reg_we[i])
               wr_req_desc_6_axuser_8_reg[i] <= uc2rb_wr_req_desc_6_axuser_8_reg[i];
             else 
               wr_req_desc_6_axuser_8_reg[i] <= wr_req_desc_6_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_9_reg_we[i])
               wr_req_desc_6_axuser_9_reg[i] <= uc2rb_wr_req_desc_6_axuser_9_reg[i];
             else 
               wr_req_desc_6_axuser_9_reg[i] <= wr_req_desc_6_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_10_reg_we[i])
               wr_req_desc_6_axuser_10_reg[i] <= uc2rb_wr_req_desc_6_axuser_10_reg[i];
             else 
               wr_req_desc_6_axuser_10_reg[i] <= wr_req_desc_6_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_11_reg_we[i])
               wr_req_desc_6_axuser_11_reg[i] <= uc2rb_wr_req_desc_6_axuser_11_reg[i];
             else 
               wr_req_desc_6_axuser_11_reg[i] <= wr_req_desc_6_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_12_reg_we[i])
               wr_req_desc_6_axuser_12_reg[i] <= uc2rb_wr_req_desc_6_axuser_12_reg[i];
             else 
               wr_req_desc_6_axuser_12_reg[i] <= wr_req_desc_6_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_13_reg_we[i])
               wr_req_desc_6_axuser_13_reg[i] <= uc2rb_wr_req_desc_6_axuser_13_reg[i];
             else 
               wr_req_desc_6_axuser_13_reg[i] <= wr_req_desc_6_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_14_reg_we[i])
               wr_req_desc_6_axuser_14_reg[i] <= uc2rb_wr_req_desc_6_axuser_14_reg[i];
             else 
               wr_req_desc_6_axuser_14_reg[i] <= wr_req_desc_6_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_6_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_axuser_15_reg_we[i])
               wr_req_desc_6_axuser_15_reg[i] <= uc2rb_wr_req_desc_6_axuser_15_reg[i];
             else 
               wr_req_desc_6_axuser_15_reg[i] <= wr_req_desc_6_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_0_reg_we[i])
               wr_req_desc_6_wuser_0_reg[i] <= uc2rb_wr_req_desc_6_wuser_0_reg[i];
             else 
               wr_req_desc_6_wuser_0_reg[i] <= wr_req_desc_6_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_1_reg_we[i])
               wr_req_desc_6_wuser_1_reg[i] <= uc2rb_wr_req_desc_6_wuser_1_reg[i];
             else 
               wr_req_desc_6_wuser_1_reg[i] <= wr_req_desc_6_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_2_reg_we[i])
               wr_req_desc_6_wuser_2_reg[i] <= uc2rb_wr_req_desc_6_wuser_2_reg[i];
             else 
               wr_req_desc_6_wuser_2_reg[i] <= wr_req_desc_6_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_3_reg_we[i])
               wr_req_desc_6_wuser_3_reg[i] <= uc2rb_wr_req_desc_6_wuser_3_reg[i];
             else 
               wr_req_desc_6_wuser_3_reg[i] <= wr_req_desc_6_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_4_reg_we[i])
               wr_req_desc_6_wuser_4_reg[i] <= uc2rb_wr_req_desc_6_wuser_4_reg[i];
             else 
               wr_req_desc_6_wuser_4_reg[i] <= wr_req_desc_6_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_5_reg_we[i])
               wr_req_desc_6_wuser_5_reg[i] <= uc2rb_wr_req_desc_6_wuser_5_reg[i];
             else 
               wr_req_desc_6_wuser_5_reg[i] <= wr_req_desc_6_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_6_reg_we[i])
               wr_req_desc_6_wuser_6_reg[i] <= uc2rb_wr_req_desc_6_wuser_6_reg[i];
             else 
               wr_req_desc_6_wuser_6_reg[i] <= wr_req_desc_6_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_7_reg_we[i])
               wr_req_desc_6_wuser_7_reg[i] <= uc2rb_wr_req_desc_6_wuser_7_reg[i];
             else 
               wr_req_desc_6_wuser_7_reg[i] <= wr_req_desc_6_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_8_reg_we[i])
               wr_req_desc_6_wuser_8_reg[i] <= uc2rb_wr_req_desc_6_wuser_8_reg[i];
             else 
               wr_req_desc_6_wuser_8_reg[i] <= wr_req_desc_6_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_9_reg_we[i])
               wr_req_desc_6_wuser_9_reg[i] <= uc2rb_wr_req_desc_6_wuser_9_reg[i];
             else 
               wr_req_desc_6_wuser_9_reg[i] <= wr_req_desc_6_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_10_reg_we[i])
               wr_req_desc_6_wuser_10_reg[i] <= uc2rb_wr_req_desc_6_wuser_10_reg[i];
             else 
               wr_req_desc_6_wuser_10_reg[i] <= wr_req_desc_6_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_11_reg_we[i])
               wr_req_desc_6_wuser_11_reg[i] <= uc2rb_wr_req_desc_6_wuser_11_reg[i];
             else 
               wr_req_desc_6_wuser_11_reg[i] <= wr_req_desc_6_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_12_reg_we[i])
               wr_req_desc_6_wuser_12_reg[i] <= uc2rb_wr_req_desc_6_wuser_12_reg[i];
             else 
               wr_req_desc_6_wuser_12_reg[i] <= wr_req_desc_6_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_13_reg_we[i])
               wr_req_desc_6_wuser_13_reg[i] <= uc2rb_wr_req_desc_6_wuser_13_reg[i];
             else 
               wr_req_desc_6_wuser_13_reg[i] <= wr_req_desc_6_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_14_reg_we[i])
               wr_req_desc_6_wuser_14_reg[i] <= uc2rb_wr_req_desc_6_wuser_14_reg[i];
             else 
               wr_req_desc_6_wuser_14_reg[i] <= wr_req_desc_6_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_6_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_6_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_6_wuser_15_reg_we[i])
               wr_req_desc_6_wuser_15_reg[i] <= uc2rb_wr_req_desc_6_wuser_15_reg[i];
             else 
               wr_req_desc_6_wuser_15_reg[i] <= wr_req_desc_6_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_6_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_6_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_6_resp_reg_we[i])
               sn_resp_desc_6_resp_reg[i] <= uc2rb_sn_resp_desc_6_resp_reg[i];
             else 
               sn_resp_desc_6_resp_reg[i] <= sn_resp_desc_6_resp_reg[i];
        end
     end
   //RD_REQ_DESC_7_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_txn_type_reg_we[i])
               rd_req_desc_7_txn_type_reg[i] <= uc2rb_rd_req_desc_7_txn_type_reg[i];
             else 
               rd_req_desc_7_txn_type_reg[i] <= rd_req_desc_7_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_7_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_size_reg_we[i])
               rd_req_desc_7_size_reg[i] <= uc2rb_rd_req_desc_7_size_reg[i];
             else 
               rd_req_desc_7_size_reg[i] <= rd_req_desc_7_size_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axsize_reg_we[i])
               rd_req_desc_7_axsize_reg[i] <= uc2rb_rd_req_desc_7_axsize_reg[i];
             else 
               rd_req_desc_7_axsize_reg[i] <= rd_req_desc_7_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_7_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_attr_reg_we[i])
               rd_req_desc_7_attr_reg[i] <= uc2rb_rd_req_desc_7_attr_reg[i];
             else 
               rd_req_desc_7_attr_reg[i] <= rd_req_desc_7_attr_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axaddr_0_reg_we[i])
               rd_req_desc_7_axaddr_0_reg[i] <= uc2rb_rd_req_desc_7_axaddr_0_reg[i];
             else 
               rd_req_desc_7_axaddr_0_reg[i] <= rd_req_desc_7_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axaddr_1_reg_we[i])
               rd_req_desc_7_axaddr_1_reg[i] <= uc2rb_rd_req_desc_7_axaddr_1_reg[i];
             else 
               rd_req_desc_7_axaddr_1_reg[i] <= rd_req_desc_7_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axaddr_2_reg_we[i])
               rd_req_desc_7_axaddr_2_reg[i] <= uc2rb_rd_req_desc_7_axaddr_2_reg[i];
             else 
               rd_req_desc_7_axaddr_2_reg[i] <= rd_req_desc_7_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axaddr_3_reg_we[i])
               rd_req_desc_7_axaddr_3_reg[i] <= uc2rb_rd_req_desc_7_axaddr_3_reg[i];
             else 
               rd_req_desc_7_axaddr_3_reg[i] <= rd_req_desc_7_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axid_0_reg_we[i])
               rd_req_desc_7_axid_0_reg[i] <= uc2rb_rd_req_desc_7_axid_0_reg[i];
             else 
               rd_req_desc_7_axid_0_reg[i] <= rd_req_desc_7_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axid_1_reg_we[i])
               rd_req_desc_7_axid_1_reg[i] <= uc2rb_rd_req_desc_7_axid_1_reg[i];
             else 
               rd_req_desc_7_axid_1_reg[i] <= rd_req_desc_7_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axid_2_reg_we[i])
               rd_req_desc_7_axid_2_reg[i] <= uc2rb_rd_req_desc_7_axid_2_reg[i];
             else 
               rd_req_desc_7_axid_2_reg[i] <= rd_req_desc_7_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axid_3_reg_we[i])
               rd_req_desc_7_axid_3_reg[i] <= uc2rb_rd_req_desc_7_axid_3_reg[i];
             else 
               rd_req_desc_7_axid_3_reg[i] <= rd_req_desc_7_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_0_reg_we[i])
               rd_req_desc_7_axuser_0_reg[i] <= uc2rb_rd_req_desc_7_axuser_0_reg[i];
             else 
               rd_req_desc_7_axuser_0_reg[i] <= rd_req_desc_7_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_1_reg_we[i])
               rd_req_desc_7_axuser_1_reg[i] <= uc2rb_rd_req_desc_7_axuser_1_reg[i];
             else 
               rd_req_desc_7_axuser_1_reg[i] <= rd_req_desc_7_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_2_reg_we[i])
               rd_req_desc_7_axuser_2_reg[i] <= uc2rb_rd_req_desc_7_axuser_2_reg[i];
             else 
               rd_req_desc_7_axuser_2_reg[i] <= rd_req_desc_7_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_3_reg_we[i])
               rd_req_desc_7_axuser_3_reg[i] <= uc2rb_rd_req_desc_7_axuser_3_reg[i];
             else 
               rd_req_desc_7_axuser_3_reg[i] <= rd_req_desc_7_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_4_reg_we[i])
               rd_req_desc_7_axuser_4_reg[i] <= uc2rb_rd_req_desc_7_axuser_4_reg[i];
             else 
               rd_req_desc_7_axuser_4_reg[i] <= rd_req_desc_7_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_5_reg_we[i])
               rd_req_desc_7_axuser_5_reg[i] <= uc2rb_rd_req_desc_7_axuser_5_reg[i];
             else 
               rd_req_desc_7_axuser_5_reg[i] <= rd_req_desc_7_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_6_reg_we[i])
               rd_req_desc_7_axuser_6_reg[i] <= uc2rb_rd_req_desc_7_axuser_6_reg[i];
             else 
               rd_req_desc_7_axuser_6_reg[i] <= rd_req_desc_7_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_7_reg_we[i])
               rd_req_desc_7_axuser_7_reg[i] <= uc2rb_rd_req_desc_7_axuser_7_reg[i];
             else 
               rd_req_desc_7_axuser_7_reg[i] <= rd_req_desc_7_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_8_reg_we[i])
               rd_req_desc_7_axuser_8_reg[i] <= uc2rb_rd_req_desc_7_axuser_8_reg[i];
             else 
               rd_req_desc_7_axuser_8_reg[i] <= rd_req_desc_7_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_9_reg_we[i])
               rd_req_desc_7_axuser_9_reg[i] <= uc2rb_rd_req_desc_7_axuser_9_reg[i];
             else 
               rd_req_desc_7_axuser_9_reg[i] <= rd_req_desc_7_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_10_reg_we[i])
               rd_req_desc_7_axuser_10_reg[i] <= uc2rb_rd_req_desc_7_axuser_10_reg[i];
             else 
               rd_req_desc_7_axuser_10_reg[i] <= rd_req_desc_7_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_11_reg_we[i])
               rd_req_desc_7_axuser_11_reg[i] <= uc2rb_rd_req_desc_7_axuser_11_reg[i];
             else 
               rd_req_desc_7_axuser_11_reg[i] <= rd_req_desc_7_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_12_reg_we[i])
               rd_req_desc_7_axuser_12_reg[i] <= uc2rb_rd_req_desc_7_axuser_12_reg[i];
             else 
               rd_req_desc_7_axuser_12_reg[i] <= rd_req_desc_7_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_13_reg_we[i])
               rd_req_desc_7_axuser_13_reg[i] <= uc2rb_rd_req_desc_7_axuser_13_reg[i];
             else 
               rd_req_desc_7_axuser_13_reg[i] <= rd_req_desc_7_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_14_reg_we[i])
               rd_req_desc_7_axuser_14_reg[i] <= uc2rb_rd_req_desc_7_axuser_14_reg[i];
             else 
               rd_req_desc_7_axuser_14_reg[i] <= rd_req_desc_7_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_7_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_7_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_7_axuser_15_reg_we[i])
               rd_req_desc_7_axuser_15_reg[i] <= uc2rb_rd_req_desc_7_axuser_15_reg[i];
             else 
               rd_req_desc_7_axuser_15_reg[i] <= rd_req_desc_7_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_7_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_txn_type_reg_we[i])
               wr_req_desc_7_txn_type_reg[i] <= uc2rb_wr_req_desc_7_txn_type_reg[i];
             else 
               wr_req_desc_7_txn_type_reg[i] <= wr_req_desc_7_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_7_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_size_reg_we[i])
               wr_req_desc_7_size_reg[i] <= uc2rb_wr_req_desc_7_size_reg[i];
             else 
               wr_req_desc_7_size_reg[i] <= wr_req_desc_7_size_reg[i];
        end
     end
   //WR_REQ_DESC_7_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_data_offset_reg_we[i])
               wr_req_desc_7_data_offset_reg[i] <= uc2rb_wr_req_desc_7_data_offset_reg[i];
             else 
               wr_req_desc_7_data_offset_reg[i] <= wr_req_desc_7_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axsize_reg_we[i])
               wr_req_desc_7_axsize_reg[i] <= uc2rb_wr_req_desc_7_axsize_reg[i];
             else 
               wr_req_desc_7_axsize_reg[i] <= wr_req_desc_7_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_7_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_attr_reg_we[i])
               wr_req_desc_7_attr_reg[i] <= uc2rb_wr_req_desc_7_attr_reg[i];
             else 
               wr_req_desc_7_attr_reg[i] <= wr_req_desc_7_attr_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axaddr_0_reg_we[i])
               wr_req_desc_7_axaddr_0_reg[i] <= uc2rb_wr_req_desc_7_axaddr_0_reg[i];
             else 
               wr_req_desc_7_axaddr_0_reg[i] <= wr_req_desc_7_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axaddr_1_reg_we[i])
               wr_req_desc_7_axaddr_1_reg[i] <= uc2rb_wr_req_desc_7_axaddr_1_reg[i];
             else 
               wr_req_desc_7_axaddr_1_reg[i] <= wr_req_desc_7_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axaddr_2_reg_we[i])
               wr_req_desc_7_axaddr_2_reg[i] <= uc2rb_wr_req_desc_7_axaddr_2_reg[i];
             else 
               wr_req_desc_7_axaddr_2_reg[i] <= wr_req_desc_7_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axaddr_3_reg_we[i])
               wr_req_desc_7_axaddr_3_reg[i] <= uc2rb_wr_req_desc_7_axaddr_3_reg[i];
             else 
               wr_req_desc_7_axaddr_3_reg[i] <= wr_req_desc_7_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axid_0_reg_we[i])
               wr_req_desc_7_axid_0_reg[i] <= uc2rb_wr_req_desc_7_axid_0_reg[i];
             else 
               wr_req_desc_7_axid_0_reg[i] <= wr_req_desc_7_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axid_1_reg_we[i])
               wr_req_desc_7_axid_1_reg[i] <= uc2rb_wr_req_desc_7_axid_1_reg[i];
             else 
               wr_req_desc_7_axid_1_reg[i] <= wr_req_desc_7_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axid_2_reg_we[i])
               wr_req_desc_7_axid_2_reg[i] <= uc2rb_wr_req_desc_7_axid_2_reg[i];
             else 
               wr_req_desc_7_axid_2_reg[i] <= wr_req_desc_7_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axid_3_reg_we[i])
               wr_req_desc_7_axid_3_reg[i] <= uc2rb_wr_req_desc_7_axid_3_reg[i];
             else 
               wr_req_desc_7_axid_3_reg[i] <= wr_req_desc_7_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_0_reg_we[i])
               wr_req_desc_7_axuser_0_reg[i] <= uc2rb_wr_req_desc_7_axuser_0_reg[i];
             else 
               wr_req_desc_7_axuser_0_reg[i] <= wr_req_desc_7_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_1_reg_we[i])
               wr_req_desc_7_axuser_1_reg[i] <= uc2rb_wr_req_desc_7_axuser_1_reg[i];
             else 
               wr_req_desc_7_axuser_1_reg[i] <= wr_req_desc_7_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_2_reg_we[i])
               wr_req_desc_7_axuser_2_reg[i] <= uc2rb_wr_req_desc_7_axuser_2_reg[i];
             else 
               wr_req_desc_7_axuser_2_reg[i] <= wr_req_desc_7_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_3_reg_we[i])
               wr_req_desc_7_axuser_3_reg[i] <= uc2rb_wr_req_desc_7_axuser_3_reg[i];
             else 
               wr_req_desc_7_axuser_3_reg[i] <= wr_req_desc_7_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_4_reg_we[i])
               wr_req_desc_7_axuser_4_reg[i] <= uc2rb_wr_req_desc_7_axuser_4_reg[i];
             else 
               wr_req_desc_7_axuser_4_reg[i] <= wr_req_desc_7_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_5_reg_we[i])
               wr_req_desc_7_axuser_5_reg[i] <= uc2rb_wr_req_desc_7_axuser_5_reg[i];
             else 
               wr_req_desc_7_axuser_5_reg[i] <= wr_req_desc_7_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_6_reg_we[i])
               wr_req_desc_7_axuser_6_reg[i] <= uc2rb_wr_req_desc_7_axuser_6_reg[i];
             else 
               wr_req_desc_7_axuser_6_reg[i] <= wr_req_desc_7_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_7_reg_we[i])
               wr_req_desc_7_axuser_7_reg[i] <= uc2rb_wr_req_desc_7_axuser_7_reg[i];
             else 
               wr_req_desc_7_axuser_7_reg[i] <= wr_req_desc_7_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_8_reg_we[i])
               wr_req_desc_7_axuser_8_reg[i] <= uc2rb_wr_req_desc_7_axuser_8_reg[i];
             else 
               wr_req_desc_7_axuser_8_reg[i] <= wr_req_desc_7_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_9_reg_we[i])
               wr_req_desc_7_axuser_9_reg[i] <= uc2rb_wr_req_desc_7_axuser_9_reg[i];
             else 
               wr_req_desc_7_axuser_9_reg[i] <= wr_req_desc_7_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_10_reg_we[i])
               wr_req_desc_7_axuser_10_reg[i] <= uc2rb_wr_req_desc_7_axuser_10_reg[i];
             else 
               wr_req_desc_7_axuser_10_reg[i] <= wr_req_desc_7_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_11_reg_we[i])
               wr_req_desc_7_axuser_11_reg[i] <= uc2rb_wr_req_desc_7_axuser_11_reg[i];
             else 
               wr_req_desc_7_axuser_11_reg[i] <= wr_req_desc_7_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_12_reg_we[i])
               wr_req_desc_7_axuser_12_reg[i] <= uc2rb_wr_req_desc_7_axuser_12_reg[i];
             else 
               wr_req_desc_7_axuser_12_reg[i] <= wr_req_desc_7_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_13_reg_we[i])
               wr_req_desc_7_axuser_13_reg[i] <= uc2rb_wr_req_desc_7_axuser_13_reg[i];
             else 
               wr_req_desc_7_axuser_13_reg[i] <= wr_req_desc_7_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_14_reg_we[i])
               wr_req_desc_7_axuser_14_reg[i] <= uc2rb_wr_req_desc_7_axuser_14_reg[i];
             else 
               wr_req_desc_7_axuser_14_reg[i] <= wr_req_desc_7_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_7_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_axuser_15_reg_we[i])
               wr_req_desc_7_axuser_15_reg[i] <= uc2rb_wr_req_desc_7_axuser_15_reg[i];
             else 
               wr_req_desc_7_axuser_15_reg[i] <= wr_req_desc_7_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_0_reg_we[i])
               wr_req_desc_7_wuser_0_reg[i] <= uc2rb_wr_req_desc_7_wuser_0_reg[i];
             else 
               wr_req_desc_7_wuser_0_reg[i] <= wr_req_desc_7_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_1_reg_we[i])
               wr_req_desc_7_wuser_1_reg[i] <= uc2rb_wr_req_desc_7_wuser_1_reg[i];
             else 
               wr_req_desc_7_wuser_1_reg[i] <= wr_req_desc_7_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_2_reg_we[i])
               wr_req_desc_7_wuser_2_reg[i] <= uc2rb_wr_req_desc_7_wuser_2_reg[i];
             else 
               wr_req_desc_7_wuser_2_reg[i] <= wr_req_desc_7_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_3_reg_we[i])
               wr_req_desc_7_wuser_3_reg[i] <= uc2rb_wr_req_desc_7_wuser_3_reg[i];
             else 
               wr_req_desc_7_wuser_3_reg[i] <= wr_req_desc_7_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_4_reg_we[i])
               wr_req_desc_7_wuser_4_reg[i] <= uc2rb_wr_req_desc_7_wuser_4_reg[i];
             else 
               wr_req_desc_7_wuser_4_reg[i] <= wr_req_desc_7_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_5_reg_we[i])
               wr_req_desc_7_wuser_5_reg[i] <= uc2rb_wr_req_desc_7_wuser_5_reg[i];
             else 
               wr_req_desc_7_wuser_5_reg[i] <= wr_req_desc_7_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_6_reg_we[i])
               wr_req_desc_7_wuser_6_reg[i] <= uc2rb_wr_req_desc_7_wuser_6_reg[i];
             else 
               wr_req_desc_7_wuser_6_reg[i] <= wr_req_desc_7_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_7_reg_we[i])
               wr_req_desc_7_wuser_7_reg[i] <= uc2rb_wr_req_desc_7_wuser_7_reg[i];
             else 
               wr_req_desc_7_wuser_7_reg[i] <= wr_req_desc_7_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_8_reg_we[i])
               wr_req_desc_7_wuser_8_reg[i] <= uc2rb_wr_req_desc_7_wuser_8_reg[i];
             else 
               wr_req_desc_7_wuser_8_reg[i] <= wr_req_desc_7_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_9_reg_we[i])
               wr_req_desc_7_wuser_9_reg[i] <= uc2rb_wr_req_desc_7_wuser_9_reg[i];
             else 
               wr_req_desc_7_wuser_9_reg[i] <= wr_req_desc_7_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_10_reg_we[i])
               wr_req_desc_7_wuser_10_reg[i] <= uc2rb_wr_req_desc_7_wuser_10_reg[i];
             else 
               wr_req_desc_7_wuser_10_reg[i] <= wr_req_desc_7_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_11_reg_we[i])
               wr_req_desc_7_wuser_11_reg[i] <= uc2rb_wr_req_desc_7_wuser_11_reg[i];
             else 
               wr_req_desc_7_wuser_11_reg[i] <= wr_req_desc_7_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_12_reg_we[i])
               wr_req_desc_7_wuser_12_reg[i] <= uc2rb_wr_req_desc_7_wuser_12_reg[i];
             else 
               wr_req_desc_7_wuser_12_reg[i] <= wr_req_desc_7_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_13_reg_we[i])
               wr_req_desc_7_wuser_13_reg[i] <= uc2rb_wr_req_desc_7_wuser_13_reg[i];
             else 
               wr_req_desc_7_wuser_13_reg[i] <= wr_req_desc_7_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_14_reg_we[i])
               wr_req_desc_7_wuser_14_reg[i] <= uc2rb_wr_req_desc_7_wuser_14_reg[i];
             else 
               wr_req_desc_7_wuser_14_reg[i] <= wr_req_desc_7_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_7_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_7_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_7_wuser_15_reg_we[i])
               wr_req_desc_7_wuser_15_reg[i] <= uc2rb_wr_req_desc_7_wuser_15_reg[i];
             else 
               wr_req_desc_7_wuser_15_reg[i] <= wr_req_desc_7_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_7_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_7_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_7_resp_reg_we[i])
               sn_resp_desc_7_resp_reg[i] <= uc2rb_sn_resp_desc_7_resp_reg[i];
             else 
               sn_resp_desc_7_resp_reg[i] <= sn_resp_desc_7_resp_reg[i];
        end
     end
   //RD_REQ_DESC_8_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_txn_type_reg_we[i])
               rd_req_desc_8_txn_type_reg[i] <= uc2rb_rd_req_desc_8_txn_type_reg[i];
             else 
               rd_req_desc_8_txn_type_reg[i] <= rd_req_desc_8_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_8_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_size_reg_we[i])
               rd_req_desc_8_size_reg[i] <= uc2rb_rd_req_desc_8_size_reg[i];
             else 
               rd_req_desc_8_size_reg[i] <= rd_req_desc_8_size_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axsize_reg_we[i])
               rd_req_desc_8_axsize_reg[i] <= uc2rb_rd_req_desc_8_axsize_reg[i];
             else 
               rd_req_desc_8_axsize_reg[i] <= rd_req_desc_8_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_8_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_attr_reg_we[i])
               rd_req_desc_8_attr_reg[i] <= uc2rb_rd_req_desc_8_attr_reg[i];
             else 
               rd_req_desc_8_attr_reg[i] <= rd_req_desc_8_attr_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axaddr_0_reg_we[i])
               rd_req_desc_8_axaddr_0_reg[i] <= uc2rb_rd_req_desc_8_axaddr_0_reg[i];
             else 
               rd_req_desc_8_axaddr_0_reg[i] <= rd_req_desc_8_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axaddr_1_reg_we[i])
               rd_req_desc_8_axaddr_1_reg[i] <= uc2rb_rd_req_desc_8_axaddr_1_reg[i];
             else 
               rd_req_desc_8_axaddr_1_reg[i] <= rd_req_desc_8_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axaddr_2_reg_we[i])
               rd_req_desc_8_axaddr_2_reg[i] <= uc2rb_rd_req_desc_8_axaddr_2_reg[i];
             else 
               rd_req_desc_8_axaddr_2_reg[i] <= rd_req_desc_8_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axaddr_3_reg_we[i])
               rd_req_desc_8_axaddr_3_reg[i] <= uc2rb_rd_req_desc_8_axaddr_3_reg[i];
             else 
               rd_req_desc_8_axaddr_3_reg[i] <= rd_req_desc_8_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axid_0_reg_we[i])
               rd_req_desc_8_axid_0_reg[i] <= uc2rb_rd_req_desc_8_axid_0_reg[i];
             else 
               rd_req_desc_8_axid_0_reg[i] <= rd_req_desc_8_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axid_1_reg_we[i])
               rd_req_desc_8_axid_1_reg[i] <= uc2rb_rd_req_desc_8_axid_1_reg[i];
             else 
               rd_req_desc_8_axid_1_reg[i] <= rd_req_desc_8_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axid_2_reg_we[i])
               rd_req_desc_8_axid_2_reg[i] <= uc2rb_rd_req_desc_8_axid_2_reg[i];
             else 
               rd_req_desc_8_axid_2_reg[i] <= rd_req_desc_8_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axid_3_reg_we[i])
               rd_req_desc_8_axid_3_reg[i] <= uc2rb_rd_req_desc_8_axid_3_reg[i];
             else 
               rd_req_desc_8_axid_3_reg[i] <= rd_req_desc_8_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_0_reg_we[i])
               rd_req_desc_8_axuser_0_reg[i] <= uc2rb_rd_req_desc_8_axuser_0_reg[i];
             else 
               rd_req_desc_8_axuser_0_reg[i] <= rd_req_desc_8_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_1_reg_we[i])
               rd_req_desc_8_axuser_1_reg[i] <= uc2rb_rd_req_desc_8_axuser_1_reg[i];
             else 
               rd_req_desc_8_axuser_1_reg[i] <= rd_req_desc_8_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_2_reg_we[i])
               rd_req_desc_8_axuser_2_reg[i] <= uc2rb_rd_req_desc_8_axuser_2_reg[i];
             else 
               rd_req_desc_8_axuser_2_reg[i] <= rd_req_desc_8_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_3_reg_we[i])
               rd_req_desc_8_axuser_3_reg[i] <= uc2rb_rd_req_desc_8_axuser_3_reg[i];
             else 
               rd_req_desc_8_axuser_3_reg[i] <= rd_req_desc_8_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_4_reg_we[i])
               rd_req_desc_8_axuser_4_reg[i] <= uc2rb_rd_req_desc_8_axuser_4_reg[i];
             else 
               rd_req_desc_8_axuser_4_reg[i] <= rd_req_desc_8_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_5_reg_we[i])
               rd_req_desc_8_axuser_5_reg[i] <= uc2rb_rd_req_desc_8_axuser_5_reg[i];
             else 
               rd_req_desc_8_axuser_5_reg[i] <= rd_req_desc_8_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_6_reg_we[i])
               rd_req_desc_8_axuser_6_reg[i] <= uc2rb_rd_req_desc_8_axuser_6_reg[i];
             else 
               rd_req_desc_8_axuser_6_reg[i] <= rd_req_desc_8_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_7_reg_we[i])
               rd_req_desc_8_axuser_7_reg[i] <= uc2rb_rd_req_desc_8_axuser_7_reg[i];
             else 
               rd_req_desc_8_axuser_7_reg[i] <= rd_req_desc_8_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_8_reg_we[i])
               rd_req_desc_8_axuser_8_reg[i] <= uc2rb_rd_req_desc_8_axuser_8_reg[i];
             else 
               rd_req_desc_8_axuser_8_reg[i] <= rd_req_desc_8_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_9_reg_we[i])
               rd_req_desc_8_axuser_9_reg[i] <= uc2rb_rd_req_desc_8_axuser_9_reg[i];
             else 
               rd_req_desc_8_axuser_9_reg[i] <= rd_req_desc_8_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_10_reg_we[i])
               rd_req_desc_8_axuser_10_reg[i] <= uc2rb_rd_req_desc_8_axuser_10_reg[i];
             else 
               rd_req_desc_8_axuser_10_reg[i] <= rd_req_desc_8_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_11_reg_we[i])
               rd_req_desc_8_axuser_11_reg[i] <= uc2rb_rd_req_desc_8_axuser_11_reg[i];
             else 
               rd_req_desc_8_axuser_11_reg[i] <= rd_req_desc_8_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_12_reg_we[i])
               rd_req_desc_8_axuser_12_reg[i] <= uc2rb_rd_req_desc_8_axuser_12_reg[i];
             else 
               rd_req_desc_8_axuser_12_reg[i] <= rd_req_desc_8_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_13_reg_we[i])
               rd_req_desc_8_axuser_13_reg[i] <= uc2rb_rd_req_desc_8_axuser_13_reg[i];
             else 
               rd_req_desc_8_axuser_13_reg[i] <= rd_req_desc_8_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_14_reg_we[i])
               rd_req_desc_8_axuser_14_reg[i] <= uc2rb_rd_req_desc_8_axuser_14_reg[i];
             else 
               rd_req_desc_8_axuser_14_reg[i] <= rd_req_desc_8_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_8_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_8_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_8_axuser_15_reg_we[i])
               rd_req_desc_8_axuser_15_reg[i] <= uc2rb_rd_req_desc_8_axuser_15_reg[i];
             else 
               rd_req_desc_8_axuser_15_reg[i] <= rd_req_desc_8_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_8_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_txn_type_reg_we[i])
               wr_req_desc_8_txn_type_reg[i] <= uc2rb_wr_req_desc_8_txn_type_reg[i];
             else 
               wr_req_desc_8_txn_type_reg[i] <= wr_req_desc_8_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_8_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_size_reg_we[i])
               wr_req_desc_8_size_reg[i] <= uc2rb_wr_req_desc_8_size_reg[i];
             else 
               wr_req_desc_8_size_reg[i] <= wr_req_desc_8_size_reg[i];
        end
     end
   //WR_REQ_DESC_8_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_data_offset_reg_we[i])
               wr_req_desc_8_data_offset_reg[i] <= uc2rb_wr_req_desc_8_data_offset_reg[i];
             else 
               wr_req_desc_8_data_offset_reg[i] <= wr_req_desc_8_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axsize_reg_we[i])
               wr_req_desc_8_axsize_reg[i] <= uc2rb_wr_req_desc_8_axsize_reg[i];
             else 
               wr_req_desc_8_axsize_reg[i] <= wr_req_desc_8_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_8_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_attr_reg_we[i])
               wr_req_desc_8_attr_reg[i] <= uc2rb_wr_req_desc_8_attr_reg[i];
             else 
               wr_req_desc_8_attr_reg[i] <= wr_req_desc_8_attr_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axaddr_0_reg_we[i])
               wr_req_desc_8_axaddr_0_reg[i] <= uc2rb_wr_req_desc_8_axaddr_0_reg[i];
             else 
               wr_req_desc_8_axaddr_0_reg[i] <= wr_req_desc_8_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axaddr_1_reg_we[i])
               wr_req_desc_8_axaddr_1_reg[i] <= uc2rb_wr_req_desc_8_axaddr_1_reg[i];
             else 
               wr_req_desc_8_axaddr_1_reg[i] <= wr_req_desc_8_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axaddr_2_reg_we[i])
               wr_req_desc_8_axaddr_2_reg[i] <= uc2rb_wr_req_desc_8_axaddr_2_reg[i];
             else 
               wr_req_desc_8_axaddr_2_reg[i] <= wr_req_desc_8_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axaddr_3_reg_we[i])
               wr_req_desc_8_axaddr_3_reg[i] <= uc2rb_wr_req_desc_8_axaddr_3_reg[i];
             else 
               wr_req_desc_8_axaddr_3_reg[i] <= wr_req_desc_8_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axid_0_reg_we[i])
               wr_req_desc_8_axid_0_reg[i] <= uc2rb_wr_req_desc_8_axid_0_reg[i];
             else 
               wr_req_desc_8_axid_0_reg[i] <= wr_req_desc_8_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axid_1_reg_we[i])
               wr_req_desc_8_axid_1_reg[i] <= uc2rb_wr_req_desc_8_axid_1_reg[i];
             else 
               wr_req_desc_8_axid_1_reg[i] <= wr_req_desc_8_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axid_2_reg_we[i])
               wr_req_desc_8_axid_2_reg[i] <= uc2rb_wr_req_desc_8_axid_2_reg[i];
             else 
               wr_req_desc_8_axid_2_reg[i] <= wr_req_desc_8_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axid_3_reg_we[i])
               wr_req_desc_8_axid_3_reg[i] <= uc2rb_wr_req_desc_8_axid_3_reg[i];
             else 
               wr_req_desc_8_axid_3_reg[i] <= wr_req_desc_8_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_0_reg_we[i])
               wr_req_desc_8_axuser_0_reg[i] <= uc2rb_wr_req_desc_8_axuser_0_reg[i];
             else 
               wr_req_desc_8_axuser_0_reg[i] <= wr_req_desc_8_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_1_reg_we[i])
               wr_req_desc_8_axuser_1_reg[i] <= uc2rb_wr_req_desc_8_axuser_1_reg[i];
             else 
               wr_req_desc_8_axuser_1_reg[i] <= wr_req_desc_8_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_2_reg_we[i])
               wr_req_desc_8_axuser_2_reg[i] <= uc2rb_wr_req_desc_8_axuser_2_reg[i];
             else 
               wr_req_desc_8_axuser_2_reg[i] <= wr_req_desc_8_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_3_reg_we[i])
               wr_req_desc_8_axuser_3_reg[i] <= uc2rb_wr_req_desc_8_axuser_3_reg[i];
             else 
               wr_req_desc_8_axuser_3_reg[i] <= wr_req_desc_8_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_4_reg_we[i])
               wr_req_desc_8_axuser_4_reg[i] <= uc2rb_wr_req_desc_8_axuser_4_reg[i];
             else 
               wr_req_desc_8_axuser_4_reg[i] <= wr_req_desc_8_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_5_reg_we[i])
               wr_req_desc_8_axuser_5_reg[i] <= uc2rb_wr_req_desc_8_axuser_5_reg[i];
             else 
               wr_req_desc_8_axuser_5_reg[i] <= wr_req_desc_8_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_6_reg_we[i])
               wr_req_desc_8_axuser_6_reg[i] <= uc2rb_wr_req_desc_8_axuser_6_reg[i];
             else 
               wr_req_desc_8_axuser_6_reg[i] <= wr_req_desc_8_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_7_reg_we[i])
               wr_req_desc_8_axuser_7_reg[i] <= uc2rb_wr_req_desc_8_axuser_7_reg[i];
             else 
               wr_req_desc_8_axuser_7_reg[i] <= wr_req_desc_8_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_8_reg_we[i])
               wr_req_desc_8_axuser_8_reg[i] <= uc2rb_wr_req_desc_8_axuser_8_reg[i];
             else 
               wr_req_desc_8_axuser_8_reg[i] <= wr_req_desc_8_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_9_reg_we[i])
               wr_req_desc_8_axuser_9_reg[i] <= uc2rb_wr_req_desc_8_axuser_9_reg[i];
             else 
               wr_req_desc_8_axuser_9_reg[i] <= wr_req_desc_8_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_10_reg_we[i])
               wr_req_desc_8_axuser_10_reg[i] <= uc2rb_wr_req_desc_8_axuser_10_reg[i];
             else 
               wr_req_desc_8_axuser_10_reg[i] <= wr_req_desc_8_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_11_reg_we[i])
               wr_req_desc_8_axuser_11_reg[i] <= uc2rb_wr_req_desc_8_axuser_11_reg[i];
             else 
               wr_req_desc_8_axuser_11_reg[i] <= wr_req_desc_8_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_12_reg_we[i])
               wr_req_desc_8_axuser_12_reg[i] <= uc2rb_wr_req_desc_8_axuser_12_reg[i];
             else 
               wr_req_desc_8_axuser_12_reg[i] <= wr_req_desc_8_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_13_reg_we[i])
               wr_req_desc_8_axuser_13_reg[i] <= uc2rb_wr_req_desc_8_axuser_13_reg[i];
             else 
               wr_req_desc_8_axuser_13_reg[i] <= wr_req_desc_8_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_14_reg_we[i])
               wr_req_desc_8_axuser_14_reg[i] <= uc2rb_wr_req_desc_8_axuser_14_reg[i];
             else 
               wr_req_desc_8_axuser_14_reg[i] <= wr_req_desc_8_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_8_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_axuser_15_reg_we[i])
               wr_req_desc_8_axuser_15_reg[i] <= uc2rb_wr_req_desc_8_axuser_15_reg[i];
             else 
               wr_req_desc_8_axuser_15_reg[i] <= wr_req_desc_8_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_0_reg_we[i])
               wr_req_desc_8_wuser_0_reg[i] <= uc2rb_wr_req_desc_8_wuser_0_reg[i];
             else 
               wr_req_desc_8_wuser_0_reg[i] <= wr_req_desc_8_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_1_reg_we[i])
               wr_req_desc_8_wuser_1_reg[i] <= uc2rb_wr_req_desc_8_wuser_1_reg[i];
             else 
               wr_req_desc_8_wuser_1_reg[i] <= wr_req_desc_8_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_2_reg_we[i])
               wr_req_desc_8_wuser_2_reg[i] <= uc2rb_wr_req_desc_8_wuser_2_reg[i];
             else 
               wr_req_desc_8_wuser_2_reg[i] <= wr_req_desc_8_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_3_reg_we[i])
               wr_req_desc_8_wuser_3_reg[i] <= uc2rb_wr_req_desc_8_wuser_3_reg[i];
             else 
               wr_req_desc_8_wuser_3_reg[i] <= wr_req_desc_8_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_4_reg_we[i])
               wr_req_desc_8_wuser_4_reg[i] <= uc2rb_wr_req_desc_8_wuser_4_reg[i];
             else 
               wr_req_desc_8_wuser_4_reg[i] <= wr_req_desc_8_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_5_reg_we[i])
               wr_req_desc_8_wuser_5_reg[i] <= uc2rb_wr_req_desc_8_wuser_5_reg[i];
             else 
               wr_req_desc_8_wuser_5_reg[i] <= wr_req_desc_8_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_6_reg_we[i])
               wr_req_desc_8_wuser_6_reg[i] <= uc2rb_wr_req_desc_8_wuser_6_reg[i];
             else 
               wr_req_desc_8_wuser_6_reg[i] <= wr_req_desc_8_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_7_reg_we[i])
               wr_req_desc_8_wuser_7_reg[i] <= uc2rb_wr_req_desc_8_wuser_7_reg[i];
             else 
               wr_req_desc_8_wuser_7_reg[i] <= wr_req_desc_8_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_8_reg_we[i])
               wr_req_desc_8_wuser_8_reg[i] <= uc2rb_wr_req_desc_8_wuser_8_reg[i];
             else 
               wr_req_desc_8_wuser_8_reg[i] <= wr_req_desc_8_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_9_reg_we[i])
               wr_req_desc_8_wuser_9_reg[i] <= uc2rb_wr_req_desc_8_wuser_9_reg[i];
             else 
               wr_req_desc_8_wuser_9_reg[i] <= wr_req_desc_8_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_10_reg_we[i])
               wr_req_desc_8_wuser_10_reg[i] <= uc2rb_wr_req_desc_8_wuser_10_reg[i];
             else 
               wr_req_desc_8_wuser_10_reg[i] <= wr_req_desc_8_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_11_reg_we[i])
               wr_req_desc_8_wuser_11_reg[i] <= uc2rb_wr_req_desc_8_wuser_11_reg[i];
             else 
               wr_req_desc_8_wuser_11_reg[i] <= wr_req_desc_8_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_12_reg_we[i])
               wr_req_desc_8_wuser_12_reg[i] <= uc2rb_wr_req_desc_8_wuser_12_reg[i];
             else 
               wr_req_desc_8_wuser_12_reg[i] <= wr_req_desc_8_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_13_reg_we[i])
               wr_req_desc_8_wuser_13_reg[i] <= uc2rb_wr_req_desc_8_wuser_13_reg[i];
             else 
               wr_req_desc_8_wuser_13_reg[i] <= wr_req_desc_8_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_14_reg_we[i])
               wr_req_desc_8_wuser_14_reg[i] <= uc2rb_wr_req_desc_8_wuser_14_reg[i];
             else 
               wr_req_desc_8_wuser_14_reg[i] <= wr_req_desc_8_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_8_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_8_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_8_wuser_15_reg_we[i])
               wr_req_desc_8_wuser_15_reg[i] <= uc2rb_wr_req_desc_8_wuser_15_reg[i];
             else 
               wr_req_desc_8_wuser_15_reg[i] <= wr_req_desc_8_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_8_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_8_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_8_resp_reg_we[i])
               sn_resp_desc_8_resp_reg[i] <= uc2rb_sn_resp_desc_8_resp_reg[i];
             else 
               sn_resp_desc_8_resp_reg[i] <= sn_resp_desc_8_resp_reg[i];
        end
     end
   //RD_REQ_DESC_9_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_txn_type_reg_we[i])
               rd_req_desc_9_txn_type_reg[i] <= uc2rb_rd_req_desc_9_txn_type_reg[i];
             else 
               rd_req_desc_9_txn_type_reg[i] <= rd_req_desc_9_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_9_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_size_reg_we[i])
               rd_req_desc_9_size_reg[i] <= uc2rb_rd_req_desc_9_size_reg[i];
             else 
               rd_req_desc_9_size_reg[i] <= rd_req_desc_9_size_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axsize_reg_we[i])
               rd_req_desc_9_axsize_reg[i] <= uc2rb_rd_req_desc_9_axsize_reg[i];
             else 
               rd_req_desc_9_axsize_reg[i] <= rd_req_desc_9_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_9_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_attr_reg_we[i])
               rd_req_desc_9_attr_reg[i] <= uc2rb_rd_req_desc_9_attr_reg[i];
             else 
               rd_req_desc_9_attr_reg[i] <= rd_req_desc_9_attr_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axaddr_0_reg_we[i])
               rd_req_desc_9_axaddr_0_reg[i] <= uc2rb_rd_req_desc_9_axaddr_0_reg[i];
             else 
               rd_req_desc_9_axaddr_0_reg[i] <= rd_req_desc_9_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axaddr_1_reg_we[i])
               rd_req_desc_9_axaddr_1_reg[i] <= uc2rb_rd_req_desc_9_axaddr_1_reg[i];
             else 
               rd_req_desc_9_axaddr_1_reg[i] <= rd_req_desc_9_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axaddr_2_reg_we[i])
               rd_req_desc_9_axaddr_2_reg[i] <= uc2rb_rd_req_desc_9_axaddr_2_reg[i];
             else 
               rd_req_desc_9_axaddr_2_reg[i] <= rd_req_desc_9_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axaddr_3_reg_we[i])
               rd_req_desc_9_axaddr_3_reg[i] <= uc2rb_rd_req_desc_9_axaddr_3_reg[i];
             else 
               rd_req_desc_9_axaddr_3_reg[i] <= rd_req_desc_9_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axid_0_reg_we[i])
               rd_req_desc_9_axid_0_reg[i] <= uc2rb_rd_req_desc_9_axid_0_reg[i];
             else 
               rd_req_desc_9_axid_0_reg[i] <= rd_req_desc_9_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axid_1_reg_we[i])
               rd_req_desc_9_axid_1_reg[i] <= uc2rb_rd_req_desc_9_axid_1_reg[i];
             else 
               rd_req_desc_9_axid_1_reg[i] <= rd_req_desc_9_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axid_2_reg_we[i])
               rd_req_desc_9_axid_2_reg[i] <= uc2rb_rd_req_desc_9_axid_2_reg[i];
             else 
               rd_req_desc_9_axid_2_reg[i] <= rd_req_desc_9_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axid_3_reg_we[i])
               rd_req_desc_9_axid_3_reg[i] <= uc2rb_rd_req_desc_9_axid_3_reg[i];
             else 
               rd_req_desc_9_axid_3_reg[i] <= rd_req_desc_9_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_0_reg_we[i])
               rd_req_desc_9_axuser_0_reg[i] <= uc2rb_rd_req_desc_9_axuser_0_reg[i];
             else 
               rd_req_desc_9_axuser_0_reg[i] <= rd_req_desc_9_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_1_reg_we[i])
               rd_req_desc_9_axuser_1_reg[i] <= uc2rb_rd_req_desc_9_axuser_1_reg[i];
             else 
               rd_req_desc_9_axuser_1_reg[i] <= rd_req_desc_9_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_2_reg_we[i])
               rd_req_desc_9_axuser_2_reg[i] <= uc2rb_rd_req_desc_9_axuser_2_reg[i];
             else 
               rd_req_desc_9_axuser_2_reg[i] <= rd_req_desc_9_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_3_reg_we[i])
               rd_req_desc_9_axuser_3_reg[i] <= uc2rb_rd_req_desc_9_axuser_3_reg[i];
             else 
               rd_req_desc_9_axuser_3_reg[i] <= rd_req_desc_9_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_4_reg_we[i])
               rd_req_desc_9_axuser_4_reg[i] <= uc2rb_rd_req_desc_9_axuser_4_reg[i];
             else 
               rd_req_desc_9_axuser_4_reg[i] <= rd_req_desc_9_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_5_reg_we[i])
               rd_req_desc_9_axuser_5_reg[i] <= uc2rb_rd_req_desc_9_axuser_5_reg[i];
             else 
               rd_req_desc_9_axuser_5_reg[i] <= rd_req_desc_9_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_6_reg_we[i])
               rd_req_desc_9_axuser_6_reg[i] <= uc2rb_rd_req_desc_9_axuser_6_reg[i];
             else 
               rd_req_desc_9_axuser_6_reg[i] <= rd_req_desc_9_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_7_reg_we[i])
               rd_req_desc_9_axuser_7_reg[i] <= uc2rb_rd_req_desc_9_axuser_7_reg[i];
             else 
               rd_req_desc_9_axuser_7_reg[i] <= rd_req_desc_9_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_8_reg_we[i])
               rd_req_desc_9_axuser_8_reg[i] <= uc2rb_rd_req_desc_9_axuser_8_reg[i];
             else 
               rd_req_desc_9_axuser_8_reg[i] <= rd_req_desc_9_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_9_reg_we[i])
               rd_req_desc_9_axuser_9_reg[i] <= uc2rb_rd_req_desc_9_axuser_9_reg[i];
             else 
               rd_req_desc_9_axuser_9_reg[i] <= rd_req_desc_9_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_10_reg_we[i])
               rd_req_desc_9_axuser_10_reg[i] <= uc2rb_rd_req_desc_9_axuser_10_reg[i];
             else 
               rd_req_desc_9_axuser_10_reg[i] <= rd_req_desc_9_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_11_reg_we[i])
               rd_req_desc_9_axuser_11_reg[i] <= uc2rb_rd_req_desc_9_axuser_11_reg[i];
             else 
               rd_req_desc_9_axuser_11_reg[i] <= rd_req_desc_9_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_12_reg_we[i])
               rd_req_desc_9_axuser_12_reg[i] <= uc2rb_rd_req_desc_9_axuser_12_reg[i];
             else 
               rd_req_desc_9_axuser_12_reg[i] <= rd_req_desc_9_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_13_reg_we[i])
               rd_req_desc_9_axuser_13_reg[i] <= uc2rb_rd_req_desc_9_axuser_13_reg[i];
             else 
               rd_req_desc_9_axuser_13_reg[i] <= rd_req_desc_9_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_14_reg_we[i])
               rd_req_desc_9_axuser_14_reg[i] <= uc2rb_rd_req_desc_9_axuser_14_reg[i];
             else 
               rd_req_desc_9_axuser_14_reg[i] <= rd_req_desc_9_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_9_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_9_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_9_axuser_15_reg_we[i])
               rd_req_desc_9_axuser_15_reg[i] <= uc2rb_rd_req_desc_9_axuser_15_reg[i];
             else 
               rd_req_desc_9_axuser_15_reg[i] <= rd_req_desc_9_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_9_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_txn_type_reg_we[i])
               wr_req_desc_9_txn_type_reg[i] <= uc2rb_wr_req_desc_9_txn_type_reg[i];
             else 
               wr_req_desc_9_txn_type_reg[i] <= wr_req_desc_9_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_9_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_size_reg_we[i])
               wr_req_desc_9_size_reg[i] <= uc2rb_wr_req_desc_9_size_reg[i];
             else 
               wr_req_desc_9_size_reg[i] <= wr_req_desc_9_size_reg[i];
        end
     end
   //WR_REQ_DESC_9_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_data_offset_reg_we[i])
               wr_req_desc_9_data_offset_reg[i] <= uc2rb_wr_req_desc_9_data_offset_reg[i];
             else 
               wr_req_desc_9_data_offset_reg[i] <= wr_req_desc_9_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axsize_reg_we[i])
               wr_req_desc_9_axsize_reg[i] <= uc2rb_wr_req_desc_9_axsize_reg[i];
             else 
               wr_req_desc_9_axsize_reg[i] <= wr_req_desc_9_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_9_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_attr_reg_we[i])
               wr_req_desc_9_attr_reg[i] <= uc2rb_wr_req_desc_9_attr_reg[i];
             else 
               wr_req_desc_9_attr_reg[i] <= wr_req_desc_9_attr_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axaddr_0_reg_we[i])
               wr_req_desc_9_axaddr_0_reg[i] <= uc2rb_wr_req_desc_9_axaddr_0_reg[i];
             else 
               wr_req_desc_9_axaddr_0_reg[i] <= wr_req_desc_9_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axaddr_1_reg_we[i])
               wr_req_desc_9_axaddr_1_reg[i] <= uc2rb_wr_req_desc_9_axaddr_1_reg[i];
             else 
               wr_req_desc_9_axaddr_1_reg[i] <= wr_req_desc_9_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axaddr_2_reg_we[i])
               wr_req_desc_9_axaddr_2_reg[i] <= uc2rb_wr_req_desc_9_axaddr_2_reg[i];
             else 
               wr_req_desc_9_axaddr_2_reg[i] <= wr_req_desc_9_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axaddr_3_reg_we[i])
               wr_req_desc_9_axaddr_3_reg[i] <= uc2rb_wr_req_desc_9_axaddr_3_reg[i];
             else 
               wr_req_desc_9_axaddr_3_reg[i] <= wr_req_desc_9_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axid_0_reg_we[i])
               wr_req_desc_9_axid_0_reg[i] <= uc2rb_wr_req_desc_9_axid_0_reg[i];
             else 
               wr_req_desc_9_axid_0_reg[i] <= wr_req_desc_9_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axid_1_reg_we[i])
               wr_req_desc_9_axid_1_reg[i] <= uc2rb_wr_req_desc_9_axid_1_reg[i];
             else 
               wr_req_desc_9_axid_1_reg[i] <= wr_req_desc_9_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axid_2_reg_we[i])
               wr_req_desc_9_axid_2_reg[i] <= uc2rb_wr_req_desc_9_axid_2_reg[i];
             else 
               wr_req_desc_9_axid_2_reg[i] <= wr_req_desc_9_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axid_3_reg_we[i])
               wr_req_desc_9_axid_3_reg[i] <= uc2rb_wr_req_desc_9_axid_3_reg[i];
             else 
               wr_req_desc_9_axid_3_reg[i] <= wr_req_desc_9_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_0_reg_we[i])
               wr_req_desc_9_axuser_0_reg[i] <= uc2rb_wr_req_desc_9_axuser_0_reg[i];
             else 
               wr_req_desc_9_axuser_0_reg[i] <= wr_req_desc_9_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_1_reg_we[i])
               wr_req_desc_9_axuser_1_reg[i] <= uc2rb_wr_req_desc_9_axuser_1_reg[i];
             else 
               wr_req_desc_9_axuser_1_reg[i] <= wr_req_desc_9_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_2_reg_we[i])
               wr_req_desc_9_axuser_2_reg[i] <= uc2rb_wr_req_desc_9_axuser_2_reg[i];
             else 
               wr_req_desc_9_axuser_2_reg[i] <= wr_req_desc_9_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_3_reg_we[i])
               wr_req_desc_9_axuser_3_reg[i] <= uc2rb_wr_req_desc_9_axuser_3_reg[i];
             else 
               wr_req_desc_9_axuser_3_reg[i] <= wr_req_desc_9_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_4_reg_we[i])
               wr_req_desc_9_axuser_4_reg[i] <= uc2rb_wr_req_desc_9_axuser_4_reg[i];
             else 
               wr_req_desc_9_axuser_4_reg[i] <= wr_req_desc_9_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_5_reg_we[i])
               wr_req_desc_9_axuser_5_reg[i] <= uc2rb_wr_req_desc_9_axuser_5_reg[i];
             else 
               wr_req_desc_9_axuser_5_reg[i] <= wr_req_desc_9_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_6_reg_we[i])
               wr_req_desc_9_axuser_6_reg[i] <= uc2rb_wr_req_desc_9_axuser_6_reg[i];
             else 
               wr_req_desc_9_axuser_6_reg[i] <= wr_req_desc_9_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_7_reg_we[i])
               wr_req_desc_9_axuser_7_reg[i] <= uc2rb_wr_req_desc_9_axuser_7_reg[i];
             else 
               wr_req_desc_9_axuser_7_reg[i] <= wr_req_desc_9_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_8_reg_we[i])
               wr_req_desc_9_axuser_8_reg[i] <= uc2rb_wr_req_desc_9_axuser_8_reg[i];
             else 
               wr_req_desc_9_axuser_8_reg[i] <= wr_req_desc_9_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_9_reg_we[i])
               wr_req_desc_9_axuser_9_reg[i] <= uc2rb_wr_req_desc_9_axuser_9_reg[i];
             else 
               wr_req_desc_9_axuser_9_reg[i] <= wr_req_desc_9_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_10_reg_we[i])
               wr_req_desc_9_axuser_10_reg[i] <= uc2rb_wr_req_desc_9_axuser_10_reg[i];
             else 
               wr_req_desc_9_axuser_10_reg[i] <= wr_req_desc_9_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_11_reg_we[i])
               wr_req_desc_9_axuser_11_reg[i] <= uc2rb_wr_req_desc_9_axuser_11_reg[i];
             else 
               wr_req_desc_9_axuser_11_reg[i] <= wr_req_desc_9_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_12_reg_we[i])
               wr_req_desc_9_axuser_12_reg[i] <= uc2rb_wr_req_desc_9_axuser_12_reg[i];
             else 
               wr_req_desc_9_axuser_12_reg[i] <= wr_req_desc_9_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_13_reg_we[i])
               wr_req_desc_9_axuser_13_reg[i] <= uc2rb_wr_req_desc_9_axuser_13_reg[i];
             else 
               wr_req_desc_9_axuser_13_reg[i] <= wr_req_desc_9_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_14_reg_we[i])
               wr_req_desc_9_axuser_14_reg[i] <= uc2rb_wr_req_desc_9_axuser_14_reg[i];
             else 
               wr_req_desc_9_axuser_14_reg[i] <= wr_req_desc_9_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_9_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_axuser_15_reg_we[i])
               wr_req_desc_9_axuser_15_reg[i] <= uc2rb_wr_req_desc_9_axuser_15_reg[i];
             else 
               wr_req_desc_9_axuser_15_reg[i] <= wr_req_desc_9_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_0_reg_we[i])
               wr_req_desc_9_wuser_0_reg[i] <= uc2rb_wr_req_desc_9_wuser_0_reg[i];
             else 
               wr_req_desc_9_wuser_0_reg[i] <= wr_req_desc_9_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_1_reg_we[i])
               wr_req_desc_9_wuser_1_reg[i] <= uc2rb_wr_req_desc_9_wuser_1_reg[i];
             else 
               wr_req_desc_9_wuser_1_reg[i] <= wr_req_desc_9_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_2_reg_we[i])
               wr_req_desc_9_wuser_2_reg[i] <= uc2rb_wr_req_desc_9_wuser_2_reg[i];
             else 
               wr_req_desc_9_wuser_2_reg[i] <= wr_req_desc_9_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_3_reg_we[i])
               wr_req_desc_9_wuser_3_reg[i] <= uc2rb_wr_req_desc_9_wuser_3_reg[i];
             else 
               wr_req_desc_9_wuser_3_reg[i] <= wr_req_desc_9_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_4_reg_we[i])
               wr_req_desc_9_wuser_4_reg[i] <= uc2rb_wr_req_desc_9_wuser_4_reg[i];
             else 
               wr_req_desc_9_wuser_4_reg[i] <= wr_req_desc_9_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_5_reg_we[i])
               wr_req_desc_9_wuser_5_reg[i] <= uc2rb_wr_req_desc_9_wuser_5_reg[i];
             else 
               wr_req_desc_9_wuser_5_reg[i] <= wr_req_desc_9_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_6_reg_we[i])
               wr_req_desc_9_wuser_6_reg[i] <= uc2rb_wr_req_desc_9_wuser_6_reg[i];
             else 
               wr_req_desc_9_wuser_6_reg[i] <= wr_req_desc_9_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_7_reg_we[i])
               wr_req_desc_9_wuser_7_reg[i] <= uc2rb_wr_req_desc_9_wuser_7_reg[i];
             else 
               wr_req_desc_9_wuser_7_reg[i] <= wr_req_desc_9_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_8_reg_we[i])
               wr_req_desc_9_wuser_8_reg[i] <= uc2rb_wr_req_desc_9_wuser_8_reg[i];
             else 
               wr_req_desc_9_wuser_8_reg[i] <= wr_req_desc_9_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_9_reg_we[i])
               wr_req_desc_9_wuser_9_reg[i] <= uc2rb_wr_req_desc_9_wuser_9_reg[i];
             else 
               wr_req_desc_9_wuser_9_reg[i] <= wr_req_desc_9_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_10_reg_we[i])
               wr_req_desc_9_wuser_10_reg[i] <= uc2rb_wr_req_desc_9_wuser_10_reg[i];
             else 
               wr_req_desc_9_wuser_10_reg[i] <= wr_req_desc_9_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_11_reg_we[i])
               wr_req_desc_9_wuser_11_reg[i] <= uc2rb_wr_req_desc_9_wuser_11_reg[i];
             else 
               wr_req_desc_9_wuser_11_reg[i] <= wr_req_desc_9_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_12_reg_we[i])
               wr_req_desc_9_wuser_12_reg[i] <= uc2rb_wr_req_desc_9_wuser_12_reg[i];
             else 
               wr_req_desc_9_wuser_12_reg[i] <= wr_req_desc_9_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_13_reg_we[i])
               wr_req_desc_9_wuser_13_reg[i] <= uc2rb_wr_req_desc_9_wuser_13_reg[i];
             else 
               wr_req_desc_9_wuser_13_reg[i] <= wr_req_desc_9_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_14_reg_we[i])
               wr_req_desc_9_wuser_14_reg[i] <= uc2rb_wr_req_desc_9_wuser_14_reg[i];
             else 
               wr_req_desc_9_wuser_14_reg[i] <= wr_req_desc_9_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_9_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_9_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_9_wuser_15_reg_we[i])
               wr_req_desc_9_wuser_15_reg[i] <= uc2rb_wr_req_desc_9_wuser_15_reg[i];
             else 
               wr_req_desc_9_wuser_15_reg[i] <= wr_req_desc_9_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_9_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_9_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_9_resp_reg_we[i])
               sn_resp_desc_9_resp_reg[i] <= uc2rb_sn_resp_desc_9_resp_reg[i];
             else 
               sn_resp_desc_9_resp_reg[i] <= sn_resp_desc_9_resp_reg[i];
        end
     end
   //RD_REQ_DESC_A_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_txn_type_reg_we[i])
               rd_req_desc_a_txn_type_reg[i] <= uc2rb_rd_req_desc_a_txn_type_reg[i];
             else 
               rd_req_desc_a_txn_type_reg[i] <= rd_req_desc_a_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_A_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_size_reg_we[i])
               rd_req_desc_a_size_reg[i] <= uc2rb_rd_req_desc_a_size_reg[i];
             else 
               rd_req_desc_a_size_reg[i] <= rd_req_desc_a_size_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axsize_reg_we[i])
               rd_req_desc_a_axsize_reg[i] <= uc2rb_rd_req_desc_a_axsize_reg[i];
             else 
               rd_req_desc_a_axsize_reg[i] <= rd_req_desc_a_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_A_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_attr_reg_we[i])
               rd_req_desc_a_attr_reg[i] <= uc2rb_rd_req_desc_a_attr_reg[i];
             else 
               rd_req_desc_a_attr_reg[i] <= rd_req_desc_a_attr_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axaddr_0_reg_we[i])
               rd_req_desc_a_axaddr_0_reg[i] <= uc2rb_rd_req_desc_a_axaddr_0_reg[i];
             else 
               rd_req_desc_a_axaddr_0_reg[i] <= rd_req_desc_a_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axaddr_1_reg_we[i])
               rd_req_desc_a_axaddr_1_reg[i] <= uc2rb_rd_req_desc_a_axaddr_1_reg[i];
             else 
               rd_req_desc_a_axaddr_1_reg[i] <= rd_req_desc_a_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axaddr_2_reg_we[i])
               rd_req_desc_a_axaddr_2_reg[i] <= uc2rb_rd_req_desc_a_axaddr_2_reg[i];
             else 
               rd_req_desc_a_axaddr_2_reg[i] <= rd_req_desc_a_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axaddr_3_reg_we[i])
               rd_req_desc_a_axaddr_3_reg[i] <= uc2rb_rd_req_desc_a_axaddr_3_reg[i];
             else 
               rd_req_desc_a_axaddr_3_reg[i] <= rd_req_desc_a_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axid_0_reg_we[i])
               rd_req_desc_a_axid_0_reg[i] <= uc2rb_rd_req_desc_a_axid_0_reg[i];
             else 
               rd_req_desc_a_axid_0_reg[i] <= rd_req_desc_a_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axid_1_reg_we[i])
               rd_req_desc_a_axid_1_reg[i] <= uc2rb_rd_req_desc_a_axid_1_reg[i];
             else 
               rd_req_desc_a_axid_1_reg[i] <= rd_req_desc_a_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axid_2_reg_we[i])
               rd_req_desc_a_axid_2_reg[i] <= uc2rb_rd_req_desc_a_axid_2_reg[i];
             else 
               rd_req_desc_a_axid_2_reg[i] <= rd_req_desc_a_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axid_3_reg_we[i])
               rd_req_desc_a_axid_3_reg[i] <= uc2rb_rd_req_desc_a_axid_3_reg[i];
             else 
               rd_req_desc_a_axid_3_reg[i] <= rd_req_desc_a_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_0_reg_we[i])
               rd_req_desc_a_axuser_0_reg[i] <= uc2rb_rd_req_desc_a_axuser_0_reg[i];
             else 
               rd_req_desc_a_axuser_0_reg[i] <= rd_req_desc_a_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_1_reg_we[i])
               rd_req_desc_a_axuser_1_reg[i] <= uc2rb_rd_req_desc_a_axuser_1_reg[i];
             else 
               rd_req_desc_a_axuser_1_reg[i] <= rd_req_desc_a_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_2_reg_we[i])
               rd_req_desc_a_axuser_2_reg[i] <= uc2rb_rd_req_desc_a_axuser_2_reg[i];
             else 
               rd_req_desc_a_axuser_2_reg[i] <= rd_req_desc_a_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_3_reg_we[i])
               rd_req_desc_a_axuser_3_reg[i] <= uc2rb_rd_req_desc_a_axuser_3_reg[i];
             else 
               rd_req_desc_a_axuser_3_reg[i] <= rd_req_desc_a_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_4_reg_we[i])
               rd_req_desc_a_axuser_4_reg[i] <= uc2rb_rd_req_desc_a_axuser_4_reg[i];
             else 
               rd_req_desc_a_axuser_4_reg[i] <= rd_req_desc_a_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_5_reg_we[i])
               rd_req_desc_a_axuser_5_reg[i] <= uc2rb_rd_req_desc_a_axuser_5_reg[i];
             else 
               rd_req_desc_a_axuser_5_reg[i] <= rd_req_desc_a_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_6_reg_we[i])
               rd_req_desc_a_axuser_6_reg[i] <= uc2rb_rd_req_desc_a_axuser_6_reg[i];
             else 
               rd_req_desc_a_axuser_6_reg[i] <= rd_req_desc_a_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_7_reg_we[i])
               rd_req_desc_a_axuser_7_reg[i] <= uc2rb_rd_req_desc_a_axuser_7_reg[i];
             else 
               rd_req_desc_a_axuser_7_reg[i] <= rd_req_desc_a_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_8_reg_we[i])
               rd_req_desc_a_axuser_8_reg[i] <= uc2rb_rd_req_desc_a_axuser_8_reg[i];
             else 
               rd_req_desc_a_axuser_8_reg[i] <= rd_req_desc_a_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_9_reg_we[i])
               rd_req_desc_a_axuser_9_reg[i] <= uc2rb_rd_req_desc_a_axuser_9_reg[i];
             else 
               rd_req_desc_a_axuser_9_reg[i] <= rd_req_desc_a_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_10_reg_we[i])
               rd_req_desc_a_axuser_10_reg[i] <= uc2rb_rd_req_desc_a_axuser_10_reg[i];
             else 
               rd_req_desc_a_axuser_10_reg[i] <= rd_req_desc_a_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_11_reg_we[i])
               rd_req_desc_a_axuser_11_reg[i] <= uc2rb_rd_req_desc_a_axuser_11_reg[i];
             else 
               rd_req_desc_a_axuser_11_reg[i] <= rd_req_desc_a_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_12_reg_we[i])
               rd_req_desc_a_axuser_12_reg[i] <= uc2rb_rd_req_desc_a_axuser_12_reg[i];
             else 
               rd_req_desc_a_axuser_12_reg[i] <= rd_req_desc_a_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_13_reg_we[i])
               rd_req_desc_a_axuser_13_reg[i] <= uc2rb_rd_req_desc_a_axuser_13_reg[i];
             else 
               rd_req_desc_a_axuser_13_reg[i] <= rd_req_desc_a_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_14_reg_we[i])
               rd_req_desc_a_axuser_14_reg[i] <= uc2rb_rd_req_desc_a_axuser_14_reg[i];
             else 
               rd_req_desc_a_axuser_14_reg[i] <= rd_req_desc_a_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_A_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_a_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_a_axuser_15_reg_we[i])
               rd_req_desc_a_axuser_15_reg[i] <= uc2rb_rd_req_desc_a_axuser_15_reg[i];
             else 
               rd_req_desc_a_axuser_15_reg[i] <= rd_req_desc_a_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_A_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_txn_type_reg_we[i])
               wr_req_desc_a_txn_type_reg[i] <= uc2rb_wr_req_desc_a_txn_type_reg[i];
             else 
               wr_req_desc_a_txn_type_reg[i] <= wr_req_desc_a_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_A_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_size_reg_we[i])
               wr_req_desc_a_size_reg[i] <= uc2rb_wr_req_desc_a_size_reg[i];
             else 
               wr_req_desc_a_size_reg[i] <= wr_req_desc_a_size_reg[i];
        end
     end
   //WR_REQ_DESC_A_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_data_offset_reg_we[i])
               wr_req_desc_a_data_offset_reg[i] <= uc2rb_wr_req_desc_a_data_offset_reg[i];
             else 
               wr_req_desc_a_data_offset_reg[i] <= wr_req_desc_a_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axsize_reg_we[i])
               wr_req_desc_a_axsize_reg[i] <= uc2rb_wr_req_desc_a_axsize_reg[i];
             else 
               wr_req_desc_a_axsize_reg[i] <= wr_req_desc_a_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_A_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_attr_reg_we[i])
               wr_req_desc_a_attr_reg[i] <= uc2rb_wr_req_desc_a_attr_reg[i];
             else 
               wr_req_desc_a_attr_reg[i] <= wr_req_desc_a_attr_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axaddr_0_reg_we[i])
               wr_req_desc_a_axaddr_0_reg[i] <= uc2rb_wr_req_desc_a_axaddr_0_reg[i];
             else 
               wr_req_desc_a_axaddr_0_reg[i] <= wr_req_desc_a_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axaddr_1_reg_we[i])
               wr_req_desc_a_axaddr_1_reg[i] <= uc2rb_wr_req_desc_a_axaddr_1_reg[i];
             else 
               wr_req_desc_a_axaddr_1_reg[i] <= wr_req_desc_a_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axaddr_2_reg_we[i])
               wr_req_desc_a_axaddr_2_reg[i] <= uc2rb_wr_req_desc_a_axaddr_2_reg[i];
             else 
               wr_req_desc_a_axaddr_2_reg[i] <= wr_req_desc_a_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axaddr_3_reg_we[i])
               wr_req_desc_a_axaddr_3_reg[i] <= uc2rb_wr_req_desc_a_axaddr_3_reg[i];
             else 
               wr_req_desc_a_axaddr_3_reg[i] <= wr_req_desc_a_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axid_0_reg_we[i])
               wr_req_desc_a_axid_0_reg[i] <= uc2rb_wr_req_desc_a_axid_0_reg[i];
             else 
               wr_req_desc_a_axid_0_reg[i] <= wr_req_desc_a_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axid_1_reg_we[i])
               wr_req_desc_a_axid_1_reg[i] <= uc2rb_wr_req_desc_a_axid_1_reg[i];
             else 
               wr_req_desc_a_axid_1_reg[i] <= wr_req_desc_a_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axid_2_reg_we[i])
               wr_req_desc_a_axid_2_reg[i] <= uc2rb_wr_req_desc_a_axid_2_reg[i];
             else 
               wr_req_desc_a_axid_2_reg[i] <= wr_req_desc_a_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axid_3_reg_we[i])
               wr_req_desc_a_axid_3_reg[i] <= uc2rb_wr_req_desc_a_axid_3_reg[i];
             else 
               wr_req_desc_a_axid_3_reg[i] <= wr_req_desc_a_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_0_reg_we[i])
               wr_req_desc_a_axuser_0_reg[i] <= uc2rb_wr_req_desc_a_axuser_0_reg[i];
             else 
               wr_req_desc_a_axuser_0_reg[i] <= wr_req_desc_a_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_1_reg_we[i])
               wr_req_desc_a_axuser_1_reg[i] <= uc2rb_wr_req_desc_a_axuser_1_reg[i];
             else 
               wr_req_desc_a_axuser_1_reg[i] <= wr_req_desc_a_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_2_reg_we[i])
               wr_req_desc_a_axuser_2_reg[i] <= uc2rb_wr_req_desc_a_axuser_2_reg[i];
             else 
               wr_req_desc_a_axuser_2_reg[i] <= wr_req_desc_a_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_3_reg_we[i])
               wr_req_desc_a_axuser_3_reg[i] <= uc2rb_wr_req_desc_a_axuser_3_reg[i];
             else 
               wr_req_desc_a_axuser_3_reg[i] <= wr_req_desc_a_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_4_reg_we[i])
               wr_req_desc_a_axuser_4_reg[i] <= uc2rb_wr_req_desc_a_axuser_4_reg[i];
             else 
               wr_req_desc_a_axuser_4_reg[i] <= wr_req_desc_a_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_5_reg_we[i])
               wr_req_desc_a_axuser_5_reg[i] <= uc2rb_wr_req_desc_a_axuser_5_reg[i];
             else 
               wr_req_desc_a_axuser_5_reg[i] <= wr_req_desc_a_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_6_reg_we[i])
               wr_req_desc_a_axuser_6_reg[i] <= uc2rb_wr_req_desc_a_axuser_6_reg[i];
             else 
               wr_req_desc_a_axuser_6_reg[i] <= wr_req_desc_a_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_7_reg_we[i])
               wr_req_desc_a_axuser_7_reg[i] <= uc2rb_wr_req_desc_a_axuser_7_reg[i];
             else 
               wr_req_desc_a_axuser_7_reg[i] <= wr_req_desc_a_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_8_reg_we[i])
               wr_req_desc_a_axuser_8_reg[i] <= uc2rb_wr_req_desc_a_axuser_8_reg[i];
             else 
               wr_req_desc_a_axuser_8_reg[i] <= wr_req_desc_a_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_9_reg_we[i])
               wr_req_desc_a_axuser_9_reg[i] <= uc2rb_wr_req_desc_a_axuser_9_reg[i];
             else 
               wr_req_desc_a_axuser_9_reg[i] <= wr_req_desc_a_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_10_reg_we[i])
               wr_req_desc_a_axuser_10_reg[i] <= uc2rb_wr_req_desc_a_axuser_10_reg[i];
             else 
               wr_req_desc_a_axuser_10_reg[i] <= wr_req_desc_a_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_11_reg_we[i])
               wr_req_desc_a_axuser_11_reg[i] <= uc2rb_wr_req_desc_a_axuser_11_reg[i];
             else 
               wr_req_desc_a_axuser_11_reg[i] <= wr_req_desc_a_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_12_reg_we[i])
               wr_req_desc_a_axuser_12_reg[i] <= uc2rb_wr_req_desc_a_axuser_12_reg[i];
             else 
               wr_req_desc_a_axuser_12_reg[i] <= wr_req_desc_a_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_13_reg_we[i])
               wr_req_desc_a_axuser_13_reg[i] <= uc2rb_wr_req_desc_a_axuser_13_reg[i];
             else 
               wr_req_desc_a_axuser_13_reg[i] <= wr_req_desc_a_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_14_reg_we[i])
               wr_req_desc_a_axuser_14_reg[i] <= uc2rb_wr_req_desc_a_axuser_14_reg[i];
             else 
               wr_req_desc_a_axuser_14_reg[i] <= wr_req_desc_a_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_A_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_axuser_15_reg_we[i])
               wr_req_desc_a_axuser_15_reg[i] <= uc2rb_wr_req_desc_a_axuser_15_reg[i];
             else 
               wr_req_desc_a_axuser_15_reg[i] <= wr_req_desc_a_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_0_reg_we[i])
               wr_req_desc_a_wuser_0_reg[i] <= uc2rb_wr_req_desc_a_wuser_0_reg[i];
             else 
               wr_req_desc_a_wuser_0_reg[i] <= wr_req_desc_a_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_1_reg_we[i])
               wr_req_desc_a_wuser_1_reg[i] <= uc2rb_wr_req_desc_a_wuser_1_reg[i];
             else 
               wr_req_desc_a_wuser_1_reg[i] <= wr_req_desc_a_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_2_reg_we[i])
               wr_req_desc_a_wuser_2_reg[i] <= uc2rb_wr_req_desc_a_wuser_2_reg[i];
             else 
               wr_req_desc_a_wuser_2_reg[i] <= wr_req_desc_a_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_3_reg_we[i])
               wr_req_desc_a_wuser_3_reg[i] <= uc2rb_wr_req_desc_a_wuser_3_reg[i];
             else 
               wr_req_desc_a_wuser_3_reg[i] <= wr_req_desc_a_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_4_reg_we[i])
               wr_req_desc_a_wuser_4_reg[i] <= uc2rb_wr_req_desc_a_wuser_4_reg[i];
             else 
               wr_req_desc_a_wuser_4_reg[i] <= wr_req_desc_a_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_5_reg_we[i])
               wr_req_desc_a_wuser_5_reg[i] <= uc2rb_wr_req_desc_a_wuser_5_reg[i];
             else 
               wr_req_desc_a_wuser_5_reg[i] <= wr_req_desc_a_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_6_reg_we[i])
               wr_req_desc_a_wuser_6_reg[i] <= uc2rb_wr_req_desc_a_wuser_6_reg[i];
             else 
               wr_req_desc_a_wuser_6_reg[i] <= wr_req_desc_a_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_7_reg_we[i])
               wr_req_desc_a_wuser_7_reg[i] <= uc2rb_wr_req_desc_a_wuser_7_reg[i];
             else 
               wr_req_desc_a_wuser_7_reg[i] <= wr_req_desc_a_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_8_reg_we[i])
               wr_req_desc_a_wuser_8_reg[i] <= uc2rb_wr_req_desc_a_wuser_8_reg[i];
             else 
               wr_req_desc_a_wuser_8_reg[i] <= wr_req_desc_a_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_9_reg_we[i])
               wr_req_desc_a_wuser_9_reg[i] <= uc2rb_wr_req_desc_a_wuser_9_reg[i];
             else 
               wr_req_desc_a_wuser_9_reg[i] <= wr_req_desc_a_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_10_reg_we[i])
               wr_req_desc_a_wuser_10_reg[i] <= uc2rb_wr_req_desc_a_wuser_10_reg[i];
             else 
               wr_req_desc_a_wuser_10_reg[i] <= wr_req_desc_a_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_11_reg_we[i])
               wr_req_desc_a_wuser_11_reg[i] <= uc2rb_wr_req_desc_a_wuser_11_reg[i];
             else 
               wr_req_desc_a_wuser_11_reg[i] <= wr_req_desc_a_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_12_reg_we[i])
               wr_req_desc_a_wuser_12_reg[i] <= uc2rb_wr_req_desc_a_wuser_12_reg[i];
             else 
               wr_req_desc_a_wuser_12_reg[i] <= wr_req_desc_a_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_13_reg_we[i])
               wr_req_desc_a_wuser_13_reg[i] <= uc2rb_wr_req_desc_a_wuser_13_reg[i];
             else 
               wr_req_desc_a_wuser_13_reg[i] <= wr_req_desc_a_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_14_reg_we[i])
               wr_req_desc_a_wuser_14_reg[i] <= uc2rb_wr_req_desc_a_wuser_14_reg[i];
             else 
               wr_req_desc_a_wuser_14_reg[i] <= wr_req_desc_a_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_A_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_a_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_a_wuser_15_reg_we[i])
               wr_req_desc_a_wuser_15_reg[i] <= uc2rb_wr_req_desc_a_wuser_15_reg[i];
             else 
               wr_req_desc_a_wuser_15_reg[i] <= wr_req_desc_a_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_A_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_a_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_a_resp_reg_we[i])
               sn_resp_desc_a_resp_reg[i] <= uc2rb_sn_resp_desc_a_resp_reg[i];
             else 
               sn_resp_desc_a_resp_reg[i] <= sn_resp_desc_a_resp_reg[i];
        end
     end
   //RD_REQ_DESC_B_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_txn_type_reg_we[i])
               rd_req_desc_b_txn_type_reg[i] <= uc2rb_rd_req_desc_b_txn_type_reg[i];
             else 
               rd_req_desc_b_txn_type_reg[i] <= rd_req_desc_b_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_B_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_size_reg_we[i])
               rd_req_desc_b_size_reg[i] <= uc2rb_rd_req_desc_b_size_reg[i];
             else 
               rd_req_desc_b_size_reg[i] <= rd_req_desc_b_size_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axsize_reg_we[i])
               rd_req_desc_b_axsize_reg[i] <= uc2rb_rd_req_desc_b_axsize_reg[i];
             else 
               rd_req_desc_b_axsize_reg[i] <= rd_req_desc_b_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_B_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_attr_reg_we[i])
               rd_req_desc_b_attr_reg[i] <= uc2rb_rd_req_desc_b_attr_reg[i];
             else 
               rd_req_desc_b_attr_reg[i] <= rd_req_desc_b_attr_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axaddr_0_reg_we[i])
               rd_req_desc_b_axaddr_0_reg[i] <= uc2rb_rd_req_desc_b_axaddr_0_reg[i];
             else 
               rd_req_desc_b_axaddr_0_reg[i] <= rd_req_desc_b_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axaddr_1_reg_we[i])
               rd_req_desc_b_axaddr_1_reg[i] <= uc2rb_rd_req_desc_b_axaddr_1_reg[i];
             else 
               rd_req_desc_b_axaddr_1_reg[i] <= rd_req_desc_b_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axaddr_2_reg_we[i])
               rd_req_desc_b_axaddr_2_reg[i] <= uc2rb_rd_req_desc_b_axaddr_2_reg[i];
             else 
               rd_req_desc_b_axaddr_2_reg[i] <= rd_req_desc_b_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axaddr_3_reg_we[i])
               rd_req_desc_b_axaddr_3_reg[i] <= uc2rb_rd_req_desc_b_axaddr_3_reg[i];
             else 
               rd_req_desc_b_axaddr_3_reg[i] <= rd_req_desc_b_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axid_0_reg_we[i])
               rd_req_desc_b_axid_0_reg[i] <= uc2rb_rd_req_desc_b_axid_0_reg[i];
             else 
               rd_req_desc_b_axid_0_reg[i] <= rd_req_desc_b_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axid_1_reg_we[i])
               rd_req_desc_b_axid_1_reg[i] <= uc2rb_rd_req_desc_b_axid_1_reg[i];
             else 
               rd_req_desc_b_axid_1_reg[i] <= rd_req_desc_b_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axid_2_reg_we[i])
               rd_req_desc_b_axid_2_reg[i] <= uc2rb_rd_req_desc_b_axid_2_reg[i];
             else 
               rd_req_desc_b_axid_2_reg[i] <= rd_req_desc_b_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axid_3_reg_we[i])
               rd_req_desc_b_axid_3_reg[i] <= uc2rb_rd_req_desc_b_axid_3_reg[i];
             else 
               rd_req_desc_b_axid_3_reg[i] <= rd_req_desc_b_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_0_reg_we[i])
               rd_req_desc_b_axuser_0_reg[i] <= uc2rb_rd_req_desc_b_axuser_0_reg[i];
             else 
               rd_req_desc_b_axuser_0_reg[i] <= rd_req_desc_b_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_1_reg_we[i])
               rd_req_desc_b_axuser_1_reg[i] <= uc2rb_rd_req_desc_b_axuser_1_reg[i];
             else 
               rd_req_desc_b_axuser_1_reg[i] <= rd_req_desc_b_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_2_reg_we[i])
               rd_req_desc_b_axuser_2_reg[i] <= uc2rb_rd_req_desc_b_axuser_2_reg[i];
             else 
               rd_req_desc_b_axuser_2_reg[i] <= rd_req_desc_b_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_3_reg_we[i])
               rd_req_desc_b_axuser_3_reg[i] <= uc2rb_rd_req_desc_b_axuser_3_reg[i];
             else 
               rd_req_desc_b_axuser_3_reg[i] <= rd_req_desc_b_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_4_reg_we[i])
               rd_req_desc_b_axuser_4_reg[i] <= uc2rb_rd_req_desc_b_axuser_4_reg[i];
             else 
               rd_req_desc_b_axuser_4_reg[i] <= rd_req_desc_b_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_5_reg_we[i])
               rd_req_desc_b_axuser_5_reg[i] <= uc2rb_rd_req_desc_b_axuser_5_reg[i];
             else 
               rd_req_desc_b_axuser_5_reg[i] <= rd_req_desc_b_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_6_reg_we[i])
               rd_req_desc_b_axuser_6_reg[i] <= uc2rb_rd_req_desc_b_axuser_6_reg[i];
             else 
               rd_req_desc_b_axuser_6_reg[i] <= rd_req_desc_b_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_7_reg_we[i])
               rd_req_desc_b_axuser_7_reg[i] <= uc2rb_rd_req_desc_b_axuser_7_reg[i];
             else 
               rd_req_desc_b_axuser_7_reg[i] <= rd_req_desc_b_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_8_reg_we[i])
               rd_req_desc_b_axuser_8_reg[i] <= uc2rb_rd_req_desc_b_axuser_8_reg[i];
             else 
               rd_req_desc_b_axuser_8_reg[i] <= rd_req_desc_b_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_9_reg_we[i])
               rd_req_desc_b_axuser_9_reg[i] <= uc2rb_rd_req_desc_b_axuser_9_reg[i];
             else 
               rd_req_desc_b_axuser_9_reg[i] <= rd_req_desc_b_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_10_reg_we[i])
               rd_req_desc_b_axuser_10_reg[i] <= uc2rb_rd_req_desc_b_axuser_10_reg[i];
             else 
               rd_req_desc_b_axuser_10_reg[i] <= rd_req_desc_b_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_11_reg_we[i])
               rd_req_desc_b_axuser_11_reg[i] <= uc2rb_rd_req_desc_b_axuser_11_reg[i];
             else 
               rd_req_desc_b_axuser_11_reg[i] <= rd_req_desc_b_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_12_reg_we[i])
               rd_req_desc_b_axuser_12_reg[i] <= uc2rb_rd_req_desc_b_axuser_12_reg[i];
             else 
               rd_req_desc_b_axuser_12_reg[i] <= rd_req_desc_b_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_13_reg_we[i])
               rd_req_desc_b_axuser_13_reg[i] <= uc2rb_rd_req_desc_b_axuser_13_reg[i];
             else 
               rd_req_desc_b_axuser_13_reg[i] <= rd_req_desc_b_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_14_reg_we[i])
               rd_req_desc_b_axuser_14_reg[i] <= uc2rb_rd_req_desc_b_axuser_14_reg[i];
             else 
               rd_req_desc_b_axuser_14_reg[i] <= rd_req_desc_b_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_B_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_b_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_b_axuser_15_reg_we[i])
               rd_req_desc_b_axuser_15_reg[i] <= uc2rb_rd_req_desc_b_axuser_15_reg[i];
             else 
               rd_req_desc_b_axuser_15_reg[i] <= rd_req_desc_b_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_B_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_txn_type_reg_we[i])
               wr_req_desc_b_txn_type_reg[i] <= uc2rb_wr_req_desc_b_txn_type_reg[i];
             else 
               wr_req_desc_b_txn_type_reg[i] <= wr_req_desc_b_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_B_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_size_reg_we[i])
               wr_req_desc_b_size_reg[i] <= uc2rb_wr_req_desc_b_size_reg[i];
             else 
               wr_req_desc_b_size_reg[i] <= wr_req_desc_b_size_reg[i];
        end
     end
   //WR_REQ_DESC_B_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_data_offset_reg_we[i])
               wr_req_desc_b_data_offset_reg[i] <= uc2rb_wr_req_desc_b_data_offset_reg[i];
             else 
               wr_req_desc_b_data_offset_reg[i] <= wr_req_desc_b_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axsize_reg_we[i])
               wr_req_desc_b_axsize_reg[i] <= uc2rb_wr_req_desc_b_axsize_reg[i];
             else 
               wr_req_desc_b_axsize_reg[i] <= wr_req_desc_b_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_B_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_attr_reg_we[i])
               wr_req_desc_b_attr_reg[i] <= uc2rb_wr_req_desc_b_attr_reg[i];
             else 
               wr_req_desc_b_attr_reg[i] <= wr_req_desc_b_attr_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axaddr_0_reg_we[i])
               wr_req_desc_b_axaddr_0_reg[i] <= uc2rb_wr_req_desc_b_axaddr_0_reg[i];
             else 
               wr_req_desc_b_axaddr_0_reg[i] <= wr_req_desc_b_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axaddr_1_reg_we[i])
               wr_req_desc_b_axaddr_1_reg[i] <= uc2rb_wr_req_desc_b_axaddr_1_reg[i];
             else 
               wr_req_desc_b_axaddr_1_reg[i] <= wr_req_desc_b_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axaddr_2_reg_we[i])
               wr_req_desc_b_axaddr_2_reg[i] <= uc2rb_wr_req_desc_b_axaddr_2_reg[i];
             else 
               wr_req_desc_b_axaddr_2_reg[i] <= wr_req_desc_b_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axaddr_3_reg_we[i])
               wr_req_desc_b_axaddr_3_reg[i] <= uc2rb_wr_req_desc_b_axaddr_3_reg[i];
             else 
               wr_req_desc_b_axaddr_3_reg[i] <= wr_req_desc_b_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axid_0_reg_we[i])
               wr_req_desc_b_axid_0_reg[i] <= uc2rb_wr_req_desc_b_axid_0_reg[i];
             else 
               wr_req_desc_b_axid_0_reg[i] <= wr_req_desc_b_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axid_1_reg_we[i])
               wr_req_desc_b_axid_1_reg[i] <= uc2rb_wr_req_desc_b_axid_1_reg[i];
             else 
               wr_req_desc_b_axid_1_reg[i] <= wr_req_desc_b_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axid_2_reg_we[i])
               wr_req_desc_b_axid_2_reg[i] <= uc2rb_wr_req_desc_b_axid_2_reg[i];
             else 
               wr_req_desc_b_axid_2_reg[i] <= wr_req_desc_b_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axid_3_reg_we[i])
               wr_req_desc_b_axid_3_reg[i] <= uc2rb_wr_req_desc_b_axid_3_reg[i];
             else 
               wr_req_desc_b_axid_3_reg[i] <= wr_req_desc_b_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_0_reg_we[i])
               wr_req_desc_b_axuser_0_reg[i] <= uc2rb_wr_req_desc_b_axuser_0_reg[i];
             else 
               wr_req_desc_b_axuser_0_reg[i] <= wr_req_desc_b_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_1_reg_we[i])
               wr_req_desc_b_axuser_1_reg[i] <= uc2rb_wr_req_desc_b_axuser_1_reg[i];
             else 
               wr_req_desc_b_axuser_1_reg[i] <= wr_req_desc_b_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_2_reg_we[i])
               wr_req_desc_b_axuser_2_reg[i] <= uc2rb_wr_req_desc_b_axuser_2_reg[i];
             else 
               wr_req_desc_b_axuser_2_reg[i] <= wr_req_desc_b_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_3_reg_we[i])
               wr_req_desc_b_axuser_3_reg[i] <= uc2rb_wr_req_desc_b_axuser_3_reg[i];
             else 
               wr_req_desc_b_axuser_3_reg[i] <= wr_req_desc_b_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_4_reg_we[i])
               wr_req_desc_b_axuser_4_reg[i] <= uc2rb_wr_req_desc_b_axuser_4_reg[i];
             else 
               wr_req_desc_b_axuser_4_reg[i] <= wr_req_desc_b_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_5_reg_we[i])
               wr_req_desc_b_axuser_5_reg[i] <= uc2rb_wr_req_desc_b_axuser_5_reg[i];
             else 
               wr_req_desc_b_axuser_5_reg[i] <= wr_req_desc_b_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_6_reg_we[i])
               wr_req_desc_b_axuser_6_reg[i] <= uc2rb_wr_req_desc_b_axuser_6_reg[i];
             else 
               wr_req_desc_b_axuser_6_reg[i] <= wr_req_desc_b_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_7_reg_we[i])
               wr_req_desc_b_axuser_7_reg[i] <= uc2rb_wr_req_desc_b_axuser_7_reg[i];
             else 
               wr_req_desc_b_axuser_7_reg[i] <= wr_req_desc_b_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_8_reg_we[i])
               wr_req_desc_b_axuser_8_reg[i] <= uc2rb_wr_req_desc_b_axuser_8_reg[i];
             else 
               wr_req_desc_b_axuser_8_reg[i] <= wr_req_desc_b_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_9_reg_we[i])
               wr_req_desc_b_axuser_9_reg[i] <= uc2rb_wr_req_desc_b_axuser_9_reg[i];
             else 
               wr_req_desc_b_axuser_9_reg[i] <= wr_req_desc_b_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_10_reg_we[i])
               wr_req_desc_b_axuser_10_reg[i] <= uc2rb_wr_req_desc_b_axuser_10_reg[i];
             else 
               wr_req_desc_b_axuser_10_reg[i] <= wr_req_desc_b_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_11_reg_we[i])
               wr_req_desc_b_axuser_11_reg[i] <= uc2rb_wr_req_desc_b_axuser_11_reg[i];
             else 
               wr_req_desc_b_axuser_11_reg[i] <= wr_req_desc_b_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_12_reg_we[i])
               wr_req_desc_b_axuser_12_reg[i] <= uc2rb_wr_req_desc_b_axuser_12_reg[i];
             else 
               wr_req_desc_b_axuser_12_reg[i] <= wr_req_desc_b_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_13_reg_we[i])
               wr_req_desc_b_axuser_13_reg[i] <= uc2rb_wr_req_desc_b_axuser_13_reg[i];
             else 
               wr_req_desc_b_axuser_13_reg[i] <= wr_req_desc_b_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_14_reg_we[i])
               wr_req_desc_b_axuser_14_reg[i] <= uc2rb_wr_req_desc_b_axuser_14_reg[i];
             else 
               wr_req_desc_b_axuser_14_reg[i] <= wr_req_desc_b_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_B_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_axuser_15_reg_we[i])
               wr_req_desc_b_axuser_15_reg[i] <= uc2rb_wr_req_desc_b_axuser_15_reg[i];
             else 
               wr_req_desc_b_axuser_15_reg[i] <= wr_req_desc_b_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_0_reg_we[i])
               wr_req_desc_b_wuser_0_reg[i] <= uc2rb_wr_req_desc_b_wuser_0_reg[i];
             else 
               wr_req_desc_b_wuser_0_reg[i] <= wr_req_desc_b_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_1_reg_we[i])
               wr_req_desc_b_wuser_1_reg[i] <= uc2rb_wr_req_desc_b_wuser_1_reg[i];
             else 
               wr_req_desc_b_wuser_1_reg[i] <= wr_req_desc_b_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_2_reg_we[i])
               wr_req_desc_b_wuser_2_reg[i] <= uc2rb_wr_req_desc_b_wuser_2_reg[i];
             else 
               wr_req_desc_b_wuser_2_reg[i] <= wr_req_desc_b_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_3_reg_we[i])
               wr_req_desc_b_wuser_3_reg[i] <= uc2rb_wr_req_desc_b_wuser_3_reg[i];
             else 
               wr_req_desc_b_wuser_3_reg[i] <= wr_req_desc_b_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_4_reg_we[i])
               wr_req_desc_b_wuser_4_reg[i] <= uc2rb_wr_req_desc_b_wuser_4_reg[i];
             else 
               wr_req_desc_b_wuser_4_reg[i] <= wr_req_desc_b_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_5_reg_we[i])
               wr_req_desc_b_wuser_5_reg[i] <= uc2rb_wr_req_desc_b_wuser_5_reg[i];
             else 
               wr_req_desc_b_wuser_5_reg[i] <= wr_req_desc_b_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_6_reg_we[i])
               wr_req_desc_b_wuser_6_reg[i] <= uc2rb_wr_req_desc_b_wuser_6_reg[i];
             else 
               wr_req_desc_b_wuser_6_reg[i] <= wr_req_desc_b_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_7_reg_we[i])
               wr_req_desc_b_wuser_7_reg[i] <= uc2rb_wr_req_desc_b_wuser_7_reg[i];
             else 
               wr_req_desc_b_wuser_7_reg[i] <= wr_req_desc_b_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_8_reg_we[i])
               wr_req_desc_b_wuser_8_reg[i] <= uc2rb_wr_req_desc_b_wuser_8_reg[i];
             else 
               wr_req_desc_b_wuser_8_reg[i] <= wr_req_desc_b_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_9_reg_we[i])
               wr_req_desc_b_wuser_9_reg[i] <= uc2rb_wr_req_desc_b_wuser_9_reg[i];
             else 
               wr_req_desc_b_wuser_9_reg[i] <= wr_req_desc_b_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_10_reg_we[i])
               wr_req_desc_b_wuser_10_reg[i] <= uc2rb_wr_req_desc_b_wuser_10_reg[i];
             else 
               wr_req_desc_b_wuser_10_reg[i] <= wr_req_desc_b_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_11_reg_we[i])
               wr_req_desc_b_wuser_11_reg[i] <= uc2rb_wr_req_desc_b_wuser_11_reg[i];
             else 
               wr_req_desc_b_wuser_11_reg[i] <= wr_req_desc_b_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_12_reg_we[i])
               wr_req_desc_b_wuser_12_reg[i] <= uc2rb_wr_req_desc_b_wuser_12_reg[i];
             else 
               wr_req_desc_b_wuser_12_reg[i] <= wr_req_desc_b_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_13_reg_we[i])
               wr_req_desc_b_wuser_13_reg[i] <= uc2rb_wr_req_desc_b_wuser_13_reg[i];
             else 
               wr_req_desc_b_wuser_13_reg[i] <= wr_req_desc_b_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_14_reg_we[i])
               wr_req_desc_b_wuser_14_reg[i] <= uc2rb_wr_req_desc_b_wuser_14_reg[i];
             else 
               wr_req_desc_b_wuser_14_reg[i] <= wr_req_desc_b_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_B_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_b_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_b_wuser_15_reg_we[i])
               wr_req_desc_b_wuser_15_reg[i] <= uc2rb_wr_req_desc_b_wuser_15_reg[i];
             else 
               wr_req_desc_b_wuser_15_reg[i] <= wr_req_desc_b_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_B_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_b_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_b_resp_reg_we[i])
               sn_resp_desc_b_resp_reg[i] <= uc2rb_sn_resp_desc_b_resp_reg[i];
             else 
               sn_resp_desc_b_resp_reg[i] <= sn_resp_desc_b_resp_reg[i];
        end
     end
   //RD_REQ_DESC_C_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_txn_type_reg_we[i])
               rd_req_desc_c_txn_type_reg[i] <= uc2rb_rd_req_desc_c_txn_type_reg[i];
             else 
               rd_req_desc_c_txn_type_reg[i] <= rd_req_desc_c_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_C_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_size_reg_we[i])
               rd_req_desc_c_size_reg[i] <= uc2rb_rd_req_desc_c_size_reg[i];
             else 
               rd_req_desc_c_size_reg[i] <= rd_req_desc_c_size_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axsize_reg_we[i])
               rd_req_desc_c_axsize_reg[i] <= uc2rb_rd_req_desc_c_axsize_reg[i];
             else 
               rd_req_desc_c_axsize_reg[i] <= rd_req_desc_c_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_C_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_attr_reg_we[i])
               rd_req_desc_c_attr_reg[i] <= uc2rb_rd_req_desc_c_attr_reg[i];
             else 
               rd_req_desc_c_attr_reg[i] <= rd_req_desc_c_attr_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axaddr_0_reg_we[i])
               rd_req_desc_c_axaddr_0_reg[i] <= uc2rb_rd_req_desc_c_axaddr_0_reg[i];
             else 
               rd_req_desc_c_axaddr_0_reg[i] <= rd_req_desc_c_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axaddr_1_reg_we[i])
               rd_req_desc_c_axaddr_1_reg[i] <= uc2rb_rd_req_desc_c_axaddr_1_reg[i];
             else 
               rd_req_desc_c_axaddr_1_reg[i] <= rd_req_desc_c_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axaddr_2_reg_we[i])
               rd_req_desc_c_axaddr_2_reg[i] <= uc2rb_rd_req_desc_c_axaddr_2_reg[i];
             else 
               rd_req_desc_c_axaddr_2_reg[i] <= rd_req_desc_c_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axaddr_3_reg_we[i])
               rd_req_desc_c_axaddr_3_reg[i] <= uc2rb_rd_req_desc_c_axaddr_3_reg[i];
             else 
               rd_req_desc_c_axaddr_3_reg[i] <= rd_req_desc_c_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axid_0_reg_we[i])
               rd_req_desc_c_axid_0_reg[i] <= uc2rb_rd_req_desc_c_axid_0_reg[i];
             else 
               rd_req_desc_c_axid_0_reg[i] <= rd_req_desc_c_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axid_1_reg_we[i])
               rd_req_desc_c_axid_1_reg[i] <= uc2rb_rd_req_desc_c_axid_1_reg[i];
             else 
               rd_req_desc_c_axid_1_reg[i] <= rd_req_desc_c_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axid_2_reg_we[i])
               rd_req_desc_c_axid_2_reg[i] <= uc2rb_rd_req_desc_c_axid_2_reg[i];
             else 
               rd_req_desc_c_axid_2_reg[i] <= rd_req_desc_c_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axid_3_reg_we[i])
               rd_req_desc_c_axid_3_reg[i] <= uc2rb_rd_req_desc_c_axid_3_reg[i];
             else 
               rd_req_desc_c_axid_3_reg[i] <= rd_req_desc_c_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_0_reg_we[i])
               rd_req_desc_c_axuser_0_reg[i] <= uc2rb_rd_req_desc_c_axuser_0_reg[i];
             else 
               rd_req_desc_c_axuser_0_reg[i] <= rd_req_desc_c_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_1_reg_we[i])
               rd_req_desc_c_axuser_1_reg[i] <= uc2rb_rd_req_desc_c_axuser_1_reg[i];
             else 
               rd_req_desc_c_axuser_1_reg[i] <= rd_req_desc_c_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_2_reg_we[i])
               rd_req_desc_c_axuser_2_reg[i] <= uc2rb_rd_req_desc_c_axuser_2_reg[i];
             else 
               rd_req_desc_c_axuser_2_reg[i] <= rd_req_desc_c_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_3_reg_we[i])
               rd_req_desc_c_axuser_3_reg[i] <= uc2rb_rd_req_desc_c_axuser_3_reg[i];
             else 
               rd_req_desc_c_axuser_3_reg[i] <= rd_req_desc_c_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_4_reg_we[i])
               rd_req_desc_c_axuser_4_reg[i] <= uc2rb_rd_req_desc_c_axuser_4_reg[i];
             else 
               rd_req_desc_c_axuser_4_reg[i] <= rd_req_desc_c_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_5_reg_we[i])
               rd_req_desc_c_axuser_5_reg[i] <= uc2rb_rd_req_desc_c_axuser_5_reg[i];
             else 
               rd_req_desc_c_axuser_5_reg[i] <= rd_req_desc_c_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_6_reg_we[i])
               rd_req_desc_c_axuser_6_reg[i] <= uc2rb_rd_req_desc_c_axuser_6_reg[i];
             else 
               rd_req_desc_c_axuser_6_reg[i] <= rd_req_desc_c_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_7_reg_we[i])
               rd_req_desc_c_axuser_7_reg[i] <= uc2rb_rd_req_desc_c_axuser_7_reg[i];
             else 
               rd_req_desc_c_axuser_7_reg[i] <= rd_req_desc_c_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_8_reg_we[i])
               rd_req_desc_c_axuser_8_reg[i] <= uc2rb_rd_req_desc_c_axuser_8_reg[i];
             else 
               rd_req_desc_c_axuser_8_reg[i] <= rd_req_desc_c_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_9_reg_we[i])
               rd_req_desc_c_axuser_9_reg[i] <= uc2rb_rd_req_desc_c_axuser_9_reg[i];
             else 
               rd_req_desc_c_axuser_9_reg[i] <= rd_req_desc_c_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_10_reg_we[i])
               rd_req_desc_c_axuser_10_reg[i] <= uc2rb_rd_req_desc_c_axuser_10_reg[i];
             else 
               rd_req_desc_c_axuser_10_reg[i] <= rd_req_desc_c_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_11_reg_we[i])
               rd_req_desc_c_axuser_11_reg[i] <= uc2rb_rd_req_desc_c_axuser_11_reg[i];
             else 
               rd_req_desc_c_axuser_11_reg[i] <= rd_req_desc_c_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_12_reg_we[i])
               rd_req_desc_c_axuser_12_reg[i] <= uc2rb_rd_req_desc_c_axuser_12_reg[i];
             else 
               rd_req_desc_c_axuser_12_reg[i] <= rd_req_desc_c_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_13_reg_we[i])
               rd_req_desc_c_axuser_13_reg[i] <= uc2rb_rd_req_desc_c_axuser_13_reg[i];
             else 
               rd_req_desc_c_axuser_13_reg[i] <= rd_req_desc_c_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_14_reg_we[i])
               rd_req_desc_c_axuser_14_reg[i] <= uc2rb_rd_req_desc_c_axuser_14_reg[i];
             else 
               rd_req_desc_c_axuser_14_reg[i] <= rd_req_desc_c_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_C_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_c_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_c_axuser_15_reg_we[i])
               rd_req_desc_c_axuser_15_reg[i] <= uc2rb_rd_req_desc_c_axuser_15_reg[i];
             else 
               rd_req_desc_c_axuser_15_reg[i] <= rd_req_desc_c_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_C_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_txn_type_reg_we[i])
               wr_req_desc_c_txn_type_reg[i] <= uc2rb_wr_req_desc_c_txn_type_reg[i];
             else 
               wr_req_desc_c_txn_type_reg[i] <= wr_req_desc_c_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_C_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_size_reg_we[i])
               wr_req_desc_c_size_reg[i] <= uc2rb_wr_req_desc_c_size_reg[i];
             else 
               wr_req_desc_c_size_reg[i] <= wr_req_desc_c_size_reg[i];
        end
     end
   //WR_REQ_DESC_C_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_data_offset_reg_we[i])
               wr_req_desc_c_data_offset_reg[i] <= uc2rb_wr_req_desc_c_data_offset_reg[i];
             else 
               wr_req_desc_c_data_offset_reg[i] <= wr_req_desc_c_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axsize_reg_we[i])
               wr_req_desc_c_axsize_reg[i] <= uc2rb_wr_req_desc_c_axsize_reg[i];
             else 
               wr_req_desc_c_axsize_reg[i] <= wr_req_desc_c_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_C_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_attr_reg_we[i])
               wr_req_desc_c_attr_reg[i] <= uc2rb_wr_req_desc_c_attr_reg[i];
             else 
               wr_req_desc_c_attr_reg[i] <= wr_req_desc_c_attr_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axaddr_0_reg_we[i])
               wr_req_desc_c_axaddr_0_reg[i] <= uc2rb_wr_req_desc_c_axaddr_0_reg[i];
             else 
               wr_req_desc_c_axaddr_0_reg[i] <= wr_req_desc_c_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axaddr_1_reg_we[i])
               wr_req_desc_c_axaddr_1_reg[i] <= uc2rb_wr_req_desc_c_axaddr_1_reg[i];
             else 
               wr_req_desc_c_axaddr_1_reg[i] <= wr_req_desc_c_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axaddr_2_reg_we[i])
               wr_req_desc_c_axaddr_2_reg[i] <= uc2rb_wr_req_desc_c_axaddr_2_reg[i];
             else 
               wr_req_desc_c_axaddr_2_reg[i] <= wr_req_desc_c_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axaddr_3_reg_we[i])
               wr_req_desc_c_axaddr_3_reg[i] <= uc2rb_wr_req_desc_c_axaddr_3_reg[i];
             else 
               wr_req_desc_c_axaddr_3_reg[i] <= wr_req_desc_c_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axid_0_reg_we[i])
               wr_req_desc_c_axid_0_reg[i] <= uc2rb_wr_req_desc_c_axid_0_reg[i];
             else 
               wr_req_desc_c_axid_0_reg[i] <= wr_req_desc_c_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axid_1_reg_we[i])
               wr_req_desc_c_axid_1_reg[i] <= uc2rb_wr_req_desc_c_axid_1_reg[i];
             else 
               wr_req_desc_c_axid_1_reg[i] <= wr_req_desc_c_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axid_2_reg_we[i])
               wr_req_desc_c_axid_2_reg[i] <= uc2rb_wr_req_desc_c_axid_2_reg[i];
             else 
               wr_req_desc_c_axid_2_reg[i] <= wr_req_desc_c_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axid_3_reg_we[i])
               wr_req_desc_c_axid_3_reg[i] <= uc2rb_wr_req_desc_c_axid_3_reg[i];
             else 
               wr_req_desc_c_axid_3_reg[i] <= wr_req_desc_c_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_0_reg_we[i])
               wr_req_desc_c_axuser_0_reg[i] <= uc2rb_wr_req_desc_c_axuser_0_reg[i];
             else 
               wr_req_desc_c_axuser_0_reg[i] <= wr_req_desc_c_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_1_reg_we[i])
               wr_req_desc_c_axuser_1_reg[i] <= uc2rb_wr_req_desc_c_axuser_1_reg[i];
             else 
               wr_req_desc_c_axuser_1_reg[i] <= wr_req_desc_c_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_2_reg_we[i])
               wr_req_desc_c_axuser_2_reg[i] <= uc2rb_wr_req_desc_c_axuser_2_reg[i];
             else 
               wr_req_desc_c_axuser_2_reg[i] <= wr_req_desc_c_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_3_reg_we[i])
               wr_req_desc_c_axuser_3_reg[i] <= uc2rb_wr_req_desc_c_axuser_3_reg[i];
             else 
               wr_req_desc_c_axuser_3_reg[i] <= wr_req_desc_c_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_4_reg_we[i])
               wr_req_desc_c_axuser_4_reg[i] <= uc2rb_wr_req_desc_c_axuser_4_reg[i];
             else 
               wr_req_desc_c_axuser_4_reg[i] <= wr_req_desc_c_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_5_reg_we[i])
               wr_req_desc_c_axuser_5_reg[i] <= uc2rb_wr_req_desc_c_axuser_5_reg[i];
             else 
               wr_req_desc_c_axuser_5_reg[i] <= wr_req_desc_c_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_6_reg_we[i])
               wr_req_desc_c_axuser_6_reg[i] <= uc2rb_wr_req_desc_c_axuser_6_reg[i];
             else 
               wr_req_desc_c_axuser_6_reg[i] <= wr_req_desc_c_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_7_reg_we[i])
               wr_req_desc_c_axuser_7_reg[i] <= uc2rb_wr_req_desc_c_axuser_7_reg[i];
             else 
               wr_req_desc_c_axuser_7_reg[i] <= wr_req_desc_c_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_8_reg_we[i])
               wr_req_desc_c_axuser_8_reg[i] <= uc2rb_wr_req_desc_c_axuser_8_reg[i];
             else 
               wr_req_desc_c_axuser_8_reg[i] <= wr_req_desc_c_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_9_reg_we[i])
               wr_req_desc_c_axuser_9_reg[i] <= uc2rb_wr_req_desc_c_axuser_9_reg[i];
             else 
               wr_req_desc_c_axuser_9_reg[i] <= wr_req_desc_c_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_10_reg_we[i])
               wr_req_desc_c_axuser_10_reg[i] <= uc2rb_wr_req_desc_c_axuser_10_reg[i];
             else 
               wr_req_desc_c_axuser_10_reg[i] <= wr_req_desc_c_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_11_reg_we[i])
               wr_req_desc_c_axuser_11_reg[i] <= uc2rb_wr_req_desc_c_axuser_11_reg[i];
             else 
               wr_req_desc_c_axuser_11_reg[i] <= wr_req_desc_c_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_12_reg_we[i])
               wr_req_desc_c_axuser_12_reg[i] <= uc2rb_wr_req_desc_c_axuser_12_reg[i];
             else 
               wr_req_desc_c_axuser_12_reg[i] <= wr_req_desc_c_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_13_reg_we[i])
               wr_req_desc_c_axuser_13_reg[i] <= uc2rb_wr_req_desc_c_axuser_13_reg[i];
             else 
               wr_req_desc_c_axuser_13_reg[i] <= wr_req_desc_c_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_14_reg_we[i])
               wr_req_desc_c_axuser_14_reg[i] <= uc2rb_wr_req_desc_c_axuser_14_reg[i];
             else 
               wr_req_desc_c_axuser_14_reg[i] <= wr_req_desc_c_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_C_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_axuser_15_reg_we[i])
               wr_req_desc_c_axuser_15_reg[i] <= uc2rb_wr_req_desc_c_axuser_15_reg[i];
             else 
               wr_req_desc_c_axuser_15_reg[i] <= wr_req_desc_c_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_0_reg_we[i])
               wr_req_desc_c_wuser_0_reg[i] <= uc2rb_wr_req_desc_c_wuser_0_reg[i];
             else 
               wr_req_desc_c_wuser_0_reg[i] <= wr_req_desc_c_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_1_reg_we[i])
               wr_req_desc_c_wuser_1_reg[i] <= uc2rb_wr_req_desc_c_wuser_1_reg[i];
             else 
               wr_req_desc_c_wuser_1_reg[i] <= wr_req_desc_c_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_2_reg_we[i])
               wr_req_desc_c_wuser_2_reg[i] <= uc2rb_wr_req_desc_c_wuser_2_reg[i];
             else 
               wr_req_desc_c_wuser_2_reg[i] <= wr_req_desc_c_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_3_reg_we[i])
               wr_req_desc_c_wuser_3_reg[i] <= uc2rb_wr_req_desc_c_wuser_3_reg[i];
             else 
               wr_req_desc_c_wuser_3_reg[i] <= wr_req_desc_c_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_4_reg_we[i])
               wr_req_desc_c_wuser_4_reg[i] <= uc2rb_wr_req_desc_c_wuser_4_reg[i];
             else 
               wr_req_desc_c_wuser_4_reg[i] <= wr_req_desc_c_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_5_reg_we[i])
               wr_req_desc_c_wuser_5_reg[i] <= uc2rb_wr_req_desc_c_wuser_5_reg[i];
             else 
               wr_req_desc_c_wuser_5_reg[i] <= wr_req_desc_c_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_6_reg_we[i])
               wr_req_desc_c_wuser_6_reg[i] <= uc2rb_wr_req_desc_c_wuser_6_reg[i];
             else 
               wr_req_desc_c_wuser_6_reg[i] <= wr_req_desc_c_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_7_reg_we[i])
               wr_req_desc_c_wuser_7_reg[i] <= uc2rb_wr_req_desc_c_wuser_7_reg[i];
             else 
               wr_req_desc_c_wuser_7_reg[i] <= wr_req_desc_c_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_8_reg_we[i])
               wr_req_desc_c_wuser_8_reg[i] <= uc2rb_wr_req_desc_c_wuser_8_reg[i];
             else 
               wr_req_desc_c_wuser_8_reg[i] <= wr_req_desc_c_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_9_reg_we[i])
               wr_req_desc_c_wuser_9_reg[i] <= uc2rb_wr_req_desc_c_wuser_9_reg[i];
             else 
               wr_req_desc_c_wuser_9_reg[i] <= wr_req_desc_c_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_10_reg_we[i])
               wr_req_desc_c_wuser_10_reg[i] <= uc2rb_wr_req_desc_c_wuser_10_reg[i];
             else 
               wr_req_desc_c_wuser_10_reg[i] <= wr_req_desc_c_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_11_reg_we[i])
               wr_req_desc_c_wuser_11_reg[i] <= uc2rb_wr_req_desc_c_wuser_11_reg[i];
             else 
               wr_req_desc_c_wuser_11_reg[i] <= wr_req_desc_c_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_12_reg_we[i])
               wr_req_desc_c_wuser_12_reg[i] <= uc2rb_wr_req_desc_c_wuser_12_reg[i];
             else 
               wr_req_desc_c_wuser_12_reg[i] <= wr_req_desc_c_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_13_reg_we[i])
               wr_req_desc_c_wuser_13_reg[i] <= uc2rb_wr_req_desc_c_wuser_13_reg[i];
             else 
               wr_req_desc_c_wuser_13_reg[i] <= wr_req_desc_c_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_14_reg_we[i])
               wr_req_desc_c_wuser_14_reg[i] <= uc2rb_wr_req_desc_c_wuser_14_reg[i];
             else 
               wr_req_desc_c_wuser_14_reg[i] <= wr_req_desc_c_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_C_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_c_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_c_wuser_15_reg_we[i])
               wr_req_desc_c_wuser_15_reg[i] <= uc2rb_wr_req_desc_c_wuser_15_reg[i];
             else 
               wr_req_desc_c_wuser_15_reg[i] <= wr_req_desc_c_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_C_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_c_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_c_resp_reg_we[i])
               sn_resp_desc_c_resp_reg[i] <= uc2rb_sn_resp_desc_c_resp_reg[i];
             else 
               sn_resp_desc_c_resp_reg[i] <= sn_resp_desc_c_resp_reg[i];
        end
     end
   //RD_REQ_DESC_D_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_txn_type_reg_we[i])
               rd_req_desc_d_txn_type_reg[i] <= uc2rb_rd_req_desc_d_txn_type_reg[i];
             else 
               rd_req_desc_d_txn_type_reg[i] <= rd_req_desc_d_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_D_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_size_reg_we[i])
               rd_req_desc_d_size_reg[i] <= uc2rb_rd_req_desc_d_size_reg[i];
             else 
               rd_req_desc_d_size_reg[i] <= rd_req_desc_d_size_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axsize_reg_we[i])
               rd_req_desc_d_axsize_reg[i] <= uc2rb_rd_req_desc_d_axsize_reg[i];
             else 
               rd_req_desc_d_axsize_reg[i] <= rd_req_desc_d_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_D_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_attr_reg_we[i])
               rd_req_desc_d_attr_reg[i] <= uc2rb_rd_req_desc_d_attr_reg[i];
             else 
               rd_req_desc_d_attr_reg[i] <= rd_req_desc_d_attr_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axaddr_0_reg_we[i])
               rd_req_desc_d_axaddr_0_reg[i] <= uc2rb_rd_req_desc_d_axaddr_0_reg[i];
             else 
               rd_req_desc_d_axaddr_0_reg[i] <= rd_req_desc_d_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axaddr_1_reg_we[i])
               rd_req_desc_d_axaddr_1_reg[i] <= uc2rb_rd_req_desc_d_axaddr_1_reg[i];
             else 
               rd_req_desc_d_axaddr_1_reg[i] <= rd_req_desc_d_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axaddr_2_reg_we[i])
               rd_req_desc_d_axaddr_2_reg[i] <= uc2rb_rd_req_desc_d_axaddr_2_reg[i];
             else 
               rd_req_desc_d_axaddr_2_reg[i] <= rd_req_desc_d_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axaddr_3_reg_we[i])
               rd_req_desc_d_axaddr_3_reg[i] <= uc2rb_rd_req_desc_d_axaddr_3_reg[i];
             else 
               rd_req_desc_d_axaddr_3_reg[i] <= rd_req_desc_d_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axid_0_reg_we[i])
               rd_req_desc_d_axid_0_reg[i] <= uc2rb_rd_req_desc_d_axid_0_reg[i];
             else 
               rd_req_desc_d_axid_0_reg[i] <= rd_req_desc_d_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axid_1_reg_we[i])
               rd_req_desc_d_axid_1_reg[i] <= uc2rb_rd_req_desc_d_axid_1_reg[i];
             else 
               rd_req_desc_d_axid_1_reg[i] <= rd_req_desc_d_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axid_2_reg_we[i])
               rd_req_desc_d_axid_2_reg[i] <= uc2rb_rd_req_desc_d_axid_2_reg[i];
             else 
               rd_req_desc_d_axid_2_reg[i] <= rd_req_desc_d_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axid_3_reg_we[i])
               rd_req_desc_d_axid_3_reg[i] <= uc2rb_rd_req_desc_d_axid_3_reg[i];
             else 
               rd_req_desc_d_axid_3_reg[i] <= rd_req_desc_d_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_0_reg_we[i])
               rd_req_desc_d_axuser_0_reg[i] <= uc2rb_rd_req_desc_d_axuser_0_reg[i];
             else 
               rd_req_desc_d_axuser_0_reg[i] <= rd_req_desc_d_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_1_reg_we[i])
               rd_req_desc_d_axuser_1_reg[i] <= uc2rb_rd_req_desc_d_axuser_1_reg[i];
             else 
               rd_req_desc_d_axuser_1_reg[i] <= rd_req_desc_d_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_2_reg_we[i])
               rd_req_desc_d_axuser_2_reg[i] <= uc2rb_rd_req_desc_d_axuser_2_reg[i];
             else 
               rd_req_desc_d_axuser_2_reg[i] <= rd_req_desc_d_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_3_reg_we[i])
               rd_req_desc_d_axuser_3_reg[i] <= uc2rb_rd_req_desc_d_axuser_3_reg[i];
             else 
               rd_req_desc_d_axuser_3_reg[i] <= rd_req_desc_d_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_4_reg_we[i])
               rd_req_desc_d_axuser_4_reg[i] <= uc2rb_rd_req_desc_d_axuser_4_reg[i];
             else 
               rd_req_desc_d_axuser_4_reg[i] <= rd_req_desc_d_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_5_reg_we[i])
               rd_req_desc_d_axuser_5_reg[i] <= uc2rb_rd_req_desc_d_axuser_5_reg[i];
             else 
               rd_req_desc_d_axuser_5_reg[i] <= rd_req_desc_d_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_6_reg_we[i])
               rd_req_desc_d_axuser_6_reg[i] <= uc2rb_rd_req_desc_d_axuser_6_reg[i];
             else 
               rd_req_desc_d_axuser_6_reg[i] <= rd_req_desc_d_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_7_reg_we[i])
               rd_req_desc_d_axuser_7_reg[i] <= uc2rb_rd_req_desc_d_axuser_7_reg[i];
             else 
               rd_req_desc_d_axuser_7_reg[i] <= rd_req_desc_d_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_8_reg_we[i])
               rd_req_desc_d_axuser_8_reg[i] <= uc2rb_rd_req_desc_d_axuser_8_reg[i];
             else 
               rd_req_desc_d_axuser_8_reg[i] <= rd_req_desc_d_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_9_reg_we[i])
               rd_req_desc_d_axuser_9_reg[i] <= uc2rb_rd_req_desc_d_axuser_9_reg[i];
             else 
               rd_req_desc_d_axuser_9_reg[i] <= rd_req_desc_d_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_10_reg_we[i])
               rd_req_desc_d_axuser_10_reg[i] <= uc2rb_rd_req_desc_d_axuser_10_reg[i];
             else 
               rd_req_desc_d_axuser_10_reg[i] <= rd_req_desc_d_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_11_reg_we[i])
               rd_req_desc_d_axuser_11_reg[i] <= uc2rb_rd_req_desc_d_axuser_11_reg[i];
             else 
               rd_req_desc_d_axuser_11_reg[i] <= rd_req_desc_d_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_12_reg_we[i])
               rd_req_desc_d_axuser_12_reg[i] <= uc2rb_rd_req_desc_d_axuser_12_reg[i];
             else 
               rd_req_desc_d_axuser_12_reg[i] <= rd_req_desc_d_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_13_reg_we[i])
               rd_req_desc_d_axuser_13_reg[i] <= uc2rb_rd_req_desc_d_axuser_13_reg[i];
             else 
               rd_req_desc_d_axuser_13_reg[i] <= rd_req_desc_d_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_14_reg_we[i])
               rd_req_desc_d_axuser_14_reg[i] <= uc2rb_rd_req_desc_d_axuser_14_reg[i];
             else 
               rd_req_desc_d_axuser_14_reg[i] <= rd_req_desc_d_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_D_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_d_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_d_axuser_15_reg_we[i])
               rd_req_desc_d_axuser_15_reg[i] <= uc2rb_rd_req_desc_d_axuser_15_reg[i];
             else 
               rd_req_desc_d_axuser_15_reg[i] <= rd_req_desc_d_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_D_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_txn_type_reg_we[i])
               wr_req_desc_d_txn_type_reg[i] <= uc2rb_wr_req_desc_d_txn_type_reg[i];
             else 
               wr_req_desc_d_txn_type_reg[i] <= wr_req_desc_d_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_D_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_size_reg_we[i])
               wr_req_desc_d_size_reg[i] <= uc2rb_wr_req_desc_d_size_reg[i];
             else 
               wr_req_desc_d_size_reg[i] <= wr_req_desc_d_size_reg[i];
        end
     end
   //WR_REQ_DESC_D_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_data_offset_reg_we[i])
               wr_req_desc_d_data_offset_reg[i] <= uc2rb_wr_req_desc_d_data_offset_reg[i];
             else 
               wr_req_desc_d_data_offset_reg[i] <= wr_req_desc_d_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axsize_reg_we[i])
               wr_req_desc_d_axsize_reg[i] <= uc2rb_wr_req_desc_d_axsize_reg[i];
             else 
               wr_req_desc_d_axsize_reg[i] <= wr_req_desc_d_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_D_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_attr_reg_we[i])
               wr_req_desc_d_attr_reg[i] <= uc2rb_wr_req_desc_d_attr_reg[i];
             else 
               wr_req_desc_d_attr_reg[i] <= wr_req_desc_d_attr_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axaddr_0_reg_we[i])
               wr_req_desc_d_axaddr_0_reg[i] <= uc2rb_wr_req_desc_d_axaddr_0_reg[i];
             else 
               wr_req_desc_d_axaddr_0_reg[i] <= wr_req_desc_d_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axaddr_1_reg_we[i])
               wr_req_desc_d_axaddr_1_reg[i] <= uc2rb_wr_req_desc_d_axaddr_1_reg[i];
             else 
               wr_req_desc_d_axaddr_1_reg[i] <= wr_req_desc_d_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axaddr_2_reg_we[i])
               wr_req_desc_d_axaddr_2_reg[i] <= uc2rb_wr_req_desc_d_axaddr_2_reg[i];
             else 
               wr_req_desc_d_axaddr_2_reg[i] <= wr_req_desc_d_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axaddr_3_reg_we[i])
               wr_req_desc_d_axaddr_3_reg[i] <= uc2rb_wr_req_desc_d_axaddr_3_reg[i];
             else 
               wr_req_desc_d_axaddr_3_reg[i] <= wr_req_desc_d_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axid_0_reg_we[i])
               wr_req_desc_d_axid_0_reg[i] <= uc2rb_wr_req_desc_d_axid_0_reg[i];
             else 
               wr_req_desc_d_axid_0_reg[i] <= wr_req_desc_d_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axid_1_reg_we[i])
               wr_req_desc_d_axid_1_reg[i] <= uc2rb_wr_req_desc_d_axid_1_reg[i];
             else 
               wr_req_desc_d_axid_1_reg[i] <= wr_req_desc_d_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axid_2_reg_we[i])
               wr_req_desc_d_axid_2_reg[i] <= uc2rb_wr_req_desc_d_axid_2_reg[i];
             else 
               wr_req_desc_d_axid_2_reg[i] <= wr_req_desc_d_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axid_3_reg_we[i])
               wr_req_desc_d_axid_3_reg[i] <= uc2rb_wr_req_desc_d_axid_3_reg[i];
             else 
               wr_req_desc_d_axid_3_reg[i] <= wr_req_desc_d_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_0_reg_we[i])
               wr_req_desc_d_axuser_0_reg[i] <= uc2rb_wr_req_desc_d_axuser_0_reg[i];
             else 
               wr_req_desc_d_axuser_0_reg[i] <= wr_req_desc_d_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_1_reg_we[i])
               wr_req_desc_d_axuser_1_reg[i] <= uc2rb_wr_req_desc_d_axuser_1_reg[i];
             else 
               wr_req_desc_d_axuser_1_reg[i] <= wr_req_desc_d_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_2_reg_we[i])
               wr_req_desc_d_axuser_2_reg[i] <= uc2rb_wr_req_desc_d_axuser_2_reg[i];
             else 
               wr_req_desc_d_axuser_2_reg[i] <= wr_req_desc_d_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_3_reg_we[i])
               wr_req_desc_d_axuser_3_reg[i] <= uc2rb_wr_req_desc_d_axuser_3_reg[i];
             else 
               wr_req_desc_d_axuser_3_reg[i] <= wr_req_desc_d_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_4_reg_we[i])
               wr_req_desc_d_axuser_4_reg[i] <= uc2rb_wr_req_desc_d_axuser_4_reg[i];
             else 
               wr_req_desc_d_axuser_4_reg[i] <= wr_req_desc_d_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_5_reg_we[i])
               wr_req_desc_d_axuser_5_reg[i] <= uc2rb_wr_req_desc_d_axuser_5_reg[i];
             else 
               wr_req_desc_d_axuser_5_reg[i] <= wr_req_desc_d_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_6_reg_we[i])
               wr_req_desc_d_axuser_6_reg[i] <= uc2rb_wr_req_desc_d_axuser_6_reg[i];
             else 
               wr_req_desc_d_axuser_6_reg[i] <= wr_req_desc_d_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_7_reg_we[i])
               wr_req_desc_d_axuser_7_reg[i] <= uc2rb_wr_req_desc_d_axuser_7_reg[i];
             else 
               wr_req_desc_d_axuser_7_reg[i] <= wr_req_desc_d_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_8_reg_we[i])
               wr_req_desc_d_axuser_8_reg[i] <= uc2rb_wr_req_desc_d_axuser_8_reg[i];
             else 
               wr_req_desc_d_axuser_8_reg[i] <= wr_req_desc_d_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_9_reg_we[i])
               wr_req_desc_d_axuser_9_reg[i] <= uc2rb_wr_req_desc_d_axuser_9_reg[i];
             else 
               wr_req_desc_d_axuser_9_reg[i] <= wr_req_desc_d_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_10_reg_we[i])
               wr_req_desc_d_axuser_10_reg[i] <= uc2rb_wr_req_desc_d_axuser_10_reg[i];
             else 
               wr_req_desc_d_axuser_10_reg[i] <= wr_req_desc_d_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_11_reg_we[i])
               wr_req_desc_d_axuser_11_reg[i] <= uc2rb_wr_req_desc_d_axuser_11_reg[i];
             else 
               wr_req_desc_d_axuser_11_reg[i] <= wr_req_desc_d_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_12_reg_we[i])
               wr_req_desc_d_axuser_12_reg[i] <= uc2rb_wr_req_desc_d_axuser_12_reg[i];
             else 
               wr_req_desc_d_axuser_12_reg[i] <= wr_req_desc_d_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_13_reg_we[i])
               wr_req_desc_d_axuser_13_reg[i] <= uc2rb_wr_req_desc_d_axuser_13_reg[i];
             else 
               wr_req_desc_d_axuser_13_reg[i] <= wr_req_desc_d_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_14_reg_we[i])
               wr_req_desc_d_axuser_14_reg[i] <= uc2rb_wr_req_desc_d_axuser_14_reg[i];
             else 
               wr_req_desc_d_axuser_14_reg[i] <= wr_req_desc_d_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_D_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_axuser_15_reg_we[i])
               wr_req_desc_d_axuser_15_reg[i] <= uc2rb_wr_req_desc_d_axuser_15_reg[i];
             else 
               wr_req_desc_d_axuser_15_reg[i] <= wr_req_desc_d_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_0_reg_we[i])
               wr_req_desc_d_wuser_0_reg[i] <= uc2rb_wr_req_desc_d_wuser_0_reg[i];
             else 
               wr_req_desc_d_wuser_0_reg[i] <= wr_req_desc_d_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_1_reg_we[i])
               wr_req_desc_d_wuser_1_reg[i] <= uc2rb_wr_req_desc_d_wuser_1_reg[i];
             else 
               wr_req_desc_d_wuser_1_reg[i] <= wr_req_desc_d_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_2_reg_we[i])
               wr_req_desc_d_wuser_2_reg[i] <= uc2rb_wr_req_desc_d_wuser_2_reg[i];
             else 
               wr_req_desc_d_wuser_2_reg[i] <= wr_req_desc_d_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_3_reg_we[i])
               wr_req_desc_d_wuser_3_reg[i] <= uc2rb_wr_req_desc_d_wuser_3_reg[i];
             else 
               wr_req_desc_d_wuser_3_reg[i] <= wr_req_desc_d_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_4_reg_we[i])
               wr_req_desc_d_wuser_4_reg[i] <= uc2rb_wr_req_desc_d_wuser_4_reg[i];
             else 
               wr_req_desc_d_wuser_4_reg[i] <= wr_req_desc_d_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_5_reg_we[i])
               wr_req_desc_d_wuser_5_reg[i] <= uc2rb_wr_req_desc_d_wuser_5_reg[i];
             else 
               wr_req_desc_d_wuser_5_reg[i] <= wr_req_desc_d_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_6_reg_we[i])
               wr_req_desc_d_wuser_6_reg[i] <= uc2rb_wr_req_desc_d_wuser_6_reg[i];
             else 
               wr_req_desc_d_wuser_6_reg[i] <= wr_req_desc_d_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_7_reg_we[i])
               wr_req_desc_d_wuser_7_reg[i] <= uc2rb_wr_req_desc_d_wuser_7_reg[i];
             else 
               wr_req_desc_d_wuser_7_reg[i] <= wr_req_desc_d_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_8_reg_we[i])
               wr_req_desc_d_wuser_8_reg[i] <= uc2rb_wr_req_desc_d_wuser_8_reg[i];
             else 
               wr_req_desc_d_wuser_8_reg[i] <= wr_req_desc_d_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_9_reg_we[i])
               wr_req_desc_d_wuser_9_reg[i] <= uc2rb_wr_req_desc_d_wuser_9_reg[i];
             else 
               wr_req_desc_d_wuser_9_reg[i] <= wr_req_desc_d_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_10_reg_we[i])
               wr_req_desc_d_wuser_10_reg[i] <= uc2rb_wr_req_desc_d_wuser_10_reg[i];
             else 
               wr_req_desc_d_wuser_10_reg[i] <= wr_req_desc_d_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_11_reg_we[i])
               wr_req_desc_d_wuser_11_reg[i] <= uc2rb_wr_req_desc_d_wuser_11_reg[i];
             else 
               wr_req_desc_d_wuser_11_reg[i] <= wr_req_desc_d_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_12_reg_we[i])
               wr_req_desc_d_wuser_12_reg[i] <= uc2rb_wr_req_desc_d_wuser_12_reg[i];
             else 
               wr_req_desc_d_wuser_12_reg[i] <= wr_req_desc_d_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_13_reg_we[i])
               wr_req_desc_d_wuser_13_reg[i] <= uc2rb_wr_req_desc_d_wuser_13_reg[i];
             else 
               wr_req_desc_d_wuser_13_reg[i] <= wr_req_desc_d_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_14_reg_we[i])
               wr_req_desc_d_wuser_14_reg[i] <= uc2rb_wr_req_desc_d_wuser_14_reg[i];
             else 
               wr_req_desc_d_wuser_14_reg[i] <= wr_req_desc_d_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_D_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_d_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_d_wuser_15_reg_we[i])
               wr_req_desc_d_wuser_15_reg[i] <= uc2rb_wr_req_desc_d_wuser_15_reg[i];
             else 
               wr_req_desc_d_wuser_15_reg[i] <= wr_req_desc_d_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_D_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_d_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_d_resp_reg_we[i])
               sn_resp_desc_d_resp_reg[i] <= uc2rb_sn_resp_desc_d_resp_reg[i];
             else 
               sn_resp_desc_d_resp_reg[i] <= sn_resp_desc_d_resp_reg[i];
        end
     end
   //RD_REQ_DESC_E_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_txn_type_reg_we[i])
               rd_req_desc_e_txn_type_reg[i] <= uc2rb_rd_req_desc_e_txn_type_reg[i];
             else 
               rd_req_desc_e_txn_type_reg[i] <= rd_req_desc_e_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_E_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_size_reg_we[i])
               rd_req_desc_e_size_reg[i] <= uc2rb_rd_req_desc_e_size_reg[i];
             else 
               rd_req_desc_e_size_reg[i] <= rd_req_desc_e_size_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axsize_reg_we[i])
               rd_req_desc_e_axsize_reg[i] <= uc2rb_rd_req_desc_e_axsize_reg[i];
             else 
               rd_req_desc_e_axsize_reg[i] <= rd_req_desc_e_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_E_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_attr_reg_we[i])
               rd_req_desc_e_attr_reg[i] <= uc2rb_rd_req_desc_e_attr_reg[i];
             else 
               rd_req_desc_e_attr_reg[i] <= rd_req_desc_e_attr_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axaddr_0_reg_we[i])
               rd_req_desc_e_axaddr_0_reg[i] <= uc2rb_rd_req_desc_e_axaddr_0_reg[i];
             else 
               rd_req_desc_e_axaddr_0_reg[i] <= rd_req_desc_e_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axaddr_1_reg_we[i])
               rd_req_desc_e_axaddr_1_reg[i] <= uc2rb_rd_req_desc_e_axaddr_1_reg[i];
             else 
               rd_req_desc_e_axaddr_1_reg[i] <= rd_req_desc_e_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axaddr_2_reg_we[i])
               rd_req_desc_e_axaddr_2_reg[i] <= uc2rb_rd_req_desc_e_axaddr_2_reg[i];
             else 
               rd_req_desc_e_axaddr_2_reg[i] <= rd_req_desc_e_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axaddr_3_reg_we[i])
               rd_req_desc_e_axaddr_3_reg[i] <= uc2rb_rd_req_desc_e_axaddr_3_reg[i];
             else 
               rd_req_desc_e_axaddr_3_reg[i] <= rd_req_desc_e_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axid_0_reg_we[i])
               rd_req_desc_e_axid_0_reg[i] <= uc2rb_rd_req_desc_e_axid_0_reg[i];
             else 
               rd_req_desc_e_axid_0_reg[i] <= rd_req_desc_e_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axid_1_reg_we[i])
               rd_req_desc_e_axid_1_reg[i] <= uc2rb_rd_req_desc_e_axid_1_reg[i];
             else 
               rd_req_desc_e_axid_1_reg[i] <= rd_req_desc_e_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axid_2_reg_we[i])
               rd_req_desc_e_axid_2_reg[i] <= uc2rb_rd_req_desc_e_axid_2_reg[i];
             else 
               rd_req_desc_e_axid_2_reg[i] <= rd_req_desc_e_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axid_3_reg_we[i])
               rd_req_desc_e_axid_3_reg[i] <= uc2rb_rd_req_desc_e_axid_3_reg[i];
             else 
               rd_req_desc_e_axid_3_reg[i] <= rd_req_desc_e_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_0_reg_we[i])
               rd_req_desc_e_axuser_0_reg[i] <= uc2rb_rd_req_desc_e_axuser_0_reg[i];
             else 
               rd_req_desc_e_axuser_0_reg[i] <= rd_req_desc_e_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_1_reg_we[i])
               rd_req_desc_e_axuser_1_reg[i] <= uc2rb_rd_req_desc_e_axuser_1_reg[i];
             else 
               rd_req_desc_e_axuser_1_reg[i] <= rd_req_desc_e_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_2_reg_we[i])
               rd_req_desc_e_axuser_2_reg[i] <= uc2rb_rd_req_desc_e_axuser_2_reg[i];
             else 
               rd_req_desc_e_axuser_2_reg[i] <= rd_req_desc_e_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_3_reg_we[i])
               rd_req_desc_e_axuser_3_reg[i] <= uc2rb_rd_req_desc_e_axuser_3_reg[i];
             else 
               rd_req_desc_e_axuser_3_reg[i] <= rd_req_desc_e_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_4_reg_we[i])
               rd_req_desc_e_axuser_4_reg[i] <= uc2rb_rd_req_desc_e_axuser_4_reg[i];
             else 
               rd_req_desc_e_axuser_4_reg[i] <= rd_req_desc_e_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_5_reg_we[i])
               rd_req_desc_e_axuser_5_reg[i] <= uc2rb_rd_req_desc_e_axuser_5_reg[i];
             else 
               rd_req_desc_e_axuser_5_reg[i] <= rd_req_desc_e_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_6_reg_we[i])
               rd_req_desc_e_axuser_6_reg[i] <= uc2rb_rd_req_desc_e_axuser_6_reg[i];
             else 
               rd_req_desc_e_axuser_6_reg[i] <= rd_req_desc_e_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_7_reg_we[i])
               rd_req_desc_e_axuser_7_reg[i] <= uc2rb_rd_req_desc_e_axuser_7_reg[i];
             else 
               rd_req_desc_e_axuser_7_reg[i] <= rd_req_desc_e_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_8_reg_we[i])
               rd_req_desc_e_axuser_8_reg[i] <= uc2rb_rd_req_desc_e_axuser_8_reg[i];
             else 
               rd_req_desc_e_axuser_8_reg[i] <= rd_req_desc_e_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_9_reg_we[i])
               rd_req_desc_e_axuser_9_reg[i] <= uc2rb_rd_req_desc_e_axuser_9_reg[i];
             else 
               rd_req_desc_e_axuser_9_reg[i] <= rd_req_desc_e_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_10_reg_we[i])
               rd_req_desc_e_axuser_10_reg[i] <= uc2rb_rd_req_desc_e_axuser_10_reg[i];
             else 
               rd_req_desc_e_axuser_10_reg[i] <= rd_req_desc_e_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_11_reg_we[i])
               rd_req_desc_e_axuser_11_reg[i] <= uc2rb_rd_req_desc_e_axuser_11_reg[i];
             else 
               rd_req_desc_e_axuser_11_reg[i] <= rd_req_desc_e_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_12_reg_we[i])
               rd_req_desc_e_axuser_12_reg[i] <= uc2rb_rd_req_desc_e_axuser_12_reg[i];
             else 
               rd_req_desc_e_axuser_12_reg[i] <= rd_req_desc_e_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_13_reg_we[i])
               rd_req_desc_e_axuser_13_reg[i] <= uc2rb_rd_req_desc_e_axuser_13_reg[i];
             else 
               rd_req_desc_e_axuser_13_reg[i] <= rd_req_desc_e_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_14_reg_we[i])
               rd_req_desc_e_axuser_14_reg[i] <= uc2rb_rd_req_desc_e_axuser_14_reg[i];
             else 
               rd_req_desc_e_axuser_14_reg[i] <= rd_req_desc_e_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_E_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_e_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_e_axuser_15_reg_we[i])
               rd_req_desc_e_axuser_15_reg[i] <= uc2rb_rd_req_desc_e_axuser_15_reg[i];
             else 
               rd_req_desc_e_axuser_15_reg[i] <= rd_req_desc_e_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_E_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_txn_type_reg_we[i])
               wr_req_desc_e_txn_type_reg[i] <= uc2rb_wr_req_desc_e_txn_type_reg[i];
             else 
               wr_req_desc_e_txn_type_reg[i] <= wr_req_desc_e_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_E_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_size_reg_we[i])
               wr_req_desc_e_size_reg[i] <= uc2rb_wr_req_desc_e_size_reg[i];
             else 
               wr_req_desc_e_size_reg[i] <= wr_req_desc_e_size_reg[i];
        end
     end
   //WR_REQ_DESC_E_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_data_offset_reg_we[i])
               wr_req_desc_e_data_offset_reg[i] <= uc2rb_wr_req_desc_e_data_offset_reg[i];
             else 
               wr_req_desc_e_data_offset_reg[i] <= wr_req_desc_e_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axsize_reg_we[i])
               wr_req_desc_e_axsize_reg[i] <= uc2rb_wr_req_desc_e_axsize_reg[i];
             else 
               wr_req_desc_e_axsize_reg[i] <= wr_req_desc_e_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_E_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_attr_reg_we[i])
               wr_req_desc_e_attr_reg[i] <= uc2rb_wr_req_desc_e_attr_reg[i];
             else 
               wr_req_desc_e_attr_reg[i] <= wr_req_desc_e_attr_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axaddr_0_reg_we[i])
               wr_req_desc_e_axaddr_0_reg[i] <= uc2rb_wr_req_desc_e_axaddr_0_reg[i];
             else 
               wr_req_desc_e_axaddr_0_reg[i] <= wr_req_desc_e_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axaddr_1_reg_we[i])
               wr_req_desc_e_axaddr_1_reg[i] <= uc2rb_wr_req_desc_e_axaddr_1_reg[i];
             else 
               wr_req_desc_e_axaddr_1_reg[i] <= wr_req_desc_e_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axaddr_2_reg_we[i])
               wr_req_desc_e_axaddr_2_reg[i] <= uc2rb_wr_req_desc_e_axaddr_2_reg[i];
             else 
               wr_req_desc_e_axaddr_2_reg[i] <= wr_req_desc_e_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axaddr_3_reg_we[i])
               wr_req_desc_e_axaddr_3_reg[i] <= uc2rb_wr_req_desc_e_axaddr_3_reg[i];
             else 
               wr_req_desc_e_axaddr_3_reg[i] <= wr_req_desc_e_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axid_0_reg_we[i])
               wr_req_desc_e_axid_0_reg[i] <= uc2rb_wr_req_desc_e_axid_0_reg[i];
             else 
               wr_req_desc_e_axid_0_reg[i] <= wr_req_desc_e_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axid_1_reg_we[i])
               wr_req_desc_e_axid_1_reg[i] <= uc2rb_wr_req_desc_e_axid_1_reg[i];
             else 
               wr_req_desc_e_axid_1_reg[i] <= wr_req_desc_e_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axid_2_reg_we[i])
               wr_req_desc_e_axid_2_reg[i] <= uc2rb_wr_req_desc_e_axid_2_reg[i];
             else 
               wr_req_desc_e_axid_2_reg[i] <= wr_req_desc_e_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axid_3_reg_we[i])
               wr_req_desc_e_axid_3_reg[i] <= uc2rb_wr_req_desc_e_axid_3_reg[i];
             else 
               wr_req_desc_e_axid_3_reg[i] <= wr_req_desc_e_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_0_reg_we[i])
               wr_req_desc_e_axuser_0_reg[i] <= uc2rb_wr_req_desc_e_axuser_0_reg[i];
             else 
               wr_req_desc_e_axuser_0_reg[i] <= wr_req_desc_e_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_1_reg_we[i])
               wr_req_desc_e_axuser_1_reg[i] <= uc2rb_wr_req_desc_e_axuser_1_reg[i];
             else 
               wr_req_desc_e_axuser_1_reg[i] <= wr_req_desc_e_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_2_reg_we[i])
               wr_req_desc_e_axuser_2_reg[i] <= uc2rb_wr_req_desc_e_axuser_2_reg[i];
             else 
               wr_req_desc_e_axuser_2_reg[i] <= wr_req_desc_e_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_3_reg_we[i])
               wr_req_desc_e_axuser_3_reg[i] <= uc2rb_wr_req_desc_e_axuser_3_reg[i];
             else 
               wr_req_desc_e_axuser_3_reg[i] <= wr_req_desc_e_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_4_reg_we[i])
               wr_req_desc_e_axuser_4_reg[i] <= uc2rb_wr_req_desc_e_axuser_4_reg[i];
             else 
               wr_req_desc_e_axuser_4_reg[i] <= wr_req_desc_e_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_5_reg_we[i])
               wr_req_desc_e_axuser_5_reg[i] <= uc2rb_wr_req_desc_e_axuser_5_reg[i];
             else 
               wr_req_desc_e_axuser_5_reg[i] <= wr_req_desc_e_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_6_reg_we[i])
               wr_req_desc_e_axuser_6_reg[i] <= uc2rb_wr_req_desc_e_axuser_6_reg[i];
             else 
               wr_req_desc_e_axuser_6_reg[i] <= wr_req_desc_e_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_7_reg_we[i])
               wr_req_desc_e_axuser_7_reg[i] <= uc2rb_wr_req_desc_e_axuser_7_reg[i];
             else 
               wr_req_desc_e_axuser_7_reg[i] <= wr_req_desc_e_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_8_reg_we[i])
               wr_req_desc_e_axuser_8_reg[i] <= uc2rb_wr_req_desc_e_axuser_8_reg[i];
             else 
               wr_req_desc_e_axuser_8_reg[i] <= wr_req_desc_e_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_9_reg_we[i])
               wr_req_desc_e_axuser_9_reg[i] <= uc2rb_wr_req_desc_e_axuser_9_reg[i];
             else 
               wr_req_desc_e_axuser_9_reg[i] <= wr_req_desc_e_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_10_reg_we[i])
               wr_req_desc_e_axuser_10_reg[i] <= uc2rb_wr_req_desc_e_axuser_10_reg[i];
             else 
               wr_req_desc_e_axuser_10_reg[i] <= wr_req_desc_e_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_11_reg_we[i])
               wr_req_desc_e_axuser_11_reg[i] <= uc2rb_wr_req_desc_e_axuser_11_reg[i];
             else 
               wr_req_desc_e_axuser_11_reg[i] <= wr_req_desc_e_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_12_reg_we[i])
               wr_req_desc_e_axuser_12_reg[i] <= uc2rb_wr_req_desc_e_axuser_12_reg[i];
             else 
               wr_req_desc_e_axuser_12_reg[i] <= wr_req_desc_e_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_13_reg_we[i])
               wr_req_desc_e_axuser_13_reg[i] <= uc2rb_wr_req_desc_e_axuser_13_reg[i];
             else 
               wr_req_desc_e_axuser_13_reg[i] <= wr_req_desc_e_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_14_reg_we[i])
               wr_req_desc_e_axuser_14_reg[i] <= uc2rb_wr_req_desc_e_axuser_14_reg[i];
             else 
               wr_req_desc_e_axuser_14_reg[i] <= wr_req_desc_e_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_E_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_axuser_15_reg_we[i])
               wr_req_desc_e_axuser_15_reg[i] <= uc2rb_wr_req_desc_e_axuser_15_reg[i];
             else 
               wr_req_desc_e_axuser_15_reg[i] <= wr_req_desc_e_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_0_reg_we[i])
               wr_req_desc_e_wuser_0_reg[i] <= uc2rb_wr_req_desc_e_wuser_0_reg[i];
             else 
               wr_req_desc_e_wuser_0_reg[i] <= wr_req_desc_e_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_1_reg_we[i])
               wr_req_desc_e_wuser_1_reg[i] <= uc2rb_wr_req_desc_e_wuser_1_reg[i];
             else 
               wr_req_desc_e_wuser_1_reg[i] <= wr_req_desc_e_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_2_reg_we[i])
               wr_req_desc_e_wuser_2_reg[i] <= uc2rb_wr_req_desc_e_wuser_2_reg[i];
             else 
               wr_req_desc_e_wuser_2_reg[i] <= wr_req_desc_e_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_3_reg_we[i])
               wr_req_desc_e_wuser_3_reg[i] <= uc2rb_wr_req_desc_e_wuser_3_reg[i];
             else 
               wr_req_desc_e_wuser_3_reg[i] <= wr_req_desc_e_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_4_reg_we[i])
               wr_req_desc_e_wuser_4_reg[i] <= uc2rb_wr_req_desc_e_wuser_4_reg[i];
             else 
               wr_req_desc_e_wuser_4_reg[i] <= wr_req_desc_e_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_5_reg_we[i])
               wr_req_desc_e_wuser_5_reg[i] <= uc2rb_wr_req_desc_e_wuser_5_reg[i];
             else 
               wr_req_desc_e_wuser_5_reg[i] <= wr_req_desc_e_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_6_reg_we[i])
               wr_req_desc_e_wuser_6_reg[i] <= uc2rb_wr_req_desc_e_wuser_6_reg[i];
             else 
               wr_req_desc_e_wuser_6_reg[i] <= wr_req_desc_e_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_7_reg_we[i])
               wr_req_desc_e_wuser_7_reg[i] <= uc2rb_wr_req_desc_e_wuser_7_reg[i];
             else 
               wr_req_desc_e_wuser_7_reg[i] <= wr_req_desc_e_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_8_reg_we[i])
               wr_req_desc_e_wuser_8_reg[i] <= uc2rb_wr_req_desc_e_wuser_8_reg[i];
             else 
               wr_req_desc_e_wuser_8_reg[i] <= wr_req_desc_e_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_9_reg_we[i])
               wr_req_desc_e_wuser_9_reg[i] <= uc2rb_wr_req_desc_e_wuser_9_reg[i];
             else 
               wr_req_desc_e_wuser_9_reg[i] <= wr_req_desc_e_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_10_reg_we[i])
               wr_req_desc_e_wuser_10_reg[i] <= uc2rb_wr_req_desc_e_wuser_10_reg[i];
             else 
               wr_req_desc_e_wuser_10_reg[i] <= wr_req_desc_e_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_11_reg_we[i])
               wr_req_desc_e_wuser_11_reg[i] <= uc2rb_wr_req_desc_e_wuser_11_reg[i];
             else 
               wr_req_desc_e_wuser_11_reg[i] <= wr_req_desc_e_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_12_reg_we[i])
               wr_req_desc_e_wuser_12_reg[i] <= uc2rb_wr_req_desc_e_wuser_12_reg[i];
             else 
               wr_req_desc_e_wuser_12_reg[i] <= wr_req_desc_e_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_13_reg_we[i])
               wr_req_desc_e_wuser_13_reg[i] <= uc2rb_wr_req_desc_e_wuser_13_reg[i];
             else 
               wr_req_desc_e_wuser_13_reg[i] <= wr_req_desc_e_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_14_reg_we[i])
               wr_req_desc_e_wuser_14_reg[i] <= uc2rb_wr_req_desc_e_wuser_14_reg[i];
             else 
               wr_req_desc_e_wuser_14_reg[i] <= wr_req_desc_e_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_E_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_e_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_e_wuser_15_reg_we[i])
               wr_req_desc_e_wuser_15_reg[i] <= uc2rb_wr_req_desc_e_wuser_15_reg[i];
             else 
               wr_req_desc_e_wuser_15_reg[i] <= wr_req_desc_e_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_E_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_e_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_e_resp_reg_we[i])
               sn_resp_desc_e_resp_reg[i] <= uc2rb_sn_resp_desc_e_resp_reg[i];
             else 
               sn_resp_desc_e_resp_reg[i] <= sn_resp_desc_e_resp_reg[i];
        end
     end
   //RD_REQ_DESC_F_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_txn_type_reg_we[i])
               rd_req_desc_f_txn_type_reg[i] <= uc2rb_rd_req_desc_f_txn_type_reg[i];
             else 
               rd_req_desc_f_txn_type_reg[i] <= rd_req_desc_f_txn_type_reg[i];
        end
     end
   //RD_REQ_DESC_F_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_size_reg_we[i])
               rd_req_desc_f_size_reg[i] <= uc2rb_rd_req_desc_f_size_reg[i];
             else 
               rd_req_desc_f_size_reg[i] <= rd_req_desc_f_size_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axsize_reg_we[i])
               rd_req_desc_f_axsize_reg[i] <= uc2rb_rd_req_desc_f_axsize_reg[i];
             else 
               rd_req_desc_f_axsize_reg[i] <= rd_req_desc_f_axsize_reg[i];
        end
     end
   //RD_REQ_DESC_F_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_attr_reg_we[i])
               rd_req_desc_f_attr_reg[i] <= uc2rb_rd_req_desc_f_attr_reg[i];
             else 
               rd_req_desc_f_attr_reg[i] <= rd_req_desc_f_attr_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axaddr_0_reg_we[i])
               rd_req_desc_f_axaddr_0_reg[i] <= uc2rb_rd_req_desc_f_axaddr_0_reg[i];
             else 
               rd_req_desc_f_axaddr_0_reg[i] <= rd_req_desc_f_axaddr_0_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axaddr_1_reg_we[i])
               rd_req_desc_f_axaddr_1_reg[i] <= uc2rb_rd_req_desc_f_axaddr_1_reg[i];
             else 
               rd_req_desc_f_axaddr_1_reg[i] <= rd_req_desc_f_axaddr_1_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axaddr_2_reg_we[i])
               rd_req_desc_f_axaddr_2_reg[i] <= uc2rb_rd_req_desc_f_axaddr_2_reg[i];
             else 
               rd_req_desc_f_axaddr_2_reg[i] <= rd_req_desc_f_axaddr_2_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axaddr_3_reg_we[i])
               rd_req_desc_f_axaddr_3_reg[i] <= uc2rb_rd_req_desc_f_axaddr_3_reg[i];
             else 
               rd_req_desc_f_axaddr_3_reg[i] <= rd_req_desc_f_axaddr_3_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axid_0_reg_we[i])
               rd_req_desc_f_axid_0_reg[i] <= uc2rb_rd_req_desc_f_axid_0_reg[i];
             else 
               rd_req_desc_f_axid_0_reg[i] <= rd_req_desc_f_axid_0_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axid_1_reg_we[i])
               rd_req_desc_f_axid_1_reg[i] <= uc2rb_rd_req_desc_f_axid_1_reg[i];
             else 
               rd_req_desc_f_axid_1_reg[i] <= rd_req_desc_f_axid_1_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axid_2_reg_we[i])
               rd_req_desc_f_axid_2_reg[i] <= uc2rb_rd_req_desc_f_axid_2_reg[i];
             else 
               rd_req_desc_f_axid_2_reg[i] <= rd_req_desc_f_axid_2_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axid_3_reg_we[i])
               rd_req_desc_f_axid_3_reg[i] <= uc2rb_rd_req_desc_f_axid_3_reg[i];
             else 
               rd_req_desc_f_axid_3_reg[i] <= rd_req_desc_f_axid_3_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_0_reg_we[i])
               rd_req_desc_f_axuser_0_reg[i] <= uc2rb_rd_req_desc_f_axuser_0_reg[i];
             else 
               rd_req_desc_f_axuser_0_reg[i] <= rd_req_desc_f_axuser_0_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_1_reg_we[i])
               rd_req_desc_f_axuser_1_reg[i] <= uc2rb_rd_req_desc_f_axuser_1_reg[i];
             else 
               rd_req_desc_f_axuser_1_reg[i] <= rd_req_desc_f_axuser_1_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_2_reg_we[i])
               rd_req_desc_f_axuser_2_reg[i] <= uc2rb_rd_req_desc_f_axuser_2_reg[i];
             else 
               rd_req_desc_f_axuser_2_reg[i] <= rd_req_desc_f_axuser_2_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_3_reg_we[i])
               rd_req_desc_f_axuser_3_reg[i] <= uc2rb_rd_req_desc_f_axuser_3_reg[i];
             else 
               rd_req_desc_f_axuser_3_reg[i] <= rd_req_desc_f_axuser_3_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_4_reg_we[i])
               rd_req_desc_f_axuser_4_reg[i] <= uc2rb_rd_req_desc_f_axuser_4_reg[i];
             else 
               rd_req_desc_f_axuser_4_reg[i] <= rd_req_desc_f_axuser_4_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_5_reg_we[i])
               rd_req_desc_f_axuser_5_reg[i] <= uc2rb_rd_req_desc_f_axuser_5_reg[i];
             else 
               rd_req_desc_f_axuser_5_reg[i] <= rd_req_desc_f_axuser_5_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_6_reg_we[i])
               rd_req_desc_f_axuser_6_reg[i] <= uc2rb_rd_req_desc_f_axuser_6_reg[i];
             else 
               rd_req_desc_f_axuser_6_reg[i] <= rd_req_desc_f_axuser_6_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_7_reg_we[i])
               rd_req_desc_f_axuser_7_reg[i] <= uc2rb_rd_req_desc_f_axuser_7_reg[i];
             else 
               rd_req_desc_f_axuser_7_reg[i] <= rd_req_desc_f_axuser_7_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_8_reg_we[i])
               rd_req_desc_f_axuser_8_reg[i] <= uc2rb_rd_req_desc_f_axuser_8_reg[i];
             else 
               rd_req_desc_f_axuser_8_reg[i] <= rd_req_desc_f_axuser_8_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_9_reg_we[i])
               rd_req_desc_f_axuser_9_reg[i] <= uc2rb_rd_req_desc_f_axuser_9_reg[i];
             else 
               rd_req_desc_f_axuser_9_reg[i] <= rd_req_desc_f_axuser_9_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_10_reg_we[i])
               rd_req_desc_f_axuser_10_reg[i] <= uc2rb_rd_req_desc_f_axuser_10_reg[i];
             else 
               rd_req_desc_f_axuser_10_reg[i] <= rd_req_desc_f_axuser_10_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_11_reg_we[i])
               rd_req_desc_f_axuser_11_reg[i] <= uc2rb_rd_req_desc_f_axuser_11_reg[i];
             else 
               rd_req_desc_f_axuser_11_reg[i] <= rd_req_desc_f_axuser_11_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_12_reg_we[i])
               rd_req_desc_f_axuser_12_reg[i] <= uc2rb_rd_req_desc_f_axuser_12_reg[i];
             else 
               rd_req_desc_f_axuser_12_reg[i] <= rd_req_desc_f_axuser_12_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_13_reg_we[i])
               rd_req_desc_f_axuser_13_reg[i] <= uc2rb_rd_req_desc_f_axuser_13_reg[i];
             else 
               rd_req_desc_f_axuser_13_reg[i] <= rd_req_desc_f_axuser_13_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_14_reg_we[i])
               rd_req_desc_f_axuser_14_reg[i] <= uc2rb_rd_req_desc_f_axuser_14_reg[i];
             else 
               rd_req_desc_f_axuser_14_reg[i] <= rd_req_desc_f_axuser_14_reg[i];
        end
     end
   //RD_REQ_DESC_F_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             rd_req_desc_f_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_rd_req_desc_f_axuser_15_reg_we[i])
               rd_req_desc_f_axuser_15_reg[i] <= uc2rb_rd_req_desc_f_axuser_15_reg[i];
             else 
               rd_req_desc_f_axuser_15_reg[i] <= rd_req_desc_f_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_F_TXN_TYPE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_txn_type_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_txn_type_reg_we[i])
               wr_req_desc_f_txn_type_reg[i] <= uc2rb_wr_req_desc_f_txn_type_reg[i];
             else 
               wr_req_desc_f_txn_type_reg[i] <= wr_req_desc_f_txn_type_reg[i];
        end
     end
   //WR_REQ_DESC_F_SIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_size_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_size_reg_we[i])
               wr_req_desc_f_size_reg[i] <= uc2rb_wr_req_desc_f_size_reg[i];
             else 
               wr_req_desc_f_size_reg[i] <= wr_req_desc_f_size_reg[i];
        end
     end
   //WR_REQ_DESC_F_DATA_OFFSET_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_data_offset_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_data_offset_reg_we[i])
               wr_req_desc_f_data_offset_reg[i] <= uc2rb_wr_req_desc_f_data_offset_reg[i];
             else 
               wr_req_desc_f_data_offset_reg[i] <= wr_req_desc_f_data_offset_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXSIZE_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axsize_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axsize_reg_we[i])
               wr_req_desc_f_axsize_reg[i] <= uc2rb_wr_req_desc_f_axsize_reg[i];
             else 
               wr_req_desc_f_axsize_reg[i] <= wr_req_desc_f_axsize_reg[i];
        end
     end
   //WR_REQ_DESC_F_ATTR_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_attr_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_attr_reg_we[i])
               wr_req_desc_f_attr_reg[i] <= uc2rb_wr_req_desc_f_attr_reg[i];
             else 
               wr_req_desc_f_attr_reg[i] <= wr_req_desc_f_attr_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXADDR_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axaddr_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axaddr_0_reg_we[i])
               wr_req_desc_f_axaddr_0_reg[i] <= uc2rb_wr_req_desc_f_axaddr_0_reg[i];
             else 
               wr_req_desc_f_axaddr_0_reg[i] <= wr_req_desc_f_axaddr_0_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXADDR_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axaddr_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axaddr_1_reg_we[i])
               wr_req_desc_f_axaddr_1_reg[i] <= uc2rb_wr_req_desc_f_axaddr_1_reg[i];
             else 
               wr_req_desc_f_axaddr_1_reg[i] <= wr_req_desc_f_axaddr_1_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXADDR_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axaddr_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axaddr_2_reg_we[i])
               wr_req_desc_f_axaddr_2_reg[i] <= uc2rb_wr_req_desc_f_axaddr_2_reg[i];
             else 
               wr_req_desc_f_axaddr_2_reg[i] <= wr_req_desc_f_axaddr_2_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXADDR_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axaddr_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axaddr_3_reg_we[i])
               wr_req_desc_f_axaddr_3_reg[i] <= uc2rb_wr_req_desc_f_axaddr_3_reg[i];
             else 
               wr_req_desc_f_axaddr_3_reg[i] <= wr_req_desc_f_axaddr_3_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXID_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axid_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axid_0_reg_we[i])
               wr_req_desc_f_axid_0_reg[i] <= uc2rb_wr_req_desc_f_axid_0_reg[i];
             else 
               wr_req_desc_f_axid_0_reg[i] <= wr_req_desc_f_axid_0_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXID_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axid_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axid_1_reg_we[i])
               wr_req_desc_f_axid_1_reg[i] <= uc2rb_wr_req_desc_f_axid_1_reg[i];
             else 
               wr_req_desc_f_axid_1_reg[i] <= wr_req_desc_f_axid_1_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXID_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axid_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axid_2_reg_we[i])
               wr_req_desc_f_axid_2_reg[i] <= uc2rb_wr_req_desc_f_axid_2_reg[i];
             else 
               wr_req_desc_f_axid_2_reg[i] <= wr_req_desc_f_axid_2_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXID_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axid_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axid_3_reg_we[i])
               wr_req_desc_f_axid_3_reg[i] <= uc2rb_wr_req_desc_f_axid_3_reg[i];
             else 
               wr_req_desc_f_axid_3_reg[i] <= wr_req_desc_f_axid_3_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_0_reg_we[i])
               wr_req_desc_f_axuser_0_reg[i] <= uc2rb_wr_req_desc_f_axuser_0_reg[i];
             else 
               wr_req_desc_f_axuser_0_reg[i] <= wr_req_desc_f_axuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_1_reg_we[i])
               wr_req_desc_f_axuser_1_reg[i] <= uc2rb_wr_req_desc_f_axuser_1_reg[i];
             else 
               wr_req_desc_f_axuser_1_reg[i] <= wr_req_desc_f_axuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_2_reg_we[i])
               wr_req_desc_f_axuser_2_reg[i] <= uc2rb_wr_req_desc_f_axuser_2_reg[i];
             else 
               wr_req_desc_f_axuser_2_reg[i] <= wr_req_desc_f_axuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_3_reg_we[i])
               wr_req_desc_f_axuser_3_reg[i] <= uc2rb_wr_req_desc_f_axuser_3_reg[i];
             else 
               wr_req_desc_f_axuser_3_reg[i] <= wr_req_desc_f_axuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_4_reg_we[i])
               wr_req_desc_f_axuser_4_reg[i] <= uc2rb_wr_req_desc_f_axuser_4_reg[i];
             else 
               wr_req_desc_f_axuser_4_reg[i] <= wr_req_desc_f_axuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_5_reg_we[i])
               wr_req_desc_f_axuser_5_reg[i] <= uc2rb_wr_req_desc_f_axuser_5_reg[i];
             else 
               wr_req_desc_f_axuser_5_reg[i] <= wr_req_desc_f_axuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_6_reg_we[i])
               wr_req_desc_f_axuser_6_reg[i] <= uc2rb_wr_req_desc_f_axuser_6_reg[i];
             else 
               wr_req_desc_f_axuser_6_reg[i] <= wr_req_desc_f_axuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_7_reg_we[i])
               wr_req_desc_f_axuser_7_reg[i] <= uc2rb_wr_req_desc_f_axuser_7_reg[i];
             else 
               wr_req_desc_f_axuser_7_reg[i] <= wr_req_desc_f_axuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_8_reg_we[i])
               wr_req_desc_f_axuser_8_reg[i] <= uc2rb_wr_req_desc_f_axuser_8_reg[i];
             else 
               wr_req_desc_f_axuser_8_reg[i] <= wr_req_desc_f_axuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_9_reg_we[i])
               wr_req_desc_f_axuser_9_reg[i] <= uc2rb_wr_req_desc_f_axuser_9_reg[i];
             else 
               wr_req_desc_f_axuser_9_reg[i] <= wr_req_desc_f_axuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_10_reg_we[i])
               wr_req_desc_f_axuser_10_reg[i] <= uc2rb_wr_req_desc_f_axuser_10_reg[i];
             else 
               wr_req_desc_f_axuser_10_reg[i] <= wr_req_desc_f_axuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_11_reg_we[i])
               wr_req_desc_f_axuser_11_reg[i] <= uc2rb_wr_req_desc_f_axuser_11_reg[i];
             else 
               wr_req_desc_f_axuser_11_reg[i] <= wr_req_desc_f_axuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_12_reg_we[i])
               wr_req_desc_f_axuser_12_reg[i] <= uc2rb_wr_req_desc_f_axuser_12_reg[i];
             else 
               wr_req_desc_f_axuser_12_reg[i] <= wr_req_desc_f_axuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_13_reg_we[i])
               wr_req_desc_f_axuser_13_reg[i] <= uc2rb_wr_req_desc_f_axuser_13_reg[i];
             else 
               wr_req_desc_f_axuser_13_reg[i] <= wr_req_desc_f_axuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_14_reg_we[i])
               wr_req_desc_f_axuser_14_reg[i] <= uc2rb_wr_req_desc_f_axuser_14_reg[i];
             else 
               wr_req_desc_f_axuser_14_reg[i] <= wr_req_desc_f_axuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_F_AXUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_axuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_axuser_15_reg_we[i])
               wr_req_desc_f_axuser_15_reg[i] <= uc2rb_wr_req_desc_f_axuser_15_reg[i];
             else 
               wr_req_desc_f_axuser_15_reg[i] <= wr_req_desc_f_axuser_15_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_0_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_0_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_0_reg_we[i])
               wr_req_desc_f_wuser_0_reg[i] <= uc2rb_wr_req_desc_f_wuser_0_reg[i];
             else 
               wr_req_desc_f_wuser_0_reg[i] <= wr_req_desc_f_wuser_0_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_1_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_1_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_1_reg_we[i])
               wr_req_desc_f_wuser_1_reg[i] <= uc2rb_wr_req_desc_f_wuser_1_reg[i];
             else 
               wr_req_desc_f_wuser_1_reg[i] <= wr_req_desc_f_wuser_1_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_2_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_2_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_2_reg_we[i])
               wr_req_desc_f_wuser_2_reg[i] <= uc2rb_wr_req_desc_f_wuser_2_reg[i];
             else 
               wr_req_desc_f_wuser_2_reg[i] <= wr_req_desc_f_wuser_2_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_3_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_3_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_3_reg_we[i])
               wr_req_desc_f_wuser_3_reg[i] <= uc2rb_wr_req_desc_f_wuser_3_reg[i];
             else 
               wr_req_desc_f_wuser_3_reg[i] <= wr_req_desc_f_wuser_3_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_4_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_4_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_4_reg_we[i])
               wr_req_desc_f_wuser_4_reg[i] <= uc2rb_wr_req_desc_f_wuser_4_reg[i];
             else 
               wr_req_desc_f_wuser_4_reg[i] <= wr_req_desc_f_wuser_4_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_5_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_5_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_5_reg_we[i])
               wr_req_desc_f_wuser_5_reg[i] <= uc2rb_wr_req_desc_f_wuser_5_reg[i];
             else 
               wr_req_desc_f_wuser_5_reg[i] <= wr_req_desc_f_wuser_5_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_6_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_6_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_6_reg_we[i])
               wr_req_desc_f_wuser_6_reg[i] <= uc2rb_wr_req_desc_f_wuser_6_reg[i];
             else 
               wr_req_desc_f_wuser_6_reg[i] <= wr_req_desc_f_wuser_6_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_7_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_7_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_7_reg_we[i])
               wr_req_desc_f_wuser_7_reg[i] <= uc2rb_wr_req_desc_f_wuser_7_reg[i];
             else 
               wr_req_desc_f_wuser_7_reg[i] <= wr_req_desc_f_wuser_7_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_8_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_8_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_8_reg_we[i])
               wr_req_desc_f_wuser_8_reg[i] <= uc2rb_wr_req_desc_f_wuser_8_reg[i];
             else 
               wr_req_desc_f_wuser_8_reg[i] <= wr_req_desc_f_wuser_8_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_9_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_9_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_9_reg_we[i])
               wr_req_desc_f_wuser_9_reg[i] <= uc2rb_wr_req_desc_f_wuser_9_reg[i];
             else 
               wr_req_desc_f_wuser_9_reg[i] <= wr_req_desc_f_wuser_9_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_10_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_10_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_10_reg_we[i])
               wr_req_desc_f_wuser_10_reg[i] <= uc2rb_wr_req_desc_f_wuser_10_reg[i];
             else 
               wr_req_desc_f_wuser_10_reg[i] <= wr_req_desc_f_wuser_10_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_11_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_11_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_11_reg_we[i])
               wr_req_desc_f_wuser_11_reg[i] <= uc2rb_wr_req_desc_f_wuser_11_reg[i];
             else 
               wr_req_desc_f_wuser_11_reg[i] <= wr_req_desc_f_wuser_11_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_12_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_12_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_12_reg_we[i])
               wr_req_desc_f_wuser_12_reg[i] <= uc2rb_wr_req_desc_f_wuser_12_reg[i];
             else 
               wr_req_desc_f_wuser_12_reg[i] <= wr_req_desc_f_wuser_12_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_13_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_13_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_13_reg_we[i])
               wr_req_desc_f_wuser_13_reg[i] <= uc2rb_wr_req_desc_f_wuser_13_reg[i];
             else 
               wr_req_desc_f_wuser_13_reg[i] <= wr_req_desc_f_wuser_13_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_14_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_14_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_14_reg_we[i])
               wr_req_desc_f_wuser_14_reg[i] <= uc2rb_wr_req_desc_f_wuser_14_reg[i];
             else 
               wr_req_desc_f_wuser_14_reg[i] <= wr_req_desc_f_wuser_14_reg[i];
        end
     end
   //WR_REQ_DESC_F_WUSER_15_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             wr_req_desc_f_wuser_15_reg[i] <= 1'h0;
           else 
             if (uc2rb_wr_req_desc_f_wuser_15_reg_we[i])
               wr_req_desc_f_wuser_15_reg[i] <= uc2rb_wr_req_desc_f_wuser_15_reg[i];
             else 
               wr_req_desc_f_wuser_15_reg[i] <= wr_req_desc_f_wuser_15_reg[i];
        end
     end
   //SN_RESP_DESC_F_RESP_REG
   always @( posedge clk )
     begin
        for (i = 0; i < 32 ; i = i + 1) begin
           if (~rst_n)
             sn_resp_desc_f_resp_reg[i] <= 1'h0;
           else 
             if (uc2rb_sn_resp_desc_f_resp_reg_we[i])
               sn_resp_desc_f_resp_reg[i] <= uc2rb_sn_resp_desc_f_resp_reg[i];
             else 
               sn_resp_desc_f_resp_reg[i] <= sn_resp_desc_f_resp_reg[i];
        end
     end


   // RAMS


   always @(posedge clk)
     begin
	if ( ~rst_n)
          begin
             wdata_ram_addr   <= 'h0;     
          end
	else begin
           if (~mode_select_reg[0]) begin
              if (~axi_araddr[BRIDGE_MSB] && axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2])begin //AXI RD targeted to WDATA RAM
		 if (~wdata_ram_rd_en) begin
                    if (arvalid_pending_pulse)begin
                       wdata_ram_rd_en <= 1'b1;
                       if (S_ACE_USR_XX_DATA_WIDTH == 128)
			 wdata_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:4];
                       else if (S_ACE_USR_XX_DATA_WIDTH == 64)
			 wdata_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:3];
                       else if (S_ACE_USR_XX_DATA_WIDTH == 32)                    
			 wdata_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:2];
                    end
                    else begin
                       wdata_ram_addr   <= 'h0;
                       wdata_ram_rd_en  <= 1'b0;
                    end // else: !if(arvalid_pending_pulse)
		 end // if (~wdata_ram_rd_en)
		 else begin
                    wdata_ram_addr   <= 'h0;
                    wdata_ram_rd_en  <= 1'b0;
		 end // else: !if(~wdata_ram_rd_en)
              end 
              else begin
                 wdata_ram_addr   <= 'h0;
                 wdata_ram_rd_en  <= 1'b0;
              end // else: !if(~axi_araddr[16] && axi_araddr[15] && ~axi_araddr[14])
           end
           else begin
              wdata_ram_addr   <= hm2rb_rd_addr;
              wdata_ram_rd_en  <= 1'b1;
           end // else: !if(~mode_select_reg[0])
	end // else: !if( ~rst_n)
     end // always @ (posedge clk)
   
   
   always @( posedge clk )
     begin
        if ( rst_n == 1'b0 )
          begin
             wdata_ram_data_ready  <= 0;
             wdata_ram_data_ready_1  <= 0;
             wdata_ram_data_ready_2  <= 0;
          end 
        else
          if (~axi_araddr[BRIDGE_MSB] && axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2]) begin
             wdata_ram_data_ready_1 <= wdata_ram_rd_en;
             wdata_ram_data_ready_2 <= wdata_ram_data_ready_1;
             wdata_ram_data_ready <= wdata_ram_data_ready_2;
          end
          else begin
             wdata_ram_data_ready  <= 0;
             wdata_ram_data_ready_1  <= 0;
             wdata_ram_data_ready_2  <= 0;
          end
     end // always @ ( posedge clk )
   




   // Output register or memory read data
   always @( posedge clk )
     begin
        if ( rst_n == 1'b0 )
          begin
             axi_rdata  <= 0;
          end 
        
        
        else if (axi_rvalid) 
          begin    
             axi_rdata  <= axi_rdata;
          end 


        else 
          begin    
             // When there is a valid read address (S_AXI_ARVALID) with 
             // acceptance of read address by the slave (axi_arready), 
             // output the read dada 
             if (~axi_araddr[BRIDGE_MSB] && axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2] && (~mode_select_reg[0]) )begin  //WDATA RAM
                if (wdata_ram_data_ready) begin
                   if (S_ACE_USR_XX_DATA_WIDTH == 128)begin
                      case (axi_araddr[3:2])
                        2'b00: axi_rdata <= wdata_ram_data[31:0];     //data from WDATA RAM
                        2'b01: axi_rdata <= wdata_ram_data[63:32];
                        2'b10: axi_rdata <= wdata_ram_data[95:64];
                        2'b11: axi_rdata <= wdata_ram_data[127:96];
                      endcase // case (axi_araddr[3:2])
                   end
                   else begin
                      if (S_ACE_USR_XX_DATA_WIDTH == 64)begin
                         case (axi_araddr[2])
                           1'b0: axi_rdata <= wdata_ram_data[31:0];
                           1'b1: axi_rdata <= wdata_ram_data[63:32];
                         endcase // case (axi_araddr[2])
                      end
                      else begin 
                         if (S_ACE_USR_XX_DATA_WIDTH == 32)                    
                           axi_rdata <= wdata_ram_data;
                      end
                   end // else: !if(S_ACE_USR_XX_DATA_WIDTH == 128)
                end
                else begin
	           axi_rdata <= axi_rdata;
                end // else: !if(wdata_ram_data_ready)
             end
             else if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && ~axi_araddr[BRIDGE_MSB-2] && (~mode_select_reg[0]) )begin //WSTRB RAM
                if (wstrb_ram_data_ready) begin
                   if (S_ACE_USR_XX_DATA_WIDTH == 128)begin
                      case (axi_araddr[3:2])
                        2'b00: axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[3]} }, { 8{wstrb_ram_data[2]} }, { 8{wstrb_ram_data[1]} }, { 8{wstrb_ram_data[0]} } } : {28'b0,wstrb_ram_data[3:0] } ;     //data from WSTRB RAM
                        2'b01: axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[7]} }, { 8{wstrb_ram_data[6]} }, { 8{wstrb_ram_data[5]} }, { 8{wstrb_ram_data[4]} } } : {28'b0,wstrb_ram_data[7:4]};
                        2'b10: axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[11]} }, { 8{wstrb_ram_data[10]} }, { 8{wstrb_ram_data[9]} }, { 8{wstrb_ram_data[8]} } } : {28'b0,wstrb_ram_data[11:8]};
                        2'b11: axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[15]} }, { 8{wstrb_ram_data[14]} }, { 8{wstrb_ram_data[13]} }, { 8{wstrb_ram_data[12]} } } : {28'b0,wstrb_ram_data[15:12]};
                      endcase // case (axi_araddr[3:2])
                   end
                   else begin
                      if (S_ACE_USR_XX_DATA_WIDTH == 64)begin
                         case (axi_araddr[2])
                           1'b0: axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[3]} }, { 8{wstrb_ram_data[2]} }, { 8{wstrb_ram_data[1]} }, { 8{wstrb_ram_data[0]} } } : {28'b0,wstrb_ram_data[3:0]};
                           1'b1: axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[7]} }, { 8{wstrb_ram_data[6]} }, { 8{wstrb_ram_data[5]} }, { 8{wstrb_ram_data[4]} } } : {28'b0,wstrb_ram_data[7:4]};
                         endcase // case (axi_araddr[2])
                      end
                      else begin 
                         if (S_ACE_USR_XX_DATA_WIDTH == 32)                    
                           axi_rdata <= (EXTEND_WSTRB==1) ? { { 8{wstrb_ram_data[3]} }, { 8{wstrb_ram_data[2]} }, { 8{wstrb_ram_data[1]} }, { 8{wstrb_ram_data[0]} } } : {28'b0,  wstrb_ram_data[3:0] };
                      end
                   end // else: !if(S_ACE_USR_XX_DATA_WIDTH == 128)
                end
                else
		  axi_rdata <= axi_rdata;
             end // if (axi_araddr[16] && ~axi_araddr[15] && ~axi_araddr[14])
             else if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2] && ~(|axi_araddr[BRIDGE_MSB-3:BRIDGE_MSB-6]))begin //CDDATA RAM
                if (cddata_ram_data_ready) begin
                   if (S_ACE_USR_SN_DATA_WIDTH == 128)begin
                      case (axi_araddr[3:2])
                        2'b00: axi_rdata <= cddata_ram_data[31:0];     //data from WDATA RAM
                        2'b01: axi_rdata <= cddata_ram_data[63:32];
                        2'b10: axi_rdata <= cddata_ram_data[95:64];
                        2'b11: axi_rdata <= cddata_ram_data[127:96];
                      endcase // case (axi_araddr[3:2])
                   end
                   else begin
                      if (S_ACE_USR_SN_DATA_WIDTH == 64)begin
                         case (axi_araddr[2])
                           1'b0: axi_rdata <= cddata_ram_data[31:0];
                           1'b1: axi_rdata <= cddata_ram_data[63:32];
                         endcase // case (axi_araddr[2])
                      end
                      else begin 
                         if (S_ACE_USR_SN_DATA_WIDTH == 32)                    
                           axi_rdata <= cddata_ram_data;
                      end
                   end // else: !if(S_ACE_USR_SN_DATA_WIDTH == 128)
                end
                else begin
	           axi_rdata <= axi_rdata;
                end // else: !if(cddata_ram_data_ready)
             end // if (axi_araddr[16] && ~axi_araddr[15] && ~axi_araddr[14])
             
             else begin
                rb2hm_rd_data <= wdata_ram_data;
                rb2hm_rd_wstrb <= wstrb_ram_data;

                if (match_fifo_pop_desc==1'b1) begin

                   if ( (~|axi_araddr[BRIDGE_MSB:10]) && (axi_araddr[9:0]==`RD_REQ_FIFO_POP_DESC_REG_ADDR) )begin  //fifo_pop_desc 
                      axi_rdata <= {rd_req_fifo_out_valid,{(32-(`CLOG2(XX_MAX_DESC))-1){1'b0}},rd_req_fifo_out[(`CLOG2(XX_MAX_DESC))-1:0]};
                   end
                   else if ( (~|axi_araddr[BRIDGE_MSB:10]) && (axi_araddr[9:0]==`WR_REQ_FIFO_POP_DESC_REG_ADDR) )begin  //fifo_pop_desc 
                      axi_rdata <= {wr_req_fifo_out_valid,{(32-(`CLOG2(XX_MAX_DESC))-1){1'b0}},wr_req_fifo_out[(`CLOG2(XX_MAX_DESC))-1:0]};
                   end
                   else if ( (~|axi_araddr[BRIDGE_MSB:10]) && (axi_araddr[9:0]==`SN_RESP_FIFO_POP_DESC_REG_ADDR) )begin  //fifo_pop_desc 
                      axi_rdata <= {sn_resp_fifo_out_valid,{(32-(`CLOG2(SN_MAX_DESC))-1){1'b0}},sn_resp_fifo_out[(`CLOG2(SN_MAX_DESC))-1:0]};
                   end
                   else if ( (~|axi_araddr[BRIDGE_MSB:10]) && (axi_araddr[9:0]==`SN_DATA_FIFO_POP_DESC_REG_ADDR) )begin  //fifo_pop_desc 
                      axi_rdata <= {sn_data_fifo_out_valid,{(32-(`CLOG2(SN_MAX_DESC))-1){1'b0}},sn_data_fifo_out[(`CLOG2(SN_MAX_DESC))-1:0]};
                   end              
                   
                end          
                else begin
                   axi_rdata <= reg_data_out_pipeline;               
                end

             end // else: !if(~mode_select_reg[0])
          end
     end


   always @( posedge clk )
     begin
        if ( rst_n == 1'b0 )
          begin
             match_fifo_pop_desc <= 1'b0;
          end
        else if ( (~|axi_araddr[BRIDGE_MSB:10]) && ( (axi_araddr[9:0]==`RD_REQ_FIFO_POP_DESC_REG_ADDR) || (axi_araddr[9:0]==`WR_REQ_FIFO_POP_DESC_REG_ADDR) || (axi_araddr[9:0]==`SN_RESP_FIFO_POP_DESC_REG_ADDR) || (axi_araddr[9:0]==`SN_DATA_FIFO_POP_DESC_REG_ADDR) ) )
          begin
             match_fifo_pop_desc <= 1'b1;
          end
        else 
          begin
             match_fifo_pop_desc <= 1'b0;
          end
     end
   
   
   


   // Implement axi_rvalid generation
   // axi_rvalid is asserted for one AXI_ACLK clock cycle when both 
   // S_AXI_ARVALID and axi_arready are asserted. The slave registers 
   // data are available on the axi_rdata bus at this instance. The 
   // assertion of axi_rvalid marks the validity of read data on the 
   // bus and axi_rresp indicates the status of read transaction.axi_rvalid 
   // is deasserted on reset (active low). axi_rresp and axi_rdata are 
   // cleared to zero on reset (active low).  
   always @( posedge clk )
     begin
        if ( resetn == 1'b0 )
          begin
             axi_rvalid <= 0;
             axi_rresp  <= 0;
          end 
        else
          begin    
             if (axi_arready && s_axi_arvalid && ~axi_rvalid)
               begin
                  if (~axi_araddr[BRIDGE_MSB] && axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2]) //WDATA RAM
                    if (wdata_ram_data_ready) begin
                       axi_rvalid <= 1'b1;
                       axi_rresp  <= 2'b0; // 'OKAY' response
                    end
                    else
                      axi_rvalid <= 1'b0;
                  else begin
                     if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && ~axi_araddr[BRIDGE_MSB-2]) //WSTRB RAM
                       if (wstrb_ram_data_ready) begin
                          axi_rvalid <= 1'b1;
                          axi_rresp  <= 2'b0; // 'OKAY' response
                       end
                       else
                         axi_rvalid <= 1'b0;
                     if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2] && ~(|axi_araddr[BRIDGE_MSB-3:BRIDGE_MSB-6])) //CDDATA RAM
                       if (cddata_ram_data_ready) begin
                          axi_rvalid <= 1'b1;
                          axi_rresp  <= 2'b0; // 'OKAY' response
                       end
                       else
                         axi_rvalid <= 1'b0;
                     else begin
                        // Valid read data is available at the read data bus
                        axi_rvalid <= 1'b1;
                        axi_rresp  <= 2'b0; // 'OKAY' response
                     end // else: !if(wdata_ram_data_ready)
                  end // if (axi_arready && s_axi_arvalid && ~axi_rvalid)
               end
             else if (axi_rvalid && s_axi_rready)
               begin
                  // Read data is accepted by the master
                  axi_rvalid <= 1'b0;
               end
             
          end // else: !if( resetn == 1'b0 )
     end // always @ ( posedge clk )




   data_ram #(
              .AWIDTH (`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8))), // Address Width
              .DWIDTH (S_ACE_USR_XX_DATA_WIDTH),  // Data Width
              .OREG_A ("TRUE"),  // Optional Port A output pipeline registers
              .OREG_B ("TRUE")   // Optional Port B output pipeline registers  
              )
   u_wdata_ram (
                .clk        (clk), 
                .rst_a      (~rst_n), 
                .en_a       (uc2rb_wr_we), 
                .we_a       (1'b1), // Port A is always Write port
                .byte_en_a  (uc2rb_wr_bwe),
                .addr_a     (uc2rb_wr_addr), 
                .wr_data_a  (uc2rb_wr_data), 
                .rd_data_a  (), 
                .OREG_CE_A  (1'b1),                 
                .rst_b      (~rst_n), 
                .en_b       (wdata_ram_rd_en), 
                .we_b       (1'b0), // Port B is alwyas Read port 
                .addr_b     (wdata_ram_addr), 
                .rd_data_b  (wdata_ram_data), 
                .byte_en_b  ({(S_ACE_USR_XX_DATA_WIDTH/8){1'h0}}),
                .wr_data_b  ({(S_ACE_USR_XX_DATA_WIDTH){1'h0}}), 
                .OREG_CE_B  (1'b1));





   always @(posedge clk)
     begin
	if ( ~rst_n)
          begin
             wstrb_ram_addr   <= 'h0;     
          end
	else begin
           if (~mode_select_reg[0]) begin
              if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && ~axi_araddr[BRIDGE_MSB-2])begin //AXI RD targeted to WSTRB RAM
		 if (~wstrb_ram_rd_en) begin
                    if (arvalid_pending_pulse)begin
                       wstrb_ram_rd_en <= 1'b1;
                       if (S_ACE_USR_XX_DATA_WIDTH == 128)
			 wstrb_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:4];
                       else if (S_ACE_USR_XX_DATA_WIDTH == 64)
			 wstrb_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:3];
                       else if (S_ACE_USR_XX_DATA_WIDTH == 32)                    
			 wstrb_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:2];
                    end
                    else begin
                       wstrb_ram_addr   <= 'h0;
                       wstrb_ram_rd_en  <= 1'b0;
                    end // else: !if(arvalid_pending_pulse)
		 end // if (~wstrb_ram_rd_en)
		 else begin
                    wstrb_ram_addr   <= 'h0;
                    wstrb_ram_rd_en  <= 1'b0;
		 end // else: !if(~wstrb_ram_rd_en)
              end 
              else begin
                 wstrb_ram_addr   <= 'h0;
                 wstrb_ram_rd_en  <= 1'b0;
              end // else: !if(~axi_araddr[16] && axi_araddr[15] && ~axi_araddr[14])
           end
           else begin
              wstrb_ram_addr   <= hm2rb_rd_addr;
              wstrb_ram_rd_en  <= 1'b1;
           end // else: !if(~mode_select_reg[0])
	end // else: !if( ~rst_n)
     end // always @ (posedge clk)
   



   
   always @( posedge clk )
     begin
        if ( rst_n == 1'b0 )
          begin
             wstrb_ram_data_ready  <= 0;
             wstrb_ram_data_ready_1  <= 0;
             wstrb_ram_data_ready_2  <= 0;
          end 
        else
          if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && ~axi_araddr[BRIDGE_MSB-2]) begin
             wstrb_ram_data_ready_1 <= wstrb_ram_rd_en;
             wstrb_ram_data_ready_2 <= wstrb_ram_data_ready_1;
             wstrb_ram_data_ready <= wstrb_ram_data_ready_2;
          end
          else begin
             wstrb_ram_data_ready  <= 0;
             wstrb_ram_data_ready_1  <= 0;
             wstrb_ram_data_ready_2  <= 0;
          end
     end // always @ ( posedge clk )
   




   strb_ram #(
              .AWIDTH (`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8))), // Address Width
              .DWIDTH ((S_ACE_USR_XX_DATA_WIDTH/8)),  // Data Width
              .OREG_A ("TRUE"),  // Optional Port A output pipeline registers
              .OREG_B ("TRUE")   // Optional Port B output pipeline registers  
              )
   u_wstrb_ram (
                .clk        (clk), 
                .rst_a      (~rst_n), 
                .en_a       (uc2rb_wr_we), 
                .we_a       (1'b1), // Port A is always Write port
                .nibble_en_a  ({(S_ACE_USR_XX_DATA_WIDTH/32){1'b1}}),
                .addr_a     (uc2rb_wr_addr), 
                .wr_data_a  (uc2rb_wr_wstrb), 
                .rd_data_a  ( ), 
                .OREG_CE_A  (1'b1),                 
                .rst_b      (~rst_n), 
                .en_b       (wstrb_ram_rd_en), 
                .we_b       (1'b0), // Port B is alwyas Read port 
                .addr_b     (wstrb_ram_addr), 
                .rd_data_b  (wstrb_ram_data), 
                .nibble_en_b({(S_ACE_USR_XX_DATA_WIDTH/32){1'h0}}),   //({ ((S_ACE_USR_XX_DATA_WIDTH/8)/4) {1'h0}}),
                .wr_data_b  ({(S_ACE_USR_XX_DATA_WIDTH/8){1'h0}}), 
                .OREG_CE_B  (1'b1));



   // RD DATA RAM
   
   always @(posedge clk)
     begin
	if ( ~rst_n)
          begin
             rdata_ram_we   <= 'h0;     
             rdata_ram_addr <= 'h0;     
             rdata_ram_data <= 'h0;
             rdata_ram_bwe  <= 'h0;
          end
	else begin
           if (~mode_select_reg[0]) begin
              if (reg_wr_en) begin
		 if (~axi_awaddr[BRIDGE_MSB] && axi_awaddr[BRIDGE_MSB-1] && ~axi_awaddr[BRIDGE_MSB-2])begin //AXI WR targeted to RD DATA RAM
                    rdata_ram_we <= 1'b1;
                    if (S_ACE_USR_XX_DATA_WIDTH == 128)begin
                       rdata_ram_addr <= axi_awaddr[S_AXI_ADDR_WIDTH-1:4];
                       rdata_ram_data <= {4{s_axi_wdata}};
                       rdata_ram_bwe <= { ({4{axi_awaddr[3] && axi_awaddr[2]}} & s_axi_wstrb) , ({4{axi_awaddr[3] && ~axi_awaddr[2]}} & s_axi_wstrb) , ({4{~axi_awaddr[3] && axi_awaddr[2]}} & s_axi_wstrb) , ({4{~axi_awaddr[3] && ~axi_awaddr[2]}} & s_axi_wstrb) };
                    end
                    else if (S_ACE_USR_XX_DATA_WIDTH == 64)begin
                       rdata_ram_addr <= axi_awaddr[S_AXI_ADDR_WIDTH-1:3];
                       rdata_ram_data <= {2{s_axi_wdata}};
                       rdata_ram_bwe  <= {({4{axi_awaddr[2]}} & s_axi_wstrb),({4{~axi_awaddr[2]}} & s_axi_wstrb)};
                    end
                    else if (S_ACE_USR_XX_DATA_WIDTH == 32)begin
                       rdata_ram_addr <= axi_awaddr[S_AXI_ADDR_WIDTH-1:2];
                       rdata_ram_data <= s_axi_wdata;
                       rdata_ram_bwe  <= s_axi_wstrb;
                    end
		 end
		 else begin
                    rdata_ram_we <= 1'b0;
                    rdata_ram_addr <= 'h0;     
                    rdata_ram_data <= 'h0;
                    rdata_ram_bwe  <= 'h0;
		 end // 
              end            
              else begin 
		 rdata_ram_we <= 1'b0;
		 rdata_ram_addr <= 'h0;     
		 rdata_ram_data <= 'h0;
		 rdata_ram_bwe  <= 'h0;
              end // if (reg_wr_en)
           end
           
           else begin
              rdata_ram_we   <= hm2rb_wr_we;     
              rdata_ram_bwe  <= hm2rb_wr_bwe;
              rdata_ram_addr <= hm2rb_wr_addr;     
              rdata_ram_data <= hm2rb_wr_data;
           end // else: !if(reg_wr_en)
	end // else: !if( ~rst_n)
     end // always @ (posedge clk)
   
   
   // Registering uc2rb_rd_addr

   always @( posedge clk )
     begin
        if (~rst_n)
          uc2rb_rd_addr_reg <= 'h0;
        else 
          uc2rb_rd_addr_reg <= uc2rb_rd_addr;
     end

   data_ram #(
              .AWIDTH (`CLOG2(XX_RAM_SIZE/(S_ACE_USR_XX_DATA_WIDTH/8))), // Address Width
              .DWIDTH (S_ACE_USR_XX_DATA_WIDTH),  // Data Width
              .OREG_A ("TRUE"),  // Optional Port A output pipeline registers
              .OREG_B ("TRUE")   // Optional Port B output pipeline registers  
              )
   u_rdata_ram (
                .clk        (clk), 
                .rst_a      (~rst_n), 
                .en_a       (rdata_ram_we), 
                .we_a       (1'b1), // Port A is always Write port
                .byte_en_a  (rdata_ram_bwe),
                .addr_a     (rdata_ram_addr), 
                .wr_data_a  (rdata_ram_data), 
                .rd_data_a  (), 
                .OREG_CE_A  (1'b1),                 
                .rst_b      (~rst_n), 
                .en_b       (1'b1), 
                .we_b       (1'b0), // Port B is alwyas Read port 
                .addr_b     (uc2rb_rd_addr_reg), 
                .rd_data_b  (rb2uc_rd_data), 
                .byte_en_b  ({(S_ACE_USR_XX_DATA_WIDTH/8){1'h0}}),
                .wr_data_b  ({(S_ACE_USR_XX_DATA_WIDTH){1'h0}}), 
                .OREG_CE_B  (1'b1));

   
   

   always @(posedge clk)
     begin
	if ( ~rst_n)
          begin
             cddata_ram_addr   <= 'h0;     
          end
	else begin
           if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2] && ~(|axi_araddr[BRIDGE_MSB-3:BRIDGE_MSB-6]))begin //AXI RD targeted to CDDATA RAM
              if (~cddata_ram_rd_en) begin
                 if (arvalid_pending_pulse)begin
                    cddata_ram_rd_en <= 1'b1;
                    if (S_ACE_USR_SN_DATA_WIDTH == 128)
                      cddata_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:4];
                    else if (S_ACE_USR_SN_DATA_WIDTH == 64)
                      cddata_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:3];
                    else if (S_ACE_USR_SN_DATA_WIDTH == 32)                    
                      cddata_ram_addr <= axi_araddr[S_AXI_ADDR_WIDTH-1:2];
                    else                                   
                      cddata_ram_addr <= 'h0;
                 end
                 else begin
                    cddata_ram_addr   <= 'h0;
                    cddata_ram_rd_en  <= 1'b0;
                 end // else: !if(arvalid_pending_pulse)
              end // if (~cddata_ram_rd_en)
              else begin
                 cddata_ram_addr   <= 'h0;
                 cddata_ram_rd_en  <= 1'b0;
              end // else: !if(~cddata_ram_rd_en)
           end 
           else begin
              cddata_ram_addr   <= 'h0;
              cddata_ram_rd_en  <= 1'b0;
           end // else: !if(~axi_araddr[16] && axi_araddr[15] && ~axi_araddr[14])
	end // else: !if( ~rst_n)
     end // always @ (posedge clk)
   
   
   
   always @( posedge clk )
     begin
        if ( rst_n == 1'b0 )
          begin
             cddata_ram_data_ready  <= 0;
             cddata_ram_data_ready_1  <= 0;
             cddata_ram_data_ready_2  <= 0;
          end 
        else
          if (axi_araddr[BRIDGE_MSB] && ~axi_araddr[BRIDGE_MSB-1] && axi_araddr[BRIDGE_MSB-2] && ~(|axi_araddr[BRIDGE_MSB-3:BRIDGE_MSB-6])) begin
             cddata_ram_data_ready_1 <= cddata_ram_rd_en;
             cddata_ram_data_ready_2 <= cddata_ram_data_ready_1;
             cddata_ram_data_ready <= cddata_ram_data_ready_2;
          end
          else begin
             cddata_ram_data_ready  <= 0;
             cddata_ram_data_ready_1  <= 0;
             cddata_ram_data_ready_2  <= 0;
          end
     end // always @ ( posedge clk )
   



   
   
   



   data_ram #(
              .AWIDTH (`CLOG2(SN_RAM_SIZE/(S_ACE_USR_SN_DATA_WIDTH/8))), // Address Width
              .DWIDTH (S_ACE_USR_SN_DATA_WIDTH),  // Data Width
              .OREG_A ("TRUE"),  // Optional Port A output pipeline registers
              .OREG_B ("TRUE")   // Optional Port B output pipeline registers  
              )
   u_cddata_ram (
                 .clk        (clk), 
                 .rst_a      (~rst_n), 
                 .en_a       (uc2rb_sn_we), 
                 .we_a       (1'b1), // Port A is always Write port
                 .byte_en_a  (uc2rb_sn_bwe),
                 .addr_a     (uc2rb_sn_addr), 
                 .wr_data_a  (uc2rb_sn_data), 
                 .rd_data_a  (), 
                 .OREG_CE_A  (1'b1),                 
                 .rst_b      (~rst_n), 
                 .en_b       (cddata_ram_rd_en), 
                 .we_b       (1'b0), // Port B is alwyas Read port 
                 .addr_b     (cddata_ram_addr), 
                 .rd_data_b  (cddata_ram_data), 
                 .byte_en_b  ({(S_ACE_USR_SN_DATA_WIDTH/8){1'h0}}),
                 .wr_data_b  ({(S_ACE_USR_SN_DATA_WIDTH){1'h0}}), 
                 .OREG_CE_B  (1'b1));




   

   
endmodule // regs_slave

/* regs_slave.v ends here */
