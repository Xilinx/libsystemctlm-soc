/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *   This module directly handshakes with Register block, Host Control
 *   block. 
 *
 *
 */

`include "ace_defines_common.vh"
module ace_usr_mst_control #(

                             parameter ACE_PROTOCOL                   = "FULLACE" 
                             
                             ,parameter M_ACE_USR_ADDR_WIDTH           = 64 
                             ,parameter M_ACE_USR_XX_DATA_WIDTH        = 128       
                             ,parameter M_ACE_USR_SN_DATA_WIDTH        = 128       
                             ,parameter M_ACE_USR_ID_WIDTH             = 16 
                             ,parameter M_ACE_USR_AWUSER_WIDTH         = 32 
                             ,parameter M_ACE_USR_WUSER_WIDTH          = 32 
                             ,parameter M_ACE_USR_BUSER_WIDTH          = 32 
                             ,parameter M_ACE_USR_ARUSER_WIDTH         = 32 
                             ,parameter M_ACE_USR_RUSER_WIDTH          = 32 
                             
                             ,parameter CACHE_LINE_SIZE                = 64 
                             ,parameter XX_MAX_DESC                    = 16         
                             ,parameter SN_MAX_DESC                    = 16         
                             ,parameter XX_RAM_SIZE                    = 16384     
                             ,parameter SN_RAM_SIZE                    = 1024       

                             )(

                               //Clock and reset
                               input clk 
			       ,input resetn
   
			       //M_ACE_USR
			       ,output[M_ACE_USR_ID_WIDTH-1:0] m_ace_usr_awid 
			       ,output[M_ACE_USR_ADDR_WIDTH-1:0] m_ace_usr_awaddr 
			       ,output[7:0] m_ace_usr_awlen
			       ,output[2:0] m_ace_usr_awsize 
			       ,output[1:0] m_ace_usr_awburst 
			       ,output m_ace_usr_awlock 
			       ,output[3:0] m_ace_usr_awcache 
			       ,output[2:0] m_ace_usr_awprot 
			       ,output[3:0] m_ace_usr_awqos 
			       ,output[3:0] m_ace_usr_awregion 
			       ,output[M_ACE_USR_AWUSER_WIDTH-1:0] m_ace_usr_awuser 
			       ,output[2:0] m_ace_usr_awsnoop 
			       ,output[1:0] m_ace_usr_awdomain 
			       ,output[1:0] m_ace_usr_awbar 
			       ,output m_ace_usr_awunique 
			       ,output m_ace_usr_awvalid 
			       ,input m_ace_usr_awready 
			       ,output[M_ACE_USR_XX_DATA_WIDTH-1:0] m_ace_usr_wdata 
			       ,output[(M_ACE_USR_XX_DATA_WIDTH/8)-1:0] m_ace_usr_wstrb
			       ,output m_ace_usr_wlast 
			       ,output[M_ACE_USR_WUSER_WIDTH-1:0] m_ace_usr_wuser 
			       ,output m_ace_usr_wvalid 
			       ,input m_ace_usr_wready 
			       ,input [M_ACE_USR_ID_WIDTH-1:0] m_ace_usr_bid 
			       ,input [1:0] m_ace_usr_bresp 
			       ,input [M_ACE_USR_BUSER_WIDTH-1:0] m_ace_usr_buser 
			       ,input m_ace_usr_bvalid 
			       ,output m_ace_usr_bready 
			       ,output m_ace_usr_wack 
			       ,output[M_ACE_USR_ID_WIDTH-1:0] m_ace_usr_arid 
			       ,output[M_ACE_USR_ADDR_WIDTH-1:0] m_ace_usr_araddr 
			       ,output[7:0] m_ace_usr_arlen 
			       ,output[2:0] m_ace_usr_arsize 
			       ,output[1:0] m_ace_usr_arburst 
			       ,output m_ace_usr_arlock 
			       ,output[3:0] m_ace_usr_arcache 
			       ,output[2:0] m_ace_usr_arprot 
			       ,output[3:0] m_ace_usr_arqos 
			       ,output[3:0] m_ace_usr_arregion 
			       ,output[M_ACE_USR_ARUSER_WIDTH-1:0] m_ace_usr_aruser 
			       ,output[3:0] m_ace_usr_arsnoop 
			       ,output[1:0] m_ace_usr_ardomain 
			       ,output[1:0] m_ace_usr_arbar 
			       ,output m_ace_usr_arvalid 
			       ,input m_ace_usr_arready 
			       ,input [M_ACE_USR_ID_WIDTH-1:0] m_ace_usr_rid 
			       ,input [M_ACE_USR_XX_DATA_WIDTH-1:0] m_ace_usr_rdata 
			       ,input [3:0] m_ace_usr_rresp 
			       ,input m_ace_usr_rlast 
			       ,input [M_ACE_USR_RUSER_WIDTH-1:0] m_ace_usr_ruser 
			       ,input m_ace_usr_rvalid 
			       ,output m_ace_usr_rready 
			       ,output m_ace_usr_rack 
			       ,input [M_ACE_USR_ADDR_WIDTH-1:0] m_ace_usr_acaddr 
			       ,input [3:0] m_ace_usr_acsnoop 
			       ,input [2:0] m_ace_usr_acprot 
			       ,input m_ace_usr_acvalid 
			       ,output m_ace_usr_acready 
			       ,output [4:0] m_ace_usr_crresp 
			       ,output m_ace_usr_crvalid 
			       ,input m_ace_usr_crready 
			       ,output [M_ACE_USR_SN_DATA_WIDTH-1:0] m_ace_usr_cddata 
			       ,output m_ace_usr_cdlast 
			       ,output m_ace_usr_cdvalid 
			       ,input m_ace_usr_cdready 
   
			       ,input [31:0] bridge_identification_reg
			       ,input [31:0] last_bridge_reg
			       ,input [31:0] version_reg
			       ,input [31:0] bridge_type_reg
			       ,input [31:0] mode_select_reg
			       ,input [31:0] reset_reg
			       ,input [31:0] h2c_intr_0_reg
			       ,input [31:0] h2c_intr_1_reg
			       ,input [31:0] h2c_intr_2_reg
			       ,input [31:0] h2c_intr_3_reg
			       ,input [31:0] c2h_intr_status_0_reg
			       ,input [31:0] intr_c2h_toggle_status_0_reg
			       ,input [31:0] intr_c2h_toggle_clear_0_reg
			       ,input [31:0] intr_c2h_toggle_enable_0_reg
			       ,input [31:0] c2h_intr_status_1_reg
			       ,input [31:0] intr_c2h_toggle_status_1_reg
			       ,input [31:0] intr_c2h_toggle_clear_1_reg
			       ,input [31:0] intr_c2h_toggle_enable_1_reg
			       ,input [31:0] c2h_gpio_0_reg
			       ,input [31:0] c2h_gpio_1_reg
			       ,input [31:0] c2h_gpio_2_reg
			       ,input [31:0] c2h_gpio_3_reg
			       ,input [31:0] c2h_gpio_4_reg
			       ,input [31:0] c2h_gpio_5_reg
			       ,input [31:0] c2h_gpio_6_reg
			       ,input [31:0] c2h_gpio_7_reg
			       ,input [31:0] c2h_gpio_8_reg
			       ,input [31:0] c2h_gpio_9_reg
			       ,input [31:0] c2h_gpio_10_reg
			       ,input [31:0] c2h_gpio_11_reg
			       ,input [31:0] c2h_gpio_12_reg
			       ,input [31:0] c2h_gpio_13_reg
			       ,input [31:0] c2h_gpio_14_reg
			       ,input [31:0] c2h_gpio_15_reg
			       ,input [31:0] h2c_gpio_0_reg
			       ,input [31:0] h2c_gpio_1_reg
			       ,input [31:0] h2c_gpio_2_reg
			       ,input [31:0] h2c_gpio_3_reg
			       ,input [31:0] h2c_gpio_4_reg
			       ,input [31:0] h2c_gpio_5_reg
			       ,input [31:0] h2c_gpio_6_reg
			       ,input [31:0] h2c_gpio_7_reg
			       ,input [31:0] h2c_gpio_8_reg
			       ,input [31:0] h2c_gpio_9_reg
			       ,input [31:0] h2c_gpio_10_reg
			       ,input [31:0] h2c_gpio_11_reg
			       ,input [31:0] h2c_gpio_12_reg
			       ,input [31:0] h2c_gpio_13_reg
			       ,input [31:0] h2c_gpio_14_reg
			       ,input [31:0] h2c_gpio_15_reg
			       ,input [31:0] bridge_config_reg
			       ,input [31:0] intr_status_reg
			       ,input [31:0] intr_error_status_reg
			       ,input [31:0] intr_error_clear_reg
			       ,input [31:0] intr_error_enable_reg
			       ,input [31:0] bridge_rd_user_config_reg
			       ,input [31:0] bridge_wr_user_config_reg
			       ,input [31:0] rd_max_desc_reg
			       ,input [31:0] wr_max_desc_reg
			       ,input [31:0] sn_max_desc_reg
			       ,input [31:0] rd_req_fifo_push_desc_reg
			       ,input [31:0] rd_req_fifo_free_level_reg
			       ,input [31:0] rd_req_intr_comp_status_reg
			       ,input [31:0] rd_req_intr_comp_clear_reg
			       ,input [31:0] rd_req_intr_comp_enable_reg
			       ,input [31:0] rd_resp_free_desc_reg
			       ,input [31:0] rd_resp_fifo_pop_desc_reg
			       ,input [31:0] rd_resp_fifo_fill_level_reg
			       ,input [31:0] wr_req_fifo_push_desc_reg
			       ,input [31:0] wr_req_fifo_free_level_reg
			       ,input [31:0] wr_req_intr_comp_status_reg
			       ,input [31:0] wr_req_intr_comp_clear_reg
			       ,input [31:0] wr_req_intr_comp_enable_reg
			       ,input [31:0] wr_resp_free_desc_reg
			       ,input [31:0] wr_resp_fifo_pop_desc_reg
			       ,input [31:0] wr_resp_fifo_fill_level_reg
			       ,input [31:0] sn_req_free_desc_reg
			       ,input [31:0] sn_req_fifo_pop_desc_reg
			       ,input [31:0] sn_req_fifo_fill_level_reg
			       ,input [31:0] sn_resp_fifo_push_desc_reg
			       ,input [31:0] sn_resp_fifo_free_level_reg
			       ,input [31:0] sn_resp_intr_comp_status_reg
			       ,input [31:0] sn_resp_intr_comp_clear_reg
			       ,input [31:0] sn_resp_intr_comp_enable_reg
			       ,input [31:0] sn_data_fifo_push_desc_reg
			       ,input [31:0] sn_data_fifo_free_level_reg
			       ,input [31:0] sn_data_intr_comp_status_reg
			       ,input [31:0] sn_data_intr_comp_clear_reg
			       ,input [31:0] sn_data_intr_comp_enable_reg
			       ,input [31:0] intr_fifo_enable_reg
			       ,input [31:0] rd_req_desc_0_txn_type_reg
			       ,input [31:0] rd_req_desc_0_size_reg
			       ,input [31:0] rd_req_desc_0_axsize_reg
			       ,input [31:0] rd_req_desc_0_attr_reg
			       ,input [31:0] rd_req_desc_0_axaddr_0_reg
			       ,input [31:0] rd_req_desc_0_axaddr_1_reg
			       ,input [31:0] rd_req_desc_0_axaddr_2_reg
			       ,input [31:0] rd_req_desc_0_axaddr_3_reg
			       ,input [31:0] rd_req_desc_0_axid_0_reg
			       ,input [31:0] rd_req_desc_0_axid_1_reg
			       ,input [31:0] rd_req_desc_0_axid_2_reg
			       ,input [31:0] rd_req_desc_0_axid_3_reg
			       ,input [31:0] rd_req_desc_0_axuser_0_reg
			       ,input [31:0] rd_req_desc_0_axuser_1_reg
			       ,input [31:0] rd_req_desc_0_axuser_2_reg
			       ,input [31:0] rd_req_desc_0_axuser_3_reg
			       ,input [31:0] rd_req_desc_0_axuser_4_reg
			       ,input [31:0] rd_req_desc_0_axuser_5_reg
			       ,input [31:0] rd_req_desc_0_axuser_6_reg
			       ,input [31:0] rd_req_desc_0_axuser_7_reg
			       ,input [31:0] rd_req_desc_0_axuser_8_reg
			       ,input [31:0] rd_req_desc_0_axuser_9_reg
			       ,input [31:0] rd_req_desc_0_axuser_10_reg
			       ,input [31:0] rd_req_desc_0_axuser_11_reg
			       ,input [31:0] rd_req_desc_0_axuser_12_reg
			       ,input [31:0] rd_req_desc_0_axuser_13_reg
			       ,input [31:0] rd_req_desc_0_axuser_14_reg
			       ,input [31:0] rd_req_desc_0_axuser_15_reg
			       ,input [31:0] rd_resp_desc_0_data_offset_reg
			       ,input [31:0] rd_resp_desc_0_data_size_reg
			       ,input [31:0] rd_resp_desc_0_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_0_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_0_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_0_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_0_resp_reg
			       ,input [31:0] rd_resp_desc_0_xid_0_reg
			       ,input [31:0] rd_resp_desc_0_xid_1_reg
			       ,input [31:0] rd_resp_desc_0_xid_2_reg
			       ,input [31:0] rd_resp_desc_0_xid_3_reg
			       ,input [31:0] rd_resp_desc_0_xuser_0_reg
			       ,input [31:0] rd_resp_desc_0_xuser_1_reg
			       ,input [31:0] rd_resp_desc_0_xuser_2_reg
			       ,input [31:0] rd_resp_desc_0_xuser_3_reg
			       ,input [31:0] rd_resp_desc_0_xuser_4_reg
			       ,input [31:0] rd_resp_desc_0_xuser_5_reg
			       ,input [31:0] rd_resp_desc_0_xuser_6_reg
			       ,input [31:0] rd_resp_desc_0_xuser_7_reg
			       ,input [31:0] rd_resp_desc_0_xuser_8_reg
			       ,input [31:0] rd_resp_desc_0_xuser_9_reg
			       ,input [31:0] rd_resp_desc_0_xuser_10_reg
			       ,input [31:0] rd_resp_desc_0_xuser_11_reg
			       ,input [31:0] rd_resp_desc_0_xuser_12_reg
			       ,input [31:0] rd_resp_desc_0_xuser_13_reg
			       ,input [31:0] rd_resp_desc_0_xuser_14_reg
			       ,input [31:0] rd_resp_desc_0_xuser_15_reg
			       ,input [31:0] wr_req_desc_0_txn_type_reg
			       ,input [31:0] wr_req_desc_0_size_reg
			       ,input [31:0] wr_req_desc_0_data_offset_reg
			       ,input [31:0] wr_req_desc_0_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_0_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_0_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_0_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_0_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_0_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_0_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_0_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_0_axsize_reg
			       ,input [31:0] wr_req_desc_0_attr_reg
			       ,input [31:0] wr_req_desc_0_axaddr_0_reg
			       ,input [31:0] wr_req_desc_0_axaddr_1_reg
			       ,input [31:0] wr_req_desc_0_axaddr_2_reg
			       ,input [31:0] wr_req_desc_0_axaddr_3_reg
			       ,input [31:0] wr_req_desc_0_axid_0_reg
			       ,input [31:0] wr_req_desc_0_axid_1_reg
			       ,input [31:0] wr_req_desc_0_axid_2_reg
			       ,input [31:0] wr_req_desc_0_axid_3_reg
			       ,input [31:0] wr_req_desc_0_axuser_0_reg
			       ,input [31:0] wr_req_desc_0_axuser_1_reg
			       ,input [31:0] wr_req_desc_0_axuser_2_reg
			       ,input [31:0] wr_req_desc_0_axuser_3_reg
			       ,input [31:0] wr_req_desc_0_axuser_4_reg
			       ,input [31:0] wr_req_desc_0_axuser_5_reg
			       ,input [31:0] wr_req_desc_0_axuser_6_reg
			       ,input [31:0] wr_req_desc_0_axuser_7_reg
			       ,input [31:0] wr_req_desc_0_axuser_8_reg
			       ,input [31:0] wr_req_desc_0_axuser_9_reg
			       ,input [31:0] wr_req_desc_0_axuser_10_reg
			       ,input [31:0] wr_req_desc_0_axuser_11_reg
			       ,input [31:0] wr_req_desc_0_axuser_12_reg
			       ,input [31:0] wr_req_desc_0_axuser_13_reg
			       ,input [31:0] wr_req_desc_0_axuser_14_reg
			       ,input [31:0] wr_req_desc_0_axuser_15_reg
			       ,input [31:0] wr_req_desc_0_wuser_0_reg
			       ,input [31:0] wr_req_desc_0_wuser_1_reg
			       ,input [31:0] wr_req_desc_0_wuser_2_reg
			       ,input [31:0] wr_req_desc_0_wuser_3_reg
			       ,input [31:0] wr_req_desc_0_wuser_4_reg
			       ,input [31:0] wr_req_desc_0_wuser_5_reg
			       ,input [31:0] wr_req_desc_0_wuser_6_reg
			       ,input [31:0] wr_req_desc_0_wuser_7_reg
			       ,input [31:0] wr_req_desc_0_wuser_8_reg
			       ,input [31:0] wr_req_desc_0_wuser_9_reg
			       ,input [31:0] wr_req_desc_0_wuser_10_reg
			       ,input [31:0] wr_req_desc_0_wuser_11_reg
			       ,input [31:0] wr_req_desc_0_wuser_12_reg
			       ,input [31:0] wr_req_desc_0_wuser_13_reg
			       ,input [31:0] wr_req_desc_0_wuser_14_reg
			       ,input [31:0] wr_req_desc_0_wuser_15_reg
			       ,input [31:0] wr_resp_desc_0_resp_reg
			       ,input [31:0] wr_resp_desc_0_xid_0_reg
			       ,input [31:0] wr_resp_desc_0_xid_1_reg
			       ,input [31:0] wr_resp_desc_0_xid_2_reg
			       ,input [31:0] wr_resp_desc_0_xid_3_reg
			       ,input [31:0] wr_resp_desc_0_xuser_0_reg
			       ,input [31:0] wr_resp_desc_0_xuser_1_reg
			       ,input [31:0] wr_resp_desc_0_xuser_2_reg
			       ,input [31:0] wr_resp_desc_0_xuser_3_reg
			       ,input [31:0] wr_resp_desc_0_xuser_4_reg
			       ,input [31:0] wr_resp_desc_0_xuser_5_reg
			       ,input [31:0] wr_resp_desc_0_xuser_6_reg
			       ,input [31:0] wr_resp_desc_0_xuser_7_reg
			       ,input [31:0] wr_resp_desc_0_xuser_8_reg
			       ,input [31:0] wr_resp_desc_0_xuser_9_reg
			       ,input [31:0] wr_resp_desc_0_xuser_10_reg
			       ,input [31:0] wr_resp_desc_0_xuser_11_reg
			       ,input [31:0] wr_resp_desc_0_xuser_12_reg
			       ,input [31:0] wr_resp_desc_0_xuser_13_reg
			       ,input [31:0] wr_resp_desc_0_xuser_14_reg
			       ,input [31:0] wr_resp_desc_0_xuser_15_reg
			       ,input [31:0] sn_req_desc_0_attr_reg
			       ,input [31:0] sn_req_desc_0_acaddr_0_reg
			       ,input [31:0] sn_req_desc_0_acaddr_1_reg
			       ,input [31:0] sn_req_desc_0_acaddr_2_reg
			       ,input [31:0] sn_req_desc_0_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_0_resp_reg
			       ,input [31:0] rd_req_desc_1_txn_type_reg
			       ,input [31:0] rd_req_desc_1_size_reg
			       ,input [31:0] rd_req_desc_1_axsize_reg
			       ,input [31:0] rd_req_desc_1_attr_reg
			       ,input [31:0] rd_req_desc_1_axaddr_0_reg
			       ,input [31:0] rd_req_desc_1_axaddr_1_reg
			       ,input [31:0] rd_req_desc_1_axaddr_2_reg
			       ,input [31:0] rd_req_desc_1_axaddr_3_reg
			       ,input [31:0] rd_req_desc_1_axid_0_reg
			       ,input [31:0] rd_req_desc_1_axid_1_reg
			       ,input [31:0] rd_req_desc_1_axid_2_reg
			       ,input [31:0] rd_req_desc_1_axid_3_reg
			       ,input [31:0] rd_req_desc_1_axuser_0_reg
			       ,input [31:0] rd_req_desc_1_axuser_1_reg
			       ,input [31:0] rd_req_desc_1_axuser_2_reg
			       ,input [31:0] rd_req_desc_1_axuser_3_reg
			       ,input [31:0] rd_req_desc_1_axuser_4_reg
			       ,input [31:0] rd_req_desc_1_axuser_5_reg
			       ,input [31:0] rd_req_desc_1_axuser_6_reg
			       ,input [31:0] rd_req_desc_1_axuser_7_reg
			       ,input [31:0] rd_req_desc_1_axuser_8_reg
			       ,input [31:0] rd_req_desc_1_axuser_9_reg
			       ,input [31:0] rd_req_desc_1_axuser_10_reg
			       ,input [31:0] rd_req_desc_1_axuser_11_reg
			       ,input [31:0] rd_req_desc_1_axuser_12_reg
			       ,input [31:0] rd_req_desc_1_axuser_13_reg
			       ,input [31:0] rd_req_desc_1_axuser_14_reg
			       ,input [31:0] rd_req_desc_1_axuser_15_reg
			       ,input [31:0] rd_resp_desc_1_data_offset_reg
			       ,input [31:0] rd_resp_desc_1_data_size_reg
			       ,input [31:0] rd_resp_desc_1_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_1_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_1_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_1_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_1_resp_reg
			       ,input [31:0] rd_resp_desc_1_xid_0_reg
			       ,input [31:0] rd_resp_desc_1_xid_1_reg
			       ,input [31:0] rd_resp_desc_1_xid_2_reg
			       ,input [31:0] rd_resp_desc_1_xid_3_reg
			       ,input [31:0] rd_resp_desc_1_xuser_0_reg
			       ,input [31:0] rd_resp_desc_1_xuser_1_reg
			       ,input [31:0] rd_resp_desc_1_xuser_2_reg
			       ,input [31:0] rd_resp_desc_1_xuser_3_reg
			       ,input [31:0] rd_resp_desc_1_xuser_4_reg
			       ,input [31:0] rd_resp_desc_1_xuser_5_reg
			       ,input [31:0] rd_resp_desc_1_xuser_6_reg
			       ,input [31:0] rd_resp_desc_1_xuser_7_reg
			       ,input [31:0] rd_resp_desc_1_xuser_8_reg
			       ,input [31:0] rd_resp_desc_1_xuser_9_reg
			       ,input [31:0] rd_resp_desc_1_xuser_10_reg
			       ,input [31:0] rd_resp_desc_1_xuser_11_reg
			       ,input [31:0] rd_resp_desc_1_xuser_12_reg
			       ,input [31:0] rd_resp_desc_1_xuser_13_reg
			       ,input [31:0] rd_resp_desc_1_xuser_14_reg
			       ,input [31:0] rd_resp_desc_1_xuser_15_reg
			       ,input [31:0] wr_req_desc_1_txn_type_reg
			       ,input [31:0] wr_req_desc_1_size_reg
			       ,input [31:0] wr_req_desc_1_data_offset_reg
			       ,input [31:0] wr_req_desc_1_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_1_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_1_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_1_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_1_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_1_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_1_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_1_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_1_axsize_reg
			       ,input [31:0] wr_req_desc_1_attr_reg
			       ,input [31:0] wr_req_desc_1_axaddr_0_reg
			       ,input [31:0] wr_req_desc_1_axaddr_1_reg
			       ,input [31:0] wr_req_desc_1_axaddr_2_reg
			       ,input [31:0] wr_req_desc_1_axaddr_3_reg
			       ,input [31:0] wr_req_desc_1_axid_0_reg
			       ,input [31:0] wr_req_desc_1_axid_1_reg
			       ,input [31:0] wr_req_desc_1_axid_2_reg
			       ,input [31:0] wr_req_desc_1_axid_3_reg
			       ,input [31:0] wr_req_desc_1_axuser_0_reg
			       ,input [31:0] wr_req_desc_1_axuser_1_reg
			       ,input [31:0] wr_req_desc_1_axuser_2_reg
			       ,input [31:0] wr_req_desc_1_axuser_3_reg
			       ,input [31:0] wr_req_desc_1_axuser_4_reg
			       ,input [31:0] wr_req_desc_1_axuser_5_reg
			       ,input [31:0] wr_req_desc_1_axuser_6_reg
			       ,input [31:0] wr_req_desc_1_axuser_7_reg
			       ,input [31:0] wr_req_desc_1_axuser_8_reg
			       ,input [31:0] wr_req_desc_1_axuser_9_reg
			       ,input [31:0] wr_req_desc_1_axuser_10_reg
			       ,input [31:0] wr_req_desc_1_axuser_11_reg
			       ,input [31:0] wr_req_desc_1_axuser_12_reg
			       ,input [31:0] wr_req_desc_1_axuser_13_reg
			       ,input [31:0] wr_req_desc_1_axuser_14_reg
			       ,input [31:0] wr_req_desc_1_axuser_15_reg
			       ,input [31:0] wr_req_desc_1_wuser_0_reg
			       ,input [31:0] wr_req_desc_1_wuser_1_reg
			       ,input [31:0] wr_req_desc_1_wuser_2_reg
			       ,input [31:0] wr_req_desc_1_wuser_3_reg
			       ,input [31:0] wr_req_desc_1_wuser_4_reg
			       ,input [31:0] wr_req_desc_1_wuser_5_reg
			       ,input [31:0] wr_req_desc_1_wuser_6_reg
			       ,input [31:0] wr_req_desc_1_wuser_7_reg
			       ,input [31:0] wr_req_desc_1_wuser_8_reg
			       ,input [31:0] wr_req_desc_1_wuser_9_reg
			       ,input [31:0] wr_req_desc_1_wuser_10_reg
			       ,input [31:0] wr_req_desc_1_wuser_11_reg
			       ,input [31:0] wr_req_desc_1_wuser_12_reg
			       ,input [31:0] wr_req_desc_1_wuser_13_reg
			       ,input [31:0] wr_req_desc_1_wuser_14_reg
			       ,input [31:0] wr_req_desc_1_wuser_15_reg
			       ,input [31:0] wr_resp_desc_1_resp_reg
			       ,input [31:0] wr_resp_desc_1_xid_0_reg
			       ,input [31:0] wr_resp_desc_1_xid_1_reg
			       ,input [31:0] wr_resp_desc_1_xid_2_reg
			       ,input [31:0] wr_resp_desc_1_xid_3_reg
			       ,input [31:0] wr_resp_desc_1_xuser_0_reg
			       ,input [31:0] wr_resp_desc_1_xuser_1_reg
			       ,input [31:0] wr_resp_desc_1_xuser_2_reg
			       ,input [31:0] wr_resp_desc_1_xuser_3_reg
			       ,input [31:0] wr_resp_desc_1_xuser_4_reg
			       ,input [31:0] wr_resp_desc_1_xuser_5_reg
			       ,input [31:0] wr_resp_desc_1_xuser_6_reg
			       ,input [31:0] wr_resp_desc_1_xuser_7_reg
			       ,input [31:0] wr_resp_desc_1_xuser_8_reg
			       ,input [31:0] wr_resp_desc_1_xuser_9_reg
			       ,input [31:0] wr_resp_desc_1_xuser_10_reg
			       ,input [31:0] wr_resp_desc_1_xuser_11_reg
			       ,input [31:0] wr_resp_desc_1_xuser_12_reg
			       ,input [31:0] wr_resp_desc_1_xuser_13_reg
			       ,input [31:0] wr_resp_desc_1_xuser_14_reg
			       ,input [31:0] wr_resp_desc_1_xuser_15_reg
			       ,input [31:0] sn_req_desc_1_attr_reg
			       ,input [31:0] sn_req_desc_1_acaddr_0_reg
			       ,input [31:0] sn_req_desc_1_acaddr_1_reg
			       ,input [31:0] sn_req_desc_1_acaddr_2_reg
			       ,input [31:0] sn_req_desc_1_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_1_resp_reg
			       ,input [31:0] rd_req_desc_2_txn_type_reg
			       ,input [31:0] rd_req_desc_2_size_reg
			       ,input [31:0] rd_req_desc_2_axsize_reg
			       ,input [31:0] rd_req_desc_2_attr_reg
			       ,input [31:0] rd_req_desc_2_axaddr_0_reg
			       ,input [31:0] rd_req_desc_2_axaddr_1_reg
			       ,input [31:0] rd_req_desc_2_axaddr_2_reg
			       ,input [31:0] rd_req_desc_2_axaddr_3_reg
			       ,input [31:0] rd_req_desc_2_axid_0_reg
			       ,input [31:0] rd_req_desc_2_axid_1_reg
			       ,input [31:0] rd_req_desc_2_axid_2_reg
			       ,input [31:0] rd_req_desc_2_axid_3_reg
			       ,input [31:0] rd_req_desc_2_axuser_0_reg
			       ,input [31:0] rd_req_desc_2_axuser_1_reg
			       ,input [31:0] rd_req_desc_2_axuser_2_reg
			       ,input [31:0] rd_req_desc_2_axuser_3_reg
			       ,input [31:0] rd_req_desc_2_axuser_4_reg
			       ,input [31:0] rd_req_desc_2_axuser_5_reg
			       ,input [31:0] rd_req_desc_2_axuser_6_reg
			       ,input [31:0] rd_req_desc_2_axuser_7_reg
			       ,input [31:0] rd_req_desc_2_axuser_8_reg
			       ,input [31:0] rd_req_desc_2_axuser_9_reg
			       ,input [31:0] rd_req_desc_2_axuser_10_reg
			       ,input [31:0] rd_req_desc_2_axuser_11_reg
			       ,input [31:0] rd_req_desc_2_axuser_12_reg
			       ,input [31:0] rd_req_desc_2_axuser_13_reg
			       ,input [31:0] rd_req_desc_2_axuser_14_reg
			       ,input [31:0] rd_req_desc_2_axuser_15_reg
			       ,input [31:0] rd_resp_desc_2_data_offset_reg
			       ,input [31:0] rd_resp_desc_2_data_size_reg
			       ,input [31:0] rd_resp_desc_2_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_2_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_2_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_2_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_2_resp_reg
			       ,input [31:0] rd_resp_desc_2_xid_0_reg
			       ,input [31:0] rd_resp_desc_2_xid_1_reg
			       ,input [31:0] rd_resp_desc_2_xid_2_reg
			       ,input [31:0] rd_resp_desc_2_xid_3_reg
			       ,input [31:0] rd_resp_desc_2_xuser_0_reg
			       ,input [31:0] rd_resp_desc_2_xuser_1_reg
			       ,input [31:0] rd_resp_desc_2_xuser_2_reg
			       ,input [31:0] rd_resp_desc_2_xuser_3_reg
			       ,input [31:0] rd_resp_desc_2_xuser_4_reg
			       ,input [31:0] rd_resp_desc_2_xuser_5_reg
			       ,input [31:0] rd_resp_desc_2_xuser_6_reg
			       ,input [31:0] rd_resp_desc_2_xuser_7_reg
			       ,input [31:0] rd_resp_desc_2_xuser_8_reg
			       ,input [31:0] rd_resp_desc_2_xuser_9_reg
			       ,input [31:0] rd_resp_desc_2_xuser_10_reg
			       ,input [31:0] rd_resp_desc_2_xuser_11_reg
			       ,input [31:0] rd_resp_desc_2_xuser_12_reg
			       ,input [31:0] rd_resp_desc_2_xuser_13_reg
			       ,input [31:0] rd_resp_desc_2_xuser_14_reg
			       ,input [31:0] rd_resp_desc_2_xuser_15_reg
			       ,input [31:0] wr_req_desc_2_txn_type_reg
			       ,input [31:0] wr_req_desc_2_size_reg
			       ,input [31:0] wr_req_desc_2_data_offset_reg
			       ,input [31:0] wr_req_desc_2_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_2_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_2_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_2_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_2_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_2_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_2_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_2_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_2_axsize_reg
			       ,input [31:0] wr_req_desc_2_attr_reg
			       ,input [31:0] wr_req_desc_2_axaddr_0_reg
			       ,input [31:0] wr_req_desc_2_axaddr_1_reg
			       ,input [31:0] wr_req_desc_2_axaddr_2_reg
			       ,input [31:0] wr_req_desc_2_axaddr_3_reg
			       ,input [31:0] wr_req_desc_2_axid_0_reg
			       ,input [31:0] wr_req_desc_2_axid_1_reg
			       ,input [31:0] wr_req_desc_2_axid_2_reg
			       ,input [31:0] wr_req_desc_2_axid_3_reg
			       ,input [31:0] wr_req_desc_2_axuser_0_reg
			       ,input [31:0] wr_req_desc_2_axuser_1_reg
			       ,input [31:0] wr_req_desc_2_axuser_2_reg
			       ,input [31:0] wr_req_desc_2_axuser_3_reg
			       ,input [31:0] wr_req_desc_2_axuser_4_reg
			       ,input [31:0] wr_req_desc_2_axuser_5_reg
			       ,input [31:0] wr_req_desc_2_axuser_6_reg
			       ,input [31:0] wr_req_desc_2_axuser_7_reg
			       ,input [31:0] wr_req_desc_2_axuser_8_reg
			       ,input [31:0] wr_req_desc_2_axuser_9_reg
			       ,input [31:0] wr_req_desc_2_axuser_10_reg
			       ,input [31:0] wr_req_desc_2_axuser_11_reg
			       ,input [31:0] wr_req_desc_2_axuser_12_reg
			       ,input [31:0] wr_req_desc_2_axuser_13_reg
			       ,input [31:0] wr_req_desc_2_axuser_14_reg
			       ,input [31:0] wr_req_desc_2_axuser_15_reg
			       ,input [31:0] wr_req_desc_2_wuser_0_reg
			       ,input [31:0] wr_req_desc_2_wuser_1_reg
			       ,input [31:0] wr_req_desc_2_wuser_2_reg
			       ,input [31:0] wr_req_desc_2_wuser_3_reg
			       ,input [31:0] wr_req_desc_2_wuser_4_reg
			       ,input [31:0] wr_req_desc_2_wuser_5_reg
			       ,input [31:0] wr_req_desc_2_wuser_6_reg
			       ,input [31:0] wr_req_desc_2_wuser_7_reg
			       ,input [31:0] wr_req_desc_2_wuser_8_reg
			       ,input [31:0] wr_req_desc_2_wuser_9_reg
			       ,input [31:0] wr_req_desc_2_wuser_10_reg
			       ,input [31:0] wr_req_desc_2_wuser_11_reg
			       ,input [31:0] wr_req_desc_2_wuser_12_reg
			       ,input [31:0] wr_req_desc_2_wuser_13_reg
			       ,input [31:0] wr_req_desc_2_wuser_14_reg
			       ,input [31:0] wr_req_desc_2_wuser_15_reg
			       ,input [31:0] wr_resp_desc_2_resp_reg
			       ,input [31:0] wr_resp_desc_2_xid_0_reg
			       ,input [31:0] wr_resp_desc_2_xid_1_reg
			       ,input [31:0] wr_resp_desc_2_xid_2_reg
			       ,input [31:0] wr_resp_desc_2_xid_3_reg
			       ,input [31:0] wr_resp_desc_2_xuser_0_reg
			       ,input [31:0] wr_resp_desc_2_xuser_1_reg
			       ,input [31:0] wr_resp_desc_2_xuser_2_reg
			       ,input [31:0] wr_resp_desc_2_xuser_3_reg
			       ,input [31:0] wr_resp_desc_2_xuser_4_reg
			       ,input [31:0] wr_resp_desc_2_xuser_5_reg
			       ,input [31:0] wr_resp_desc_2_xuser_6_reg
			       ,input [31:0] wr_resp_desc_2_xuser_7_reg
			       ,input [31:0] wr_resp_desc_2_xuser_8_reg
			       ,input [31:0] wr_resp_desc_2_xuser_9_reg
			       ,input [31:0] wr_resp_desc_2_xuser_10_reg
			       ,input [31:0] wr_resp_desc_2_xuser_11_reg
			       ,input [31:0] wr_resp_desc_2_xuser_12_reg
			       ,input [31:0] wr_resp_desc_2_xuser_13_reg
			       ,input [31:0] wr_resp_desc_2_xuser_14_reg
			       ,input [31:0] wr_resp_desc_2_xuser_15_reg
			       ,input [31:0] sn_req_desc_2_attr_reg
			       ,input [31:0] sn_req_desc_2_acaddr_0_reg
			       ,input [31:0] sn_req_desc_2_acaddr_1_reg
			       ,input [31:0] sn_req_desc_2_acaddr_2_reg
			       ,input [31:0] sn_req_desc_2_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_2_resp_reg
			       ,input [31:0] rd_req_desc_3_txn_type_reg
			       ,input [31:0] rd_req_desc_3_size_reg
			       ,input [31:0] rd_req_desc_3_axsize_reg
			       ,input [31:0] rd_req_desc_3_attr_reg
			       ,input [31:0] rd_req_desc_3_axaddr_0_reg
			       ,input [31:0] rd_req_desc_3_axaddr_1_reg
			       ,input [31:0] rd_req_desc_3_axaddr_2_reg
			       ,input [31:0] rd_req_desc_3_axaddr_3_reg
			       ,input [31:0] rd_req_desc_3_axid_0_reg
			       ,input [31:0] rd_req_desc_3_axid_1_reg
			       ,input [31:0] rd_req_desc_3_axid_2_reg
			       ,input [31:0] rd_req_desc_3_axid_3_reg
			       ,input [31:0] rd_req_desc_3_axuser_0_reg
			       ,input [31:0] rd_req_desc_3_axuser_1_reg
			       ,input [31:0] rd_req_desc_3_axuser_2_reg
			       ,input [31:0] rd_req_desc_3_axuser_3_reg
			       ,input [31:0] rd_req_desc_3_axuser_4_reg
			       ,input [31:0] rd_req_desc_3_axuser_5_reg
			       ,input [31:0] rd_req_desc_3_axuser_6_reg
			       ,input [31:0] rd_req_desc_3_axuser_7_reg
			       ,input [31:0] rd_req_desc_3_axuser_8_reg
			       ,input [31:0] rd_req_desc_3_axuser_9_reg
			       ,input [31:0] rd_req_desc_3_axuser_10_reg
			       ,input [31:0] rd_req_desc_3_axuser_11_reg
			       ,input [31:0] rd_req_desc_3_axuser_12_reg
			       ,input [31:0] rd_req_desc_3_axuser_13_reg
			       ,input [31:0] rd_req_desc_3_axuser_14_reg
			       ,input [31:0] rd_req_desc_3_axuser_15_reg
			       ,input [31:0] rd_resp_desc_3_data_offset_reg
			       ,input [31:0] rd_resp_desc_3_data_size_reg
			       ,input [31:0] rd_resp_desc_3_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_3_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_3_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_3_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_3_resp_reg
			       ,input [31:0] rd_resp_desc_3_xid_0_reg
			       ,input [31:0] rd_resp_desc_3_xid_1_reg
			       ,input [31:0] rd_resp_desc_3_xid_2_reg
			       ,input [31:0] rd_resp_desc_3_xid_3_reg
			       ,input [31:0] rd_resp_desc_3_xuser_0_reg
			       ,input [31:0] rd_resp_desc_3_xuser_1_reg
			       ,input [31:0] rd_resp_desc_3_xuser_2_reg
			       ,input [31:0] rd_resp_desc_3_xuser_3_reg
			       ,input [31:0] rd_resp_desc_3_xuser_4_reg
			       ,input [31:0] rd_resp_desc_3_xuser_5_reg
			       ,input [31:0] rd_resp_desc_3_xuser_6_reg
			       ,input [31:0] rd_resp_desc_3_xuser_7_reg
			       ,input [31:0] rd_resp_desc_3_xuser_8_reg
			       ,input [31:0] rd_resp_desc_3_xuser_9_reg
			       ,input [31:0] rd_resp_desc_3_xuser_10_reg
			       ,input [31:0] rd_resp_desc_3_xuser_11_reg
			       ,input [31:0] rd_resp_desc_3_xuser_12_reg
			       ,input [31:0] rd_resp_desc_3_xuser_13_reg
			       ,input [31:0] rd_resp_desc_3_xuser_14_reg
			       ,input [31:0] rd_resp_desc_3_xuser_15_reg
			       ,input [31:0] wr_req_desc_3_txn_type_reg
			       ,input [31:0] wr_req_desc_3_size_reg
			       ,input [31:0] wr_req_desc_3_data_offset_reg
			       ,input [31:0] wr_req_desc_3_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_3_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_3_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_3_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_3_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_3_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_3_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_3_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_3_axsize_reg
			       ,input [31:0] wr_req_desc_3_attr_reg
			       ,input [31:0] wr_req_desc_3_axaddr_0_reg
			       ,input [31:0] wr_req_desc_3_axaddr_1_reg
			       ,input [31:0] wr_req_desc_3_axaddr_2_reg
			       ,input [31:0] wr_req_desc_3_axaddr_3_reg
			       ,input [31:0] wr_req_desc_3_axid_0_reg
			       ,input [31:0] wr_req_desc_3_axid_1_reg
			       ,input [31:0] wr_req_desc_3_axid_2_reg
			       ,input [31:0] wr_req_desc_3_axid_3_reg
			       ,input [31:0] wr_req_desc_3_axuser_0_reg
			       ,input [31:0] wr_req_desc_3_axuser_1_reg
			       ,input [31:0] wr_req_desc_3_axuser_2_reg
			       ,input [31:0] wr_req_desc_3_axuser_3_reg
			       ,input [31:0] wr_req_desc_3_axuser_4_reg
			       ,input [31:0] wr_req_desc_3_axuser_5_reg
			       ,input [31:0] wr_req_desc_3_axuser_6_reg
			       ,input [31:0] wr_req_desc_3_axuser_7_reg
			       ,input [31:0] wr_req_desc_3_axuser_8_reg
			       ,input [31:0] wr_req_desc_3_axuser_9_reg
			       ,input [31:0] wr_req_desc_3_axuser_10_reg
			       ,input [31:0] wr_req_desc_3_axuser_11_reg
			       ,input [31:0] wr_req_desc_3_axuser_12_reg
			       ,input [31:0] wr_req_desc_3_axuser_13_reg
			       ,input [31:0] wr_req_desc_3_axuser_14_reg
			       ,input [31:0] wr_req_desc_3_axuser_15_reg
			       ,input [31:0] wr_req_desc_3_wuser_0_reg
			       ,input [31:0] wr_req_desc_3_wuser_1_reg
			       ,input [31:0] wr_req_desc_3_wuser_2_reg
			       ,input [31:0] wr_req_desc_3_wuser_3_reg
			       ,input [31:0] wr_req_desc_3_wuser_4_reg
			       ,input [31:0] wr_req_desc_3_wuser_5_reg
			       ,input [31:0] wr_req_desc_3_wuser_6_reg
			       ,input [31:0] wr_req_desc_3_wuser_7_reg
			       ,input [31:0] wr_req_desc_3_wuser_8_reg
			       ,input [31:0] wr_req_desc_3_wuser_9_reg
			       ,input [31:0] wr_req_desc_3_wuser_10_reg
			       ,input [31:0] wr_req_desc_3_wuser_11_reg
			       ,input [31:0] wr_req_desc_3_wuser_12_reg
			       ,input [31:0] wr_req_desc_3_wuser_13_reg
			       ,input [31:0] wr_req_desc_3_wuser_14_reg
			       ,input [31:0] wr_req_desc_3_wuser_15_reg
			       ,input [31:0] wr_resp_desc_3_resp_reg
			       ,input [31:0] wr_resp_desc_3_xid_0_reg
			       ,input [31:0] wr_resp_desc_3_xid_1_reg
			       ,input [31:0] wr_resp_desc_3_xid_2_reg
			       ,input [31:0] wr_resp_desc_3_xid_3_reg
			       ,input [31:0] wr_resp_desc_3_xuser_0_reg
			       ,input [31:0] wr_resp_desc_3_xuser_1_reg
			       ,input [31:0] wr_resp_desc_3_xuser_2_reg
			       ,input [31:0] wr_resp_desc_3_xuser_3_reg
			       ,input [31:0] wr_resp_desc_3_xuser_4_reg
			       ,input [31:0] wr_resp_desc_3_xuser_5_reg
			       ,input [31:0] wr_resp_desc_3_xuser_6_reg
			       ,input [31:0] wr_resp_desc_3_xuser_7_reg
			       ,input [31:0] wr_resp_desc_3_xuser_8_reg
			       ,input [31:0] wr_resp_desc_3_xuser_9_reg
			       ,input [31:0] wr_resp_desc_3_xuser_10_reg
			       ,input [31:0] wr_resp_desc_3_xuser_11_reg
			       ,input [31:0] wr_resp_desc_3_xuser_12_reg
			       ,input [31:0] wr_resp_desc_3_xuser_13_reg
			       ,input [31:0] wr_resp_desc_3_xuser_14_reg
			       ,input [31:0] wr_resp_desc_3_xuser_15_reg
			       ,input [31:0] sn_req_desc_3_attr_reg
			       ,input [31:0] sn_req_desc_3_acaddr_0_reg
			       ,input [31:0] sn_req_desc_3_acaddr_1_reg
			       ,input [31:0] sn_req_desc_3_acaddr_2_reg
			       ,input [31:0] sn_req_desc_3_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_3_resp_reg
			       ,input [31:0] rd_req_desc_4_txn_type_reg
			       ,input [31:0] rd_req_desc_4_size_reg
			       ,input [31:0] rd_req_desc_4_axsize_reg
			       ,input [31:0] rd_req_desc_4_attr_reg
			       ,input [31:0] rd_req_desc_4_axaddr_0_reg
			       ,input [31:0] rd_req_desc_4_axaddr_1_reg
			       ,input [31:0] rd_req_desc_4_axaddr_2_reg
			       ,input [31:0] rd_req_desc_4_axaddr_3_reg
			       ,input [31:0] rd_req_desc_4_axid_0_reg
			       ,input [31:0] rd_req_desc_4_axid_1_reg
			       ,input [31:0] rd_req_desc_4_axid_2_reg
			       ,input [31:0] rd_req_desc_4_axid_3_reg
			       ,input [31:0] rd_req_desc_4_axuser_0_reg
			       ,input [31:0] rd_req_desc_4_axuser_1_reg
			       ,input [31:0] rd_req_desc_4_axuser_2_reg
			       ,input [31:0] rd_req_desc_4_axuser_3_reg
			       ,input [31:0] rd_req_desc_4_axuser_4_reg
			       ,input [31:0] rd_req_desc_4_axuser_5_reg
			       ,input [31:0] rd_req_desc_4_axuser_6_reg
			       ,input [31:0] rd_req_desc_4_axuser_7_reg
			       ,input [31:0] rd_req_desc_4_axuser_8_reg
			       ,input [31:0] rd_req_desc_4_axuser_9_reg
			       ,input [31:0] rd_req_desc_4_axuser_10_reg
			       ,input [31:0] rd_req_desc_4_axuser_11_reg
			       ,input [31:0] rd_req_desc_4_axuser_12_reg
			       ,input [31:0] rd_req_desc_4_axuser_13_reg
			       ,input [31:0] rd_req_desc_4_axuser_14_reg
			       ,input [31:0] rd_req_desc_4_axuser_15_reg
			       ,input [31:0] rd_resp_desc_4_data_offset_reg
			       ,input [31:0] rd_resp_desc_4_data_size_reg
			       ,input [31:0] rd_resp_desc_4_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_4_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_4_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_4_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_4_resp_reg
			       ,input [31:0] rd_resp_desc_4_xid_0_reg
			       ,input [31:0] rd_resp_desc_4_xid_1_reg
			       ,input [31:0] rd_resp_desc_4_xid_2_reg
			       ,input [31:0] rd_resp_desc_4_xid_3_reg
			       ,input [31:0] rd_resp_desc_4_xuser_0_reg
			       ,input [31:0] rd_resp_desc_4_xuser_1_reg
			       ,input [31:0] rd_resp_desc_4_xuser_2_reg
			       ,input [31:0] rd_resp_desc_4_xuser_3_reg
			       ,input [31:0] rd_resp_desc_4_xuser_4_reg
			       ,input [31:0] rd_resp_desc_4_xuser_5_reg
			       ,input [31:0] rd_resp_desc_4_xuser_6_reg
			       ,input [31:0] rd_resp_desc_4_xuser_7_reg
			       ,input [31:0] rd_resp_desc_4_xuser_8_reg
			       ,input [31:0] rd_resp_desc_4_xuser_9_reg
			       ,input [31:0] rd_resp_desc_4_xuser_10_reg
			       ,input [31:0] rd_resp_desc_4_xuser_11_reg
			       ,input [31:0] rd_resp_desc_4_xuser_12_reg
			       ,input [31:0] rd_resp_desc_4_xuser_13_reg
			       ,input [31:0] rd_resp_desc_4_xuser_14_reg
			       ,input [31:0] rd_resp_desc_4_xuser_15_reg
			       ,input [31:0] wr_req_desc_4_txn_type_reg
			       ,input [31:0] wr_req_desc_4_size_reg
			       ,input [31:0] wr_req_desc_4_data_offset_reg
			       ,input [31:0] wr_req_desc_4_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_4_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_4_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_4_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_4_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_4_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_4_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_4_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_4_axsize_reg
			       ,input [31:0] wr_req_desc_4_attr_reg
			       ,input [31:0] wr_req_desc_4_axaddr_0_reg
			       ,input [31:0] wr_req_desc_4_axaddr_1_reg
			       ,input [31:0] wr_req_desc_4_axaddr_2_reg
			       ,input [31:0] wr_req_desc_4_axaddr_3_reg
			       ,input [31:0] wr_req_desc_4_axid_0_reg
			       ,input [31:0] wr_req_desc_4_axid_1_reg
			       ,input [31:0] wr_req_desc_4_axid_2_reg
			       ,input [31:0] wr_req_desc_4_axid_3_reg
			       ,input [31:0] wr_req_desc_4_axuser_0_reg
			       ,input [31:0] wr_req_desc_4_axuser_1_reg
			       ,input [31:0] wr_req_desc_4_axuser_2_reg
			       ,input [31:0] wr_req_desc_4_axuser_3_reg
			       ,input [31:0] wr_req_desc_4_axuser_4_reg
			       ,input [31:0] wr_req_desc_4_axuser_5_reg
			       ,input [31:0] wr_req_desc_4_axuser_6_reg
			       ,input [31:0] wr_req_desc_4_axuser_7_reg
			       ,input [31:0] wr_req_desc_4_axuser_8_reg
			       ,input [31:0] wr_req_desc_4_axuser_9_reg
			       ,input [31:0] wr_req_desc_4_axuser_10_reg
			       ,input [31:0] wr_req_desc_4_axuser_11_reg
			       ,input [31:0] wr_req_desc_4_axuser_12_reg
			       ,input [31:0] wr_req_desc_4_axuser_13_reg
			       ,input [31:0] wr_req_desc_4_axuser_14_reg
			       ,input [31:0] wr_req_desc_4_axuser_15_reg
			       ,input [31:0] wr_req_desc_4_wuser_0_reg
			       ,input [31:0] wr_req_desc_4_wuser_1_reg
			       ,input [31:0] wr_req_desc_4_wuser_2_reg
			       ,input [31:0] wr_req_desc_4_wuser_3_reg
			       ,input [31:0] wr_req_desc_4_wuser_4_reg
			       ,input [31:0] wr_req_desc_4_wuser_5_reg
			       ,input [31:0] wr_req_desc_4_wuser_6_reg
			       ,input [31:0] wr_req_desc_4_wuser_7_reg
			       ,input [31:0] wr_req_desc_4_wuser_8_reg
			       ,input [31:0] wr_req_desc_4_wuser_9_reg
			       ,input [31:0] wr_req_desc_4_wuser_10_reg
			       ,input [31:0] wr_req_desc_4_wuser_11_reg
			       ,input [31:0] wr_req_desc_4_wuser_12_reg
			       ,input [31:0] wr_req_desc_4_wuser_13_reg
			       ,input [31:0] wr_req_desc_4_wuser_14_reg
			       ,input [31:0] wr_req_desc_4_wuser_15_reg
			       ,input [31:0] wr_resp_desc_4_resp_reg
			       ,input [31:0] wr_resp_desc_4_xid_0_reg
			       ,input [31:0] wr_resp_desc_4_xid_1_reg
			       ,input [31:0] wr_resp_desc_4_xid_2_reg
			       ,input [31:0] wr_resp_desc_4_xid_3_reg
			       ,input [31:0] wr_resp_desc_4_xuser_0_reg
			       ,input [31:0] wr_resp_desc_4_xuser_1_reg
			       ,input [31:0] wr_resp_desc_4_xuser_2_reg
			       ,input [31:0] wr_resp_desc_4_xuser_3_reg
			       ,input [31:0] wr_resp_desc_4_xuser_4_reg
			       ,input [31:0] wr_resp_desc_4_xuser_5_reg
			       ,input [31:0] wr_resp_desc_4_xuser_6_reg
			       ,input [31:0] wr_resp_desc_4_xuser_7_reg
			       ,input [31:0] wr_resp_desc_4_xuser_8_reg
			       ,input [31:0] wr_resp_desc_4_xuser_9_reg
			       ,input [31:0] wr_resp_desc_4_xuser_10_reg
			       ,input [31:0] wr_resp_desc_4_xuser_11_reg
			       ,input [31:0] wr_resp_desc_4_xuser_12_reg
			       ,input [31:0] wr_resp_desc_4_xuser_13_reg
			       ,input [31:0] wr_resp_desc_4_xuser_14_reg
			       ,input [31:0] wr_resp_desc_4_xuser_15_reg
			       ,input [31:0] sn_req_desc_4_attr_reg
			       ,input [31:0] sn_req_desc_4_acaddr_0_reg
			       ,input [31:0] sn_req_desc_4_acaddr_1_reg
			       ,input [31:0] sn_req_desc_4_acaddr_2_reg
			       ,input [31:0] sn_req_desc_4_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_4_resp_reg
			       ,input [31:0] rd_req_desc_5_txn_type_reg
			       ,input [31:0] rd_req_desc_5_size_reg
			       ,input [31:0] rd_req_desc_5_axsize_reg
			       ,input [31:0] rd_req_desc_5_attr_reg
			       ,input [31:0] rd_req_desc_5_axaddr_0_reg
			       ,input [31:0] rd_req_desc_5_axaddr_1_reg
			       ,input [31:0] rd_req_desc_5_axaddr_2_reg
			       ,input [31:0] rd_req_desc_5_axaddr_3_reg
			       ,input [31:0] rd_req_desc_5_axid_0_reg
			       ,input [31:0] rd_req_desc_5_axid_1_reg
			       ,input [31:0] rd_req_desc_5_axid_2_reg
			       ,input [31:0] rd_req_desc_5_axid_3_reg
			       ,input [31:0] rd_req_desc_5_axuser_0_reg
			       ,input [31:0] rd_req_desc_5_axuser_1_reg
			       ,input [31:0] rd_req_desc_5_axuser_2_reg
			       ,input [31:0] rd_req_desc_5_axuser_3_reg
			       ,input [31:0] rd_req_desc_5_axuser_4_reg
			       ,input [31:0] rd_req_desc_5_axuser_5_reg
			       ,input [31:0] rd_req_desc_5_axuser_6_reg
			       ,input [31:0] rd_req_desc_5_axuser_7_reg
			       ,input [31:0] rd_req_desc_5_axuser_8_reg
			       ,input [31:0] rd_req_desc_5_axuser_9_reg
			       ,input [31:0] rd_req_desc_5_axuser_10_reg
			       ,input [31:0] rd_req_desc_5_axuser_11_reg
			       ,input [31:0] rd_req_desc_5_axuser_12_reg
			       ,input [31:0] rd_req_desc_5_axuser_13_reg
			       ,input [31:0] rd_req_desc_5_axuser_14_reg
			       ,input [31:0] rd_req_desc_5_axuser_15_reg
			       ,input [31:0] rd_resp_desc_5_data_offset_reg
			       ,input [31:0] rd_resp_desc_5_data_size_reg
			       ,input [31:0] rd_resp_desc_5_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_5_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_5_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_5_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_5_resp_reg
			       ,input [31:0] rd_resp_desc_5_xid_0_reg
			       ,input [31:0] rd_resp_desc_5_xid_1_reg
			       ,input [31:0] rd_resp_desc_5_xid_2_reg
			       ,input [31:0] rd_resp_desc_5_xid_3_reg
			       ,input [31:0] rd_resp_desc_5_xuser_0_reg
			       ,input [31:0] rd_resp_desc_5_xuser_1_reg
			       ,input [31:0] rd_resp_desc_5_xuser_2_reg
			       ,input [31:0] rd_resp_desc_5_xuser_3_reg
			       ,input [31:0] rd_resp_desc_5_xuser_4_reg
			       ,input [31:0] rd_resp_desc_5_xuser_5_reg
			       ,input [31:0] rd_resp_desc_5_xuser_6_reg
			       ,input [31:0] rd_resp_desc_5_xuser_7_reg
			       ,input [31:0] rd_resp_desc_5_xuser_8_reg
			       ,input [31:0] rd_resp_desc_5_xuser_9_reg
			       ,input [31:0] rd_resp_desc_5_xuser_10_reg
			       ,input [31:0] rd_resp_desc_5_xuser_11_reg
			       ,input [31:0] rd_resp_desc_5_xuser_12_reg
			       ,input [31:0] rd_resp_desc_5_xuser_13_reg
			       ,input [31:0] rd_resp_desc_5_xuser_14_reg
			       ,input [31:0] rd_resp_desc_5_xuser_15_reg
			       ,input [31:0] wr_req_desc_5_txn_type_reg
			       ,input [31:0] wr_req_desc_5_size_reg
			       ,input [31:0] wr_req_desc_5_data_offset_reg
			       ,input [31:0] wr_req_desc_5_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_5_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_5_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_5_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_5_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_5_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_5_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_5_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_5_axsize_reg
			       ,input [31:0] wr_req_desc_5_attr_reg
			       ,input [31:0] wr_req_desc_5_axaddr_0_reg
			       ,input [31:0] wr_req_desc_5_axaddr_1_reg
			       ,input [31:0] wr_req_desc_5_axaddr_2_reg
			       ,input [31:0] wr_req_desc_5_axaddr_3_reg
			       ,input [31:0] wr_req_desc_5_axid_0_reg
			       ,input [31:0] wr_req_desc_5_axid_1_reg
			       ,input [31:0] wr_req_desc_5_axid_2_reg
			       ,input [31:0] wr_req_desc_5_axid_3_reg
			       ,input [31:0] wr_req_desc_5_axuser_0_reg
			       ,input [31:0] wr_req_desc_5_axuser_1_reg
			       ,input [31:0] wr_req_desc_5_axuser_2_reg
			       ,input [31:0] wr_req_desc_5_axuser_3_reg
			       ,input [31:0] wr_req_desc_5_axuser_4_reg
			       ,input [31:0] wr_req_desc_5_axuser_5_reg
			       ,input [31:0] wr_req_desc_5_axuser_6_reg
			       ,input [31:0] wr_req_desc_5_axuser_7_reg
			       ,input [31:0] wr_req_desc_5_axuser_8_reg
			       ,input [31:0] wr_req_desc_5_axuser_9_reg
			       ,input [31:0] wr_req_desc_5_axuser_10_reg
			       ,input [31:0] wr_req_desc_5_axuser_11_reg
			       ,input [31:0] wr_req_desc_5_axuser_12_reg
			       ,input [31:0] wr_req_desc_5_axuser_13_reg
			       ,input [31:0] wr_req_desc_5_axuser_14_reg
			       ,input [31:0] wr_req_desc_5_axuser_15_reg
			       ,input [31:0] wr_req_desc_5_wuser_0_reg
			       ,input [31:0] wr_req_desc_5_wuser_1_reg
			       ,input [31:0] wr_req_desc_5_wuser_2_reg
			       ,input [31:0] wr_req_desc_5_wuser_3_reg
			       ,input [31:0] wr_req_desc_5_wuser_4_reg
			       ,input [31:0] wr_req_desc_5_wuser_5_reg
			       ,input [31:0] wr_req_desc_5_wuser_6_reg
			       ,input [31:0] wr_req_desc_5_wuser_7_reg
			       ,input [31:0] wr_req_desc_5_wuser_8_reg
			       ,input [31:0] wr_req_desc_5_wuser_9_reg
			       ,input [31:0] wr_req_desc_5_wuser_10_reg
			       ,input [31:0] wr_req_desc_5_wuser_11_reg
			       ,input [31:0] wr_req_desc_5_wuser_12_reg
			       ,input [31:0] wr_req_desc_5_wuser_13_reg
			       ,input [31:0] wr_req_desc_5_wuser_14_reg
			       ,input [31:0] wr_req_desc_5_wuser_15_reg
			       ,input [31:0] wr_resp_desc_5_resp_reg
			       ,input [31:0] wr_resp_desc_5_xid_0_reg
			       ,input [31:0] wr_resp_desc_5_xid_1_reg
			       ,input [31:0] wr_resp_desc_5_xid_2_reg
			       ,input [31:0] wr_resp_desc_5_xid_3_reg
			       ,input [31:0] wr_resp_desc_5_xuser_0_reg
			       ,input [31:0] wr_resp_desc_5_xuser_1_reg
			       ,input [31:0] wr_resp_desc_5_xuser_2_reg
			       ,input [31:0] wr_resp_desc_5_xuser_3_reg
			       ,input [31:0] wr_resp_desc_5_xuser_4_reg
			       ,input [31:0] wr_resp_desc_5_xuser_5_reg
			       ,input [31:0] wr_resp_desc_5_xuser_6_reg
			       ,input [31:0] wr_resp_desc_5_xuser_7_reg
			       ,input [31:0] wr_resp_desc_5_xuser_8_reg
			       ,input [31:0] wr_resp_desc_5_xuser_9_reg
			       ,input [31:0] wr_resp_desc_5_xuser_10_reg
			       ,input [31:0] wr_resp_desc_5_xuser_11_reg
			       ,input [31:0] wr_resp_desc_5_xuser_12_reg
			       ,input [31:0] wr_resp_desc_5_xuser_13_reg
			       ,input [31:0] wr_resp_desc_5_xuser_14_reg
			       ,input [31:0] wr_resp_desc_5_xuser_15_reg
			       ,input [31:0] sn_req_desc_5_attr_reg
			       ,input [31:0] sn_req_desc_5_acaddr_0_reg
			       ,input [31:0] sn_req_desc_5_acaddr_1_reg
			       ,input [31:0] sn_req_desc_5_acaddr_2_reg
			       ,input [31:0] sn_req_desc_5_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_5_resp_reg
			       ,input [31:0] rd_req_desc_6_txn_type_reg
			       ,input [31:0] rd_req_desc_6_size_reg
			       ,input [31:0] rd_req_desc_6_axsize_reg
			       ,input [31:0] rd_req_desc_6_attr_reg
			       ,input [31:0] rd_req_desc_6_axaddr_0_reg
			       ,input [31:0] rd_req_desc_6_axaddr_1_reg
			       ,input [31:0] rd_req_desc_6_axaddr_2_reg
			       ,input [31:0] rd_req_desc_6_axaddr_3_reg
			       ,input [31:0] rd_req_desc_6_axid_0_reg
			       ,input [31:0] rd_req_desc_6_axid_1_reg
			       ,input [31:0] rd_req_desc_6_axid_2_reg
			       ,input [31:0] rd_req_desc_6_axid_3_reg
			       ,input [31:0] rd_req_desc_6_axuser_0_reg
			       ,input [31:0] rd_req_desc_6_axuser_1_reg
			       ,input [31:0] rd_req_desc_6_axuser_2_reg
			       ,input [31:0] rd_req_desc_6_axuser_3_reg
			       ,input [31:0] rd_req_desc_6_axuser_4_reg
			       ,input [31:0] rd_req_desc_6_axuser_5_reg
			       ,input [31:0] rd_req_desc_6_axuser_6_reg
			       ,input [31:0] rd_req_desc_6_axuser_7_reg
			       ,input [31:0] rd_req_desc_6_axuser_8_reg
			       ,input [31:0] rd_req_desc_6_axuser_9_reg
			       ,input [31:0] rd_req_desc_6_axuser_10_reg
			       ,input [31:0] rd_req_desc_6_axuser_11_reg
			       ,input [31:0] rd_req_desc_6_axuser_12_reg
			       ,input [31:0] rd_req_desc_6_axuser_13_reg
			       ,input [31:0] rd_req_desc_6_axuser_14_reg
			       ,input [31:0] rd_req_desc_6_axuser_15_reg
			       ,input [31:0] rd_resp_desc_6_data_offset_reg
			       ,input [31:0] rd_resp_desc_6_data_size_reg
			       ,input [31:0] rd_resp_desc_6_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_6_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_6_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_6_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_6_resp_reg
			       ,input [31:0] rd_resp_desc_6_xid_0_reg
			       ,input [31:0] rd_resp_desc_6_xid_1_reg
			       ,input [31:0] rd_resp_desc_6_xid_2_reg
			       ,input [31:0] rd_resp_desc_6_xid_3_reg
			       ,input [31:0] rd_resp_desc_6_xuser_0_reg
			       ,input [31:0] rd_resp_desc_6_xuser_1_reg
			       ,input [31:0] rd_resp_desc_6_xuser_2_reg
			       ,input [31:0] rd_resp_desc_6_xuser_3_reg
			       ,input [31:0] rd_resp_desc_6_xuser_4_reg
			       ,input [31:0] rd_resp_desc_6_xuser_5_reg
			       ,input [31:0] rd_resp_desc_6_xuser_6_reg
			       ,input [31:0] rd_resp_desc_6_xuser_7_reg
			       ,input [31:0] rd_resp_desc_6_xuser_8_reg
			       ,input [31:0] rd_resp_desc_6_xuser_9_reg
			       ,input [31:0] rd_resp_desc_6_xuser_10_reg
			       ,input [31:0] rd_resp_desc_6_xuser_11_reg
			       ,input [31:0] rd_resp_desc_6_xuser_12_reg
			       ,input [31:0] rd_resp_desc_6_xuser_13_reg
			       ,input [31:0] rd_resp_desc_6_xuser_14_reg
			       ,input [31:0] rd_resp_desc_6_xuser_15_reg
			       ,input [31:0] wr_req_desc_6_txn_type_reg
			       ,input [31:0] wr_req_desc_6_size_reg
			       ,input [31:0] wr_req_desc_6_data_offset_reg
			       ,input [31:0] wr_req_desc_6_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_6_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_6_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_6_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_6_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_6_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_6_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_6_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_6_axsize_reg
			       ,input [31:0] wr_req_desc_6_attr_reg
			       ,input [31:0] wr_req_desc_6_axaddr_0_reg
			       ,input [31:0] wr_req_desc_6_axaddr_1_reg
			       ,input [31:0] wr_req_desc_6_axaddr_2_reg
			       ,input [31:0] wr_req_desc_6_axaddr_3_reg
			       ,input [31:0] wr_req_desc_6_axid_0_reg
			       ,input [31:0] wr_req_desc_6_axid_1_reg
			       ,input [31:0] wr_req_desc_6_axid_2_reg
			       ,input [31:0] wr_req_desc_6_axid_3_reg
			       ,input [31:0] wr_req_desc_6_axuser_0_reg
			       ,input [31:0] wr_req_desc_6_axuser_1_reg
			       ,input [31:0] wr_req_desc_6_axuser_2_reg
			       ,input [31:0] wr_req_desc_6_axuser_3_reg
			       ,input [31:0] wr_req_desc_6_axuser_4_reg
			       ,input [31:0] wr_req_desc_6_axuser_5_reg
			       ,input [31:0] wr_req_desc_6_axuser_6_reg
			       ,input [31:0] wr_req_desc_6_axuser_7_reg
			       ,input [31:0] wr_req_desc_6_axuser_8_reg
			       ,input [31:0] wr_req_desc_6_axuser_9_reg
			       ,input [31:0] wr_req_desc_6_axuser_10_reg
			       ,input [31:0] wr_req_desc_6_axuser_11_reg
			       ,input [31:0] wr_req_desc_6_axuser_12_reg
			       ,input [31:0] wr_req_desc_6_axuser_13_reg
			       ,input [31:0] wr_req_desc_6_axuser_14_reg
			       ,input [31:0] wr_req_desc_6_axuser_15_reg
			       ,input [31:0] wr_req_desc_6_wuser_0_reg
			       ,input [31:0] wr_req_desc_6_wuser_1_reg
			       ,input [31:0] wr_req_desc_6_wuser_2_reg
			       ,input [31:0] wr_req_desc_6_wuser_3_reg
			       ,input [31:0] wr_req_desc_6_wuser_4_reg
			       ,input [31:0] wr_req_desc_6_wuser_5_reg
			       ,input [31:0] wr_req_desc_6_wuser_6_reg
			       ,input [31:0] wr_req_desc_6_wuser_7_reg
			       ,input [31:0] wr_req_desc_6_wuser_8_reg
			       ,input [31:0] wr_req_desc_6_wuser_9_reg
			       ,input [31:0] wr_req_desc_6_wuser_10_reg
			       ,input [31:0] wr_req_desc_6_wuser_11_reg
			       ,input [31:0] wr_req_desc_6_wuser_12_reg
			       ,input [31:0] wr_req_desc_6_wuser_13_reg
			       ,input [31:0] wr_req_desc_6_wuser_14_reg
			       ,input [31:0] wr_req_desc_6_wuser_15_reg
			       ,input [31:0] wr_resp_desc_6_resp_reg
			       ,input [31:0] wr_resp_desc_6_xid_0_reg
			       ,input [31:0] wr_resp_desc_6_xid_1_reg
			       ,input [31:0] wr_resp_desc_6_xid_2_reg
			       ,input [31:0] wr_resp_desc_6_xid_3_reg
			       ,input [31:0] wr_resp_desc_6_xuser_0_reg
			       ,input [31:0] wr_resp_desc_6_xuser_1_reg
			       ,input [31:0] wr_resp_desc_6_xuser_2_reg
			       ,input [31:0] wr_resp_desc_6_xuser_3_reg
			       ,input [31:0] wr_resp_desc_6_xuser_4_reg
			       ,input [31:0] wr_resp_desc_6_xuser_5_reg
			       ,input [31:0] wr_resp_desc_6_xuser_6_reg
			       ,input [31:0] wr_resp_desc_6_xuser_7_reg
			       ,input [31:0] wr_resp_desc_6_xuser_8_reg
			       ,input [31:0] wr_resp_desc_6_xuser_9_reg
			       ,input [31:0] wr_resp_desc_6_xuser_10_reg
			       ,input [31:0] wr_resp_desc_6_xuser_11_reg
			       ,input [31:0] wr_resp_desc_6_xuser_12_reg
			       ,input [31:0] wr_resp_desc_6_xuser_13_reg
			       ,input [31:0] wr_resp_desc_6_xuser_14_reg
			       ,input [31:0] wr_resp_desc_6_xuser_15_reg
			       ,input [31:0] sn_req_desc_6_attr_reg
			       ,input [31:0] sn_req_desc_6_acaddr_0_reg
			       ,input [31:0] sn_req_desc_6_acaddr_1_reg
			       ,input [31:0] sn_req_desc_6_acaddr_2_reg
			       ,input [31:0] sn_req_desc_6_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_6_resp_reg
			       ,input [31:0] rd_req_desc_7_txn_type_reg
			       ,input [31:0] rd_req_desc_7_size_reg
			       ,input [31:0] rd_req_desc_7_axsize_reg
			       ,input [31:0] rd_req_desc_7_attr_reg
			       ,input [31:0] rd_req_desc_7_axaddr_0_reg
			       ,input [31:0] rd_req_desc_7_axaddr_1_reg
			       ,input [31:0] rd_req_desc_7_axaddr_2_reg
			       ,input [31:0] rd_req_desc_7_axaddr_3_reg
			       ,input [31:0] rd_req_desc_7_axid_0_reg
			       ,input [31:0] rd_req_desc_7_axid_1_reg
			       ,input [31:0] rd_req_desc_7_axid_2_reg
			       ,input [31:0] rd_req_desc_7_axid_3_reg
			       ,input [31:0] rd_req_desc_7_axuser_0_reg
			       ,input [31:0] rd_req_desc_7_axuser_1_reg
			       ,input [31:0] rd_req_desc_7_axuser_2_reg
			       ,input [31:0] rd_req_desc_7_axuser_3_reg
			       ,input [31:0] rd_req_desc_7_axuser_4_reg
			       ,input [31:0] rd_req_desc_7_axuser_5_reg
			       ,input [31:0] rd_req_desc_7_axuser_6_reg
			       ,input [31:0] rd_req_desc_7_axuser_7_reg
			       ,input [31:0] rd_req_desc_7_axuser_8_reg
			       ,input [31:0] rd_req_desc_7_axuser_9_reg
			       ,input [31:0] rd_req_desc_7_axuser_10_reg
			       ,input [31:0] rd_req_desc_7_axuser_11_reg
			       ,input [31:0] rd_req_desc_7_axuser_12_reg
			       ,input [31:0] rd_req_desc_7_axuser_13_reg
			       ,input [31:0] rd_req_desc_7_axuser_14_reg
			       ,input [31:0] rd_req_desc_7_axuser_15_reg
			       ,input [31:0] rd_resp_desc_7_data_offset_reg
			       ,input [31:0] rd_resp_desc_7_data_size_reg
			       ,input [31:0] rd_resp_desc_7_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_7_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_7_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_7_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_7_resp_reg
			       ,input [31:0] rd_resp_desc_7_xid_0_reg
			       ,input [31:0] rd_resp_desc_7_xid_1_reg
			       ,input [31:0] rd_resp_desc_7_xid_2_reg
			       ,input [31:0] rd_resp_desc_7_xid_3_reg
			       ,input [31:0] rd_resp_desc_7_xuser_0_reg
			       ,input [31:0] rd_resp_desc_7_xuser_1_reg
			       ,input [31:0] rd_resp_desc_7_xuser_2_reg
			       ,input [31:0] rd_resp_desc_7_xuser_3_reg
			       ,input [31:0] rd_resp_desc_7_xuser_4_reg
			       ,input [31:0] rd_resp_desc_7_xuser_5_reg
			       ,input [31:0] rd_resp_desc_7_xuser_6_reg
			       ,input [31:0] rd_resp_desc_7_xuser_7_reg
			       ,input [31:0] rd_resp_desc_7_xuser_8_reg
			       ,input [31:0] rd_resp_desc_7_xuser_9_reg
			       ,input [31:0] rd_resp_desc_7_xuser_10_reg
			       ,input [31:0] rd_resp_desc_7_xuser_11_reg
			       ,input [31:0] rd_resp_desc_7_xuser_12_reg
			       ,input [31:0] rd_resp_desc_7_xuser_13_reg
			       ,input [31:0] rd_resp_desc_7_xuser_14_reg
			       ,input [31:0] rd_resp_desc_7_xuser_15_reg
			       ,input [31:0] wr_req_desc_7_txn_type_reg
			       ,input [31:0] wr_req_desc_7_size_reg
			       ,input [31:0] wr_req_desc_7_data_offset_reg
			       ,input [31:0] wr_req_desc_7_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_7_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_7_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_7_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_7_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_7_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_7_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_7_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_7_axsize_reg
			       ,input [31:0] wr_req_desc_7_attr_reg
			       ,input [31:0] wr_req_desc_7_axaddr_0_reg
			       ,input [31:0] wr_req_desc_7_axaddr_1_reg
			       ,input [31:0] wr_req_desc_7_axaddr_2_reg
			       ,input [31:0] wr_req_desc_7_axaddr_3_reg
			       ,input [31:0] wr_req_desc_7_axid_0_reg
			       ,input [31:0] wr_req_desc_7_axid_1_reg
			       ,input [31:0] wr_req_desc_7_axid_2_reg
			       ,input [31:0] wr_req_desc_7_axid_3_reg
			       ,input [31:0] wr_req_desc_7_axuser_0_reg
			       ,input [31:0] wr_req_desc_7_axuser_1_reg
			       ,input [31:0] wr_req_desc_7_axuser_2_reg
			       ,input [31:0] wr_req_desc_7_axuser_3_reg
			       ,input [31:0] wr_req_desc_7_axuser_4_reg
			       ,input [31:0] wr_req_desc_7_axuser_5_reg
			       ,input [31:0] wr_req_desc_7_axuser_6_reg
			       ,input [31:0] wr_req_desc_7_axuser_7_reg
			       ,input [31:0] wr_req_desc_7_axuser_8_reg
			       ,input [31:0] wr_req_desc_7_axuser_9_reg
			       ,input [31:0] wr_req_desc_7_axuser_10_reg
			       ,input [31:0] wr_req_desc_7_axuser_11_reg
			       ,input [31:0] wr_req_desc_7_axuser_12_reg
			       ,input [31:0] wr_req_desc_7_axuser_13_reg
			       ,input [31:0] wr_req_desc_7_axuser_14_reg
			       ,input [31:0] wr_req_desc_7_axuser_15_reg
			       ,input [31:0] wr_req_desc_7_wuser_0_reg
			       ,input [31:0] wr_req_desc_7_wuser_1_reg
			       ,input [31:0] wr_req_desc_7_wuser_2_reg
			       ,input [31:0] wr_req_desc_7_wuser_3_reg
			       ,input [31:0] wr_req_desc_7_wuser_4_reg
			       ,input [31:0] wr_req_desc_7_wuser_5_reg
			       ,input [31:0] wr_req_desc_7_wuser_6_reg
			       ,input [31:0] wr_req_desc_7_wuser_7_reg
			       ,input [31:0] wr_req_desc_7_wuser_8_reg
			       ,input [31:0] wr_req_desc_7_wuser_9_reg
			       ,input [31:0] wr_req_desc_7_wuser_10_reg
			       ,input [31:0] wr_req_desc_7_wuser_11_reg
			       ,input [31:0] wr_req_desc_7_wuser_12_reg
			       ,input [31:0] wr_req_desc_7_wuser_13_reg
			       ,input [31:0] wr_req_desc_7_wuser_14_reg
			       ,input [31:0] wr_req_desc_7_wuser_15_reg
			       ,input [31:0] wr_resp_desc_7_resp_reg
			       ,input [31:0] wr_resp_desc_7_xid_0_reg
			       ,input [31:0] wr_resp_desc_7_xid_1_reg
			       ,input [31:0] wr_resp_desc_7_xid_2_reg
			       ,input [31:0] wr_resp_desc_7_xid_3_reg
			       ,input [31:0] wr_resp_desc_7_xuser_0_reg
			       ,input [31:0] wr_resp_desc_7_xuser_1_reg
			       ,input [31:0] wr_resp_desc_7_xuser_2_reg
			       ,input [31:0] wr_resp_desc_7_xuser_3_reg
			       ,input [31:0] wr_resp_desc_7_xuser_4_reg
			       ,input [31:0] wr_resp_desc_7_xuser_5_reg
			       ,input [31:0] wr_resp_desc_7_xuser_6_reg
			       ,input [31:0] wr_resp_desc_7_xuser_7_reg
			       ,input [31:0] wr_resp_desc_7_xuser_8_reg
			       ,input [31:0] wr_resp_desc_7_xuser_9_reg
			       ,input [31:0] wr_resp_desc_7_xuser_10_reg
			       ,input [31:0] wr_resp_desc_7_xuser_11_reg
			       ,input [31:0] wr_resp_desc_7_xuser_12_reg
			       ,input [31:0] wr_resp_desc_7_xuser_13_reg
			       ,input [31:0] wr_resp_desc_7_xuser_14_reg
			       ,input [31:0] wr_resp_desc_7_xuser_15_reg
			       ,input [31:0] sn_req_desc_7_attr_reg
			       ,input [31:0] sn_req_desc_7_acaddr_0_reg
			       ,input [31:0] sn_req_desc_7_acaddr_1_reg
			       ,input [31:0] sn_req_desc_7_acaddr_2_reg
			       ,input [31:0] sn_req_desc_7_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_7_resp_reg
			       ,input [31:0] rd_req_desc_8_txn_type_reg
			       ,input [31:0] rd_req_desc_8_size_reg
			       ,input [31:0] rd_req_desc_8_axsize_reg
			       ,input [31:0] rd_req_desc_8_attr_reg
			       ,input [31:0] rd_req_desc_8_axaddr_0_reg
			       ,input [31:0] rd_req_desc_8_axaddr_1_reg
			       ,input [31:0] rd_req_desc_8_axaddr_2_reg
			       ,input [31:0] rd_req_desc_8_axaddr_3_reg
			       ,input [31:0] rd_req_desc_8_axid_0_reg
			       ,input [31:0] rd_req_desc_8_axid_1_reg
			       ,input [31:0] rd_req_desc_8_axid_2_reg
			       ,input [31:0] rd_req_desc_8_axid_3_reg
			       ,input [31:0] rd_req_desc_8_axuser_0_reg
			       ,input [31:0] rd_req_desc_8_axuser_1_reg
			       ,input [31:0] rd_req_desc_8_axuser_2_reg
			       ,input [31:0] rd_req_desc_8_axuser_3_reg
			       ,input [31:0] rd_req_desc_8_axuser_4_reg
			       ,input [31:0] rd_req_desc_8_axuser_5_reg
			       ,input [31:0] rd_req_desc_8_axuser_6_reg
			       ,input [31:0] rd_req_desc_8_axuser_7_reg
			       ,input [31:0] rd_req_desc_8_axuser_8_reg
			       ,input [31:0] rd_req_desc_8_axuser_9_reg
			       ,input [31:0] rd_req_desc_8_axuser_10_reg
			       ,input [31:0] rd_req_desc_8_axuser_11_reg
			       ,input [31:0] rd_req_desc_8_axuser_12_reg
			       ,input [31:0] rd_req_desc_8_axuser_13_reg
			       ,input [31:0] rd_req_desc_8_axuser_14_reg
			       ,input [31:0] rd_req_desc_8_axuser_15_reg
			       ,input [31:0] rd_resp_desc_8_data_offset_reg
			       ,input [31:0] rd_resp_desc_8_data_size_reg
			       ,input [31:0] rd_resp_desc_8_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_8_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_8_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_8_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_8_resp_reg
			       ,input [31:0] rd_resp_desc_8_xid_0_reg
			       ,input [31:0] rd_resp_desc_8_xid_1_reg
			       ,input [31:0] rd_resp_desc_8_xid_2_reg
			       ,input [31:0] rd_resp_desc_8_xid_3_reg
			       ,input [31:0] rd_resp_desc_8_xuser_0_reg
			       ,input [31:0] rd_resp_desc_8_xuser_1_reg
			       ,input [31:0] rd_resp_desc_8_xuser_2_reg
			       ,input [31:0] rd_resp_desc_8_xuser_3_reg
			       ,input [31:0] rd_resp_desc_8_xuser_4_reg
			       ,input [31:0] rd_resp_desc_8_xuser_5_reg
			       ,input [31:0] rd_resp_desc_8_xuser_6_reg
			       ,input [31:0] rd_resp_desc_8_xuser_7_reg
			       ,input [31:0] rd_resp_desc_8_xuser_8_reg
			       ,input [31:0] rd_resp_desc_8_xuser_9_reg
			       ,input [31:0] rd_resp_desc_8_xuser_10_reg
			       ,input [31:0] rd_resp_desc_8_xuser_11_reg
			       ,input [31:0] rd_resp_desc_8_xuser_12_reg
			       ,input [31:0] rd_resp_desc_8_xuser_13_reg
			       ,input [31:0] rd_resp_desc_8_xuser_14_reg
			       ,input [31:0] rd_resp_desc_8_xuser_15_reg
			       ,input [31:0] wr_req_desc_8_txn_type_reg
			       ,input [31:0] wr_req_desc_8_size_reg
			       ,input [31:0] wr_req_desc_8_data_offset_reg
			       ,input [31:0] wr_req_desc_8_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_8_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_8_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_8_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_8_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_8_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_8_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_8_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_8_axsize_reg
			       ,input [31:0] wr_req_desc_8_attr_reg
			       ,input [31:0] wr_req_desc_8_axaddr_0_reg
			       ,input [31:0] wr_req_desc_8_axaddr_1_reg
			       ,input [31:0] wr_req_desc_8_axaddr_2_reg
			       ,input [31:0] wr_req_desc_8_axaddr_3_reg
			       ,input [31:0] wr_req_desc_8_axid_0_reg
			       ,input [31:0] wr_req_desc_8_axid_1_reg
			       ,input [31:0] wr_req_desc_8_axid_2_reg
			       ,input [31:0] wr_req_desc_8_axid_3_reg
			       ,input [31:0] wr_req_desc_8_axuser_0_reg
			       ,input [31:0] wr_req_desc_8_axuser_1_reg
			       ,input [31:0] wr_req_desc_8_axuser_2_reg
			       ,input [31:0] wr_req_desc_8_axuser_3_reg
			       ,input [31:0] wr_req_desc_8_axuser_4_reg
			       ,input [31:0] wr_req_desc_8_axuser_5_reg
			       ,input [31:0] wr_req_desc_8_axuser_6_reg
			       ,input [31:0] wr_req_desc_8_axuser_7_reg
			       ,input [31:0] wr_req_desc_8_axuser_8_reg
			       ,input [31:0] wr_req_desc_8_axuser_9_reg
			       ,input [31:0] wr_req_desc_8_axuser_10_reg
			       ,input [31:0] wr_req_desc_8_axuser_11_reg
			       ,input [31:0] wr_req_desc_8_axuser_12_reg
			       ,input [31:0] wr_req_desc_8_axuser_13_reg
			       ,input [31:0] wr_req_desc_8_axuser_14_reg
			       ,input [31:0] wr_req_desc_8_axuser_15_reg
			       ,input [31:0] wr_req_desc_8_wuser_0_reg
			       ,input [31:0] wr_req_desc_8_wuser_1_reg
			       ,input [31:0] wr_req_desc_8_wuser_2_reg
			       ,input [31:0] wr_req_desc_8_wuser_3_reg
			       ,input [31:0] wr_req_desc_8_wuser_4_reg
			       ,input [31:0] wr_req_desc_8_wuser_5_reg
			       ,input [31:0] wr_req_desc_8_wuser_6_reg
			       ,input [31:0] wr_req_desc_8_wuser_7_reg
			       ,input [31:0] wr_req_desc_8_wuser_8_reg
			       ,input [31:0] wr_req_desc_8_wuser_9_reg
			       ,input [31:0] wr_req_desc_8_wuser_10_reg
			       ,input [31:0] wr_req_desc_8_wuser_11_reg
			       ,input [31:0] wr_req_desc_8_wuser_12_reg
			       ,input [31:0] wr_req_desc_8_wuser_13_reg
			       ,input [31:0] wr_req_desc_8_wuser_14_reg
			       ,input [31:0] wr_req_desc_8_wuser_15_reg
			       ,input [31:0] wr_resp_desc_8_resp_reg
			       ,input [31:0] wr_resp_desc_8_xid_0_reg
			       ,input [31:0] wr_resp_desc_8_xid_1_reg
			       ,input [31:0] wr_resp_desc_8_xid_2_reg
			       ,input [31:0] wr_resp_desc_8_xid_3_reg
			       ,input [31:0] wr_resp_desc_8_xuser_0_reg
			       ,input [31:0] wr_resp_desc_8_xuser_1_reg
			       ,input [31:0] wr_resp_desc_8_xuser_2_reg
			       ,input [31:0] wr_resp_desc_8_xuser_3_reg
			       ,input [31:0] wr_resp_desc_8_xuser_4_reg
			       ,input [31:0] wr_resp_desc_8_xuser_5_reg
			       ,input [31:0] wr_resp_desc_8_xuser_6_reg
			       ,input [31:0] wr_resp_desc_8_xuser_7_reg
			       ,input [31:0] wr_resp_desc_8_xuser_8_reg
			       ,input [31:0] wr_resp_desc_8_xuser_9_reg
			       ,input [31:0] wr_resp_desc_8_xuser_10_reg
			       ,input [31:0] wr_resp_desc_8_xuser_11_reg
			       ,input [31:0] wr_resp_desc_8_xuser_12_reg
			       ,input [31:0] wr_resp_desc_8_xuser_13_reg
			       ,input [31:0] wr_resp_desc_8_xuser_14_reg
			       ,input [31:0] wr_resp_desc_8_xuser_15_reg
			       ,input [31:0] sn_req_desc_8_attr_reg
			       ,input [31:0] sn_req_desc_8_acaddr_0_reg
			       ,input [31:0] sn_req_desc_8_acaddr_1_reg
			       ,input [31:0] sn_req_desc_8_acaddr_2_reg
			       ,input [31:0] sn_req_desc_8_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_8_resp_reg
			       ,input [31:0] rd_req_desc_9_txn_type_reg
			       ,input [31:0] rd_req_desc_9_size_reg
			       ,input [31:0] rd_req_desc_9_axsize_reg
			       ,input [31:0] rd_req_desc_9_attr_reg
			       ,input [31:0] rd_req_desc_9_axaddr_0_reg
			       ,input [31:0] rd_req_desc_9_axaddr_1_reg
			       ,input [31:0] rd_req_desc_9_axaddr_2_reg
			       ,input [31:0] rd_req_desc_9_axaddr_3_reg
			       ,input [31:0] rd_req_desc_9_axid_0_reg
			       ,input [31:0] rd_req_desc_9_axid_1_reg
			       ,input [31:0] rd_req_desc_9_axid_2_reg
			       ,input [31:0] rd_req_desc_9_axid_3_reg
			       ,input [31:0] rd_req_desc_9_axuser_0_reg
			       ,input [31:0] rd_req_desc_9_axuser_1_reg
			       ,input [31:0] rd_req_desc_9_axuser_2_reg
			       ,input [31:0] rd_req_desc_9_axuser_3_reg
			       ,input [31:0] rd_req_desc_9_axuser_4_reg
			       ,input [31:0] rd_req_desc_9_axuser_5_reg
			       ,input [31:0] rd_req_desc_9_axuser_6_reg
			       ,input [31:0] rd_req_desc_9_axuser_7_reg
			       ,input [31:0] rd_req_desc_9_axuser_8_reg
			       ,input [31:0] rd_req_desc_9_axuser_9_reg
			       ,input [31:0] rd_req_desc_9_axuser_10_reg
			       ,input [31:0] rd_req_desc_9_axuser_11_reg
			       ,input [31:0] rd_req_desc_9_axuser_12_reg
			       ,input [31:0] rd_req_desc_9_axuser_13_reg
			       ,input [31:0] rd_req_desc_9_axuser_14_reg
			       ,input [31:0] rd_req_desc_9_axuser_15_reg
			       ,input [31:0] rd_resp_desc_9_data_offset_reg
			       ,input [31:0] rd_resp_desc_9_data_size_reg
			       ,input [31:0] rd_resp_desc_9_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_9_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_9_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_9_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_9_resp_reg
			       ,input [31:0] rd_resp_desc_9_xid_0_reg
			       ,input [31:0] rd_resp_desc_9_xid_1_reg
			       ,input [31:0] rd_resp_desc_9_xid_2_reg
			       ,input [31:0] rd_resp_desc_9_xid_3_reg
			       ,input [31:0] rd_resp_desc_9_xuser_0_reg
			       ,input [31:0] rd_resp_desc_9_xuser_1_reg
			       ,input [31:0] rd_resp_desc_9_xuser_2_reg
			       ,input [31:0] rd_resp_desc_9_xuser_3_reg
			       ,input [31:0] rd_resp_desc_9_xuser_4_reg
			       ,input [31:0] rd_resp_desc_9_xuser_5_reg
			       ,input [31:0] rd_resp_desc_9_xuser_6_reg
			       ,input [31:0] rd_resp_desc_9_xuser_7_reg
			       ,input [31:0] rd_resp_desc_9_xuser_8_reg
			       ,input [31:0] rd_resp_desc_9_xuser_9_reg
			       ,input [31:0] rd_resp_desc_9_xuser_10_reg
			       ,input [31:0] rd_resp_desc_9_xuser_11_reg
			       ,input [31:0] rd_resp_desc_9_xuser_12_reg
			       ,input [31:0] rd_resp_desc_9_xuser_13_reg
			       ,input [31:0] rd_resp_desc_9_xuser_14_reg
			       ,input [31:0] rd_resp_desc_9_xuser_15_reg
			       ,input [31:0] wr_req_desc_9_txn_type_reg
			       ,input [31:0] wr_req_desc_9_size_reg
			       ,input [31:0] wr_req_desc_9_data_offset_reg
			       ,input [31:0] wr_req_desc_9_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_9_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_9_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_9_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_9_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_9_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_9_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_9_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_9_axsize_reg
			       ,input [31:0] wr_req_desc_9_attr_reg
			       ,input [31:0] wr_req_desc_9_axaddr_0_reg
			       ,input [31:0] wr_req_desc_9_axaddr_1_reg
			       ,input [31:0] wr_req_desc_9_axaddr_2_reg
			       ,input [31:0] wr_req_desc_9_axaddr_3_reg
			       ,input [31:0] wr_req_desc_9_axid_0_reg
			       ,input [31:0] wr_req_desc_9_axid_1_reg
			       ,input [31:0] wr_req_desc_9_axid_2_reg
			       ,input [31:0] wr_req_desc_9_axid_3_reg
			       ,input [31:0] wr_req_desc_9_axuser_0_reg
			       ,input [31:0] wr_req_desc_9_axuser_1_reg
			       ,input [31:0] wr_req_desc_9_axuser_2_reg
			       ,input [31:0] wr_req_desc_9_axuser_3_reg
			       ,input [31:0] wr_req_desc_9_axuser_4_reg
			       ,input [31:0] wr_req_desc_9_axuser_5_reg
			       ,input [31:0] wr_req_desc_9_axuser_6_reg
			       ,input [31:0] wr_req_desc_9_axuser_7_reg
			       ,input [31:0] wr_req_desc_9_axuser_8_reg
			       ,input [31:0] wr_req_desc_9_axuser_9_reg
			       ,input [31:0] wr_req_desc_9_axuser_10_reg
			       ,input [31:0] wr_req_desc_9_axuser_11_reg
			       ,input [31:0] wr_req_desc_9_axuser_12_reg
			       ,input [31:0] wr_req_desc_9_axuser_13_reg
			       ,input [31:0] wr_req_desc_9_axuser_14_reg
			       ,input [31:0] wr_req_desc_9_axuser_15_reg
			       ,input [31:0] wr_req_desc_9_wuser_0_reg
			       ,input [31:0] wr_req_desc_9_wuser_1_reg
			       ,input [31:0] wr_req_desc_9_wuser_2_reg
			       ,input [31:0] wr_req_desc_9_wuser_3_reg
			       ,input [31:0] wr_req_desc_9_wuser_4_reg
			       ,input [31:0] wr_req_desc_9_wuser_5_reg
			       ,input [31:0] wr_req_desc_9_wuser_6_reg
			       ,input [31:0] wr_req_desc_9_wuser_7_reg
			       ,input [31:0] wr_req_desc_9_wuser_8_reg
			       ,input [31:0] wr_req_desc_9_wuser_9_reg
			       ,input [31:0] wr_req_desc_9_wuser_10_reg
			       ,input [31:0] wr_req_desc_9_wuser_11_reg
			       ,input [31:0] wr_req_desc_9_wuser_12_reg
			       ,input [31:0] wr_req_desc_9_wuser_13_reg
			       ,input [31:0] wr_req_desc_9_wuser_14_reg
			       ,input [31:0] wr_req_desc_9_wuser_15_reg
			       ,input [31:0] wr_resp_desc_9_resp_reg
			       ,input [31:0] wr_resp_desc_9_xid_0_reg
			       ,input [31:0] wr_resp_desc_9_xid_1_reg
			       ,input [31:0] wr_resp_desc_9_xid_2_reg
			       ,input [31:0] wr_resp_desc_9_xid_3_reg
			       ,input [31:0] wr_resp_desc_9_xuser_0_reg
			       ,input [31:0] wr_resp_desc_9_xuser_1_reg
			       ,input [31:0] wr_resp_desc_9_xuser_2_reg
			       ,input [31:0] wr_resp_desc_9_xuser_3_reg
			       ,input [31:0] wr_resp_desc_9_xuser_4_reg
			       ,input [31:0] wr_resp_desc_9_xuser_5_reg
			       ,input [31:0] wr_resp_desc_9_xuser_6_reg
			       ,input [31:0] wr_resp_desc_9_xuser_7_reg
			       ,input [31:0] wr_resp_desc_9_xuser_8_reg
			       ,input [31:0] wr_resp_desc_9_xuser_9_reg
			       ,input [31:0] wr_resp_desc_9_xuser_10_reg
			       ,input [31:0] wr_resp_desc_9_xuser_11_reg
			       ,input [31:0] wr_resp_desc_9_xuser_12_reg
			       ,input [31:0] wr_resp_desc_9_xuser_13_reg
			       ,input [31:0] wr_resp_desc_9_xuser_14_reg
			       ,input [31:0] wr_resp_desc_9_xuser_15_reg
			       ,input [31:0] sn_req_desc_9_attr_reg
			       ,input [31:0] sn_req_desc_9_acaddr_0_reg
			       ,input [31:0] sn_req_desc_9_acaddr_1_reg
			       ,input [31:0] sn_req_desc_9_acaddr_2_reg
			       ,input [31:0] sn_req_desc_9_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_9_resp_reg
			       ,input [31:0] rd_req_desc_a_txn_type_reg
			       ,input [31:0] rd_req_desc_a_size_reg
			       ,input [31:0] rd_req_desc_a_axsize_reg
			       ,input [31:0] rd_req_desc_a_attr_reg
			       ,input [31:0] rd_req_desc_a_axaddr_0_reg
			       ,input [31:0] rd_req_desc_a_axaddr_1_reg
			       ,input [31:0] rd_req_desc_a_axaddr_2_reg
			       ,input [31:0] rd_req_desc_a_axaddr_3_reg
			       ,input [31:0] rd_req_desc_a_axid_0_reg
			       ,input [31:0] rd_req_desc_a_axid_1_reg
			       ,input [31:0] rd_req_desc_a_axid_2_reg
			       ,input [31:0] rd_req_desc_a_axid_3_reg
			       ,input [31:0] rd_req_desc_a_axuser_0_reg
			       ,input [31:0] rd_req_desc_a_axuser_1_reg
			       ,input [31:0] rd_req_desc_a_axuser_2_reg
			       ,input [31:0] rd_req_desc_a_axuser_3_reg
			       ,input [31:0] rd_req_desc_a_axuser_4_reg
			       ,input [31:0] rd_req_desc_a_axuser_5_reg
			       ,input [31:0] rd_req_desc_a_axuser_6_reg
			       ,input [31:0] rd_req_desc_a_axuser_7_reg
			       ,input [31:0] rd_req_desc_a_axuser_8_reg
			       ,input [31:0] rd_req_desc_a_axuser_9_reg
			       ,input [31:0] rd_req_desc_a_axuser_10_reg
			       ,input [31:0] rd_req_desc_a_axuser_11_reg
			       ,input [31:0] rd_req_desc_a_axuser_12_reg
			       ,input [31:0] rd_req_desc_a_axuser_13_reg
			       ,input [31:0] rd_req_desc_a_axuser_14_reg
			       ,input [31:0] rd_req_desc_a_axuser_15_reg
			       ,input [31:0] rd_resp_desc_a_data_offset_reg
			       ,input [31:0] rd_resp_desc_a_data_size_reg
			       ,input [31:0] rd_resp_desc_a_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_a_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_a_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_a_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_a_resp_reg
			       ,input [31:0] rd_resp_desc_a_xid_0_reg
			       ,input [31:0] rd_resp_desc_a_xid_1_reg
			       ,input [31:0] rd_resp_desc_a_xid_2_reg
			       ,input [31:0] rd_resp_desc_a_xid_3_reg
			       ,input [31:0] rd_resp_desc_a_xuser_0_reg
			       ,input [31:0] rd_resp_desc_a_xuser_1_reg
			       ,input [31:0] rd_resp_desc_a_xuser_2_reg
			       ,input [31:0] rd_resp_desc_a_xuser_3_reg
			       ,input [31:0] rd_resp_desc_a_xuser_4_reg
			       ,input [31:0] rd_resp_desc_a_xuser_5_reg
			       ,input [31:0] rd_resp_desc_a_xuser_6_reg
			       ,input [31:0] rd_resp_desc_a_xuser_7_reg
			       ,input [31:0] rd_resp_desc_a_xuser_8_reg
			       ,input [31:0] rd_resp_desc_a_xuser_9_reg
			       ,input [31:0] rd_resp_desc_a_xuser_10_reg
			       ,input [31:0] rd_resp_desc_a_xuser_11_reg
			       ,input [31:0] rd_resp_desc_a_xuser_12_reg
			       ,input [31:0] rd_resp_desc_a_xuser_13_reg
			       ,input [31:0] rd_resp_desc_a_xuser_14_reg
			       ,input [31:0] rd_resp_desc_a_xuser_15_reg
			       ,input [31:0] wr_req_desc_a_txn_type_reg
			       ,input [31:0] wr_req_desc_a_size_reg
			       ,input [31:0] wr_req_desc_a_data_offset_reg
			       ,input [31:0] wr_req_desc_a_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_a_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_a_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_a_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_a_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_a_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_a_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_a_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_a_axsize_reg
			       ,input [31:0] wr_req_desc_a_attr_reg
			       ,input [31:0] wr_req_desc_a_axaddr_0_reg
			       ,input [31:0] wr_req_desc_a_axaddr_1_reg
			       ,input [31:0] wr_req_desc_a_axaddr_2_reg
			       ,input [31:0] wr_req_desc_a_axaddr_3_reg
			       ,input [31:0] wr_req_desc_a_axid_0_reg
			       ,input [31:0] wr_req_desc_a_axid_1_reg
			       ,input [31:0] wr_req_desc_a_axid_2_reg
			       ,input [31:0] wr_req_desc_a_axid_3_reg
			       ,input [31:0] wr_req_desc_a_axuser_0_reg
			       ,input [31:0] wr_req_desc_a_axuser_1_reg
			       ,input [31:0] wr_req_desc_a_axuser_2_reg
			       ,input [31:0] wr_req_desc_a_axuser_3_reg
			       ,input [31:0] wr_req_desc_a_axuser_4_reg
			       ,input [31:0] wr_req_desc_a_axuser_5_reg
			       ,input [31:0] wr_req_desc_a_axuser_6_reg
			       ,input [31:0] wr_req_desc_a_axuser_7_reg
			       ,input [31:0] wr_req_desc_a_axuser_8_reg
			       ,input [31:0] wr_req_desc_a_axuser_9_reg
			       ,input [31:0] wr_req_desc_a_axuser_10_reg
			       ,input [31:0] wr_req_desc_a_axuser_11_reg
			       ,input [31:0] wr_req_desc_a_axuser_12_reg
			       ,input [31:0] wr_req_desc_a_axuser_13_reg
			       ,input [31:0] wr_req_desc_a_axuser_14_reg
			       ,input [31:0] wr_req_desc_a_axuser_15_reg
			       ,input [31:0] wr_req_desc_a_wuser_0_reg
			       ,input [31:0] wr_req_desc_a_wuser_1_reg
			       ,input [31:0] wr_req_desc_a_wuser_2_reg
			       ,input [31:0] wr_req_desc_a_wuser_3_reg
			       ,input [31:0] wr_req_desc_a_wuser_4_reg
			       ,input [31:0] wr_req_desc_a_wuser_5_reg
			       ,input [31:0] wr_req_desc_a_wuser_6_reg
			       ,input [31:0] wr_req_desc_a_wuser_7_reg
			       ,input [31:0] wr_req_desc_a_wuser_8_reg
			       ,input [31:0] wr_req_desc_a_wuser_9_reg
			       ,input [31:0] wr_req_desc_a_wuser_10_reg
			       ,input [31:0] wr_req_desc_a_wuser_11_reg
			       ,input [31:0] wr_req_desc_a_wuser_12_reg
			       ,input [31:0] wr_req_desc_a_wuser_13_reg
			       ,input [31:0] wr_req_desc_a_wuser_14_reg
			       ,input [31:0] wr_req_desc_a_wuser_15_reg
			       ,input [31:0] wr_resp_desc_a_resp_reg
			       ,input [31:0] wr_resp_desc_a_xid_0_reg
			       ,input [31:0] wr_resp_desc_a_xid_1_reg
			       ,input [31:0] wr_resp_desc_a_xid_2_reg
			       ,input [31:0] wr_resp_desc_a_xid_3_reg
			       ,input [31:0] wr_resp_desc_a_xuser_0_reg
			       ,input [31:0] wr_resp_desc_a_xuser_1_reg
			       ,input [31:0] wr_resp_desc_a_xuser_2_reg
			       ,input [31:0] wr_resp_desc_a_xuser_3_reg
			       ,input [31:0] wr_resp_desc_a_xuser_4_reg
			       ,input [31:0] wr_resp_desc_a_xuser_5_reg
			       ,input [31:0] wr_resp_desc_a_xuser_6_reg
			       ,input [31:0] wr_resp_desc_a_xuser_7_reg
			       ,input [31:0] wr_resp_desc_a_xuser_8_reg
			       ,input [31:0] wr_resp_desc_a_xuser_9_reg
			       ,input [31:0] wr_resp_desc_a_xuser_10_reg
			       ,input [31:0] wr_resp_desc_a_xuser_11_reg
			       ,input [31:0] wr_resp_desc_a_xuser_12_reg
			       ,input [31:0] wr_resp_desc_a_xuser_13_reg
			       ,input [31:0] wr_resp_desc_a_xuser_14_reg
			       ,input [31:0] wr_resp_desc_a_xuser_15_reg
			       ,input [31:0] sn_req_desc_a_attr_reg
			       ,input [31:0] sn_req_desc_a_acaddr_0_reg
			       ,input [31:0] sn_req_desc_a_acaddr_1_reg
			       ,input [31:0] sn_req_desc_a_acaddr_2_reg
			       ,input [31:0] sn_req_desc_a_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_a_resp_reg
			       ,input [31:0] rd_req_desc_b_txn_type_reg
			       ,input [31:0] rd_req_desc_b_size_reg
			       ,input [31:0] rd_req_desc_b_axsize_reg
			       ,input [31:0] rd_req_desc_b_attr_reg
			       ,input [31:0] rd_req_desc_b_axaddr_0_reg
			       ,input [31:0] rd_req_desc_b_axaddr_1_reg
			       ,input [31:0] rd_req_desc_b_axaddr_2_reg
			       ,input [31:0] rd_req_desc_b_axaddr_3_reg
			       ,input [31:0] rd_req_desc_b_axid_0_reg
			       ,input [31:0] rd_req_desc_b_axid_1_reg
			       ,input [31:0] rd_req_desc_b_axid_2_reg
			       ,input [31:0] rd_req_desc_b_axid_3_reg
			       ,input [31:0] rd_req_desc_b_axuser_0_reg
			       ,input [31:0] rd_req_desc_b_axuser_1_reg
			       ,input [31:0] rd_req_desc_b_axuser_2_reg
			       ,input [31:0] rd_req_desc_b_axuser_3_reg
			       ,input [31:0] rd_req_desc_b_axuser_4_reg
			       ,input [31:0] rd_req_desc_b_axuser_5_reg
			       ,input [31:0] rd_req_desc_b_axuser_6_reg
			       ,input [31:0] rd_req_desc_b_axuser_7_reg
			       ,input [31:0] rd_req_desc_b_axuser_8_reg
			       ,input [31:0] rd_req_desc_b_axuser_9_reg
			       ,input [31:0] rd_req_desc_b_axuser_10_reg
			       ,input [31:0] rd_req_desc_b_axuser_11_reg
			       ,input [31:0] rd_req_desc_b_axuser_12_reg
			       ,input [31:0] rd_req_desc_b_axuser_13_reg
			       ,input [31:0] rd_req_desc_b_axuser_14_reg
			       ,input [31:0] rd_req_desc_b_axuser_15_reg
			       ,input [31:0] rd_resp_desc_b_data_offset_reg
			       ,input [31:0] rd_resp_desc_b_data_size_reg
			       ,input [31:0] rd_resp_desc_b_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_b_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_b_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_b_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_b_resp_reg
			       ,input [31:0] rd_resp_desc_b_xid_0_reg
			       ,input [31:0] rd_resp_desc_b_xid_1_reg
			       ,input [31:0] rd_resp_desc_b_xid_2_reg
			       ,input [31:0] rd_resp_desc_b_xid_3_reg
			       ,input [31:0] rd_resp_desc_b_xuser_0_reg
			       ,input [31:0] rd_resp_desc_b_xuser_1_reg
			       ,input [31:0] rd_resp_desc_b_xuser_2_reg
			       ,input [31:0] rd_resp_desc_b_xuser_3_reg
			       ,input [31:0] rd_resp_desc_b_xuser_4_reg
			       ,input [31:0] rd_resp_desc_b_xuser_5_reg
			       ,input [31:0] rd_resp_desc_b_xuser_6_reg
			       ,input [31:0] rd_resp_desc_b_xuser_7_reg
			       ,input [31:0] rd_resp_desc_b_xuser_8_reg
			       ,input [31:0] rd_resp_desc_b_xuser_9_reg
			       ,input [31:0] rd_resp_desc_b_xuser_10_reg
			       ,input [31:0] rd_resp_desc_b_xuser_11_reg
			       ,input [31:0] rd_resp_desc_b_xuser_12_reg
			       ,input [31:0] rd_resp_desc_b_xuser_13_reg
			       ,input [31:0] rd_resp_desc_b_xuser_14_reg
			       ,input [31:0] rd_resp_desc_b_xuser_15_reg
			       ,input [31:0] wr_req_desc_b_txn_type_reg
			       ,input [31:0] wr_req_desc_b_size_reg
			       ,input [31:0] wr_req_desc_b_data_offset_reg
			       ,input [31:0] wr_req_desc_b_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_b_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_b_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_b_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_b_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_b_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_b_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_b_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_b_axsize_reg
			       ,input [31:0] wr_req_desc_b_attr_reg
			       ,input [31:0] wr_req_desc_b_axaddr_0_reg
			       ,input [31:0] wr_req_desc_b_axaddr_1_reg
			       ,input [31:0] wr_req_desc_b_axaddr_2_reg
			       ,input [31:0] wr_req_desc_b_axaddr_3_reg
			       ,input [31:0] wr_req_desc_b_axid_0_reg
			       ,input [31:0] wr_req_desc_b_axid_1_reg
			       ,input [31:0] wr_req_desc_b_axid_2_reg
			       ,input [31:0] wr_req_desc_b_axid_3_reg
			       ,input [31:0] wr_req_desc_b_axuser_0_reg
			       ,input [31:0] wr_req_desc_b_axuser_1_reg
			       ,input [31:0] wr_req_desc_b_axuser_2_reg
			       ,input [31:0] wr_req_desc_b_axuser_3_reg
			       ,input [31:0] wr_req_desc_b_axuser_4_reg
			       ,input [31:0] wr_req_desc_b_axuser_5_reg
			       ,input [31:0] wr_req_desc_b_axuser_6_reg
			       ,input [31:0] wr_req_desc_b_axuser_7_reg
			       ,input [31:0] wr_req_desc_b_axuser_8_reg
			       ,input [31:0] wr_req_desc_b_axuser_9_reg
			       ,input [31:0] wr_req_desc_b_axuser_10_reg
			       ,input [31:0] wr_req_desc_b_axuser_11_reg
			       ,input [31:0] wr_req_desc_b_axuser_12_reg
			       ,input [31:0] wr_req_desc_b_axuser_13_reg
			       ,input [31:0] wr_req_desc_b_axuser_14_reg
			       ,input [31:0] wr_req_desc_b_axuser_15_reg
			       ,input [31:0] wr_req_desc_b_wuser_0_reg
			       ,input [31:0] wr_req_desc_b_wuser_1_reg
			       ,input [31:0] wr_req_desc_b_wuser_2_reg
			       ,input [31:0] wr_req_desc_b_wuser_3_reg
			       ,input [31:0] wr_req_desc_b_wuser_4_reg
			       ,input [31:0] wr_req_desc_b_wuser_5_reg
			       ,input [31:0] wr_req_desc_b_wuser_6_reg
			       ,input [31:0] wr_req_desc_b_wuser_7_reg
			       ,input [31:0] wr_req_desc_b_wuser_8_reg
			       ,input [31:0] wr_req_desc_b_wuser_9_reg
			       ,input [31:0] wr_req_desc_b_wuser_10_reg
			       ,input [31:0] wr_req_desc_b_wuser_11_reg
			       ,input [31:0] wr_req_desc_b_wuser_12_reg
			       ,input [31:0] wr_req_desc_b_wuser_13_reg
			       ,input [31:0] wr_req_desc_b_wuser_14_reg
			       ,input [31:0] wr_req_desc_b_wuser_15_reg
			       ,input [31:0] wr_resp_desc_b_resp_reg
			       ,input [31:0] wr_resp_desc_b_xid_0_reg
			       ,input [31:0] wr_resp_desc_b_xid_1_reg
			       ,input [31:0] wr_resp_desc_b_xid_2_reg
			       ,input [31:0] wr_resp_desc_b_xid_3_reg
			       ,input [31:0] wr_resp_desc_b_xuser_0_reg
			       ,input [31:0] wr_resp_desc_b_xuser_1_reg
			       ,input [31:0] wr_resp_desc_b_xuser_2_reg
			       ,input [31:0] wr_resp_desc_b_xuser_3_reg
			       ,input [31:0] wr_resp_desc_b_xuser_4_reg
			       ,input [31:0] wr_resp_desc_b_xuser_5_reg
			       ,input [31:0] wr_resp_desc_b_xuser_6_reg
			       ,input [31:0] wr_resp_desc_b_xuser_7_reg
			       ,input [31:0] wr_resp_desc_b_xuser_8_reg
			       ,input [31:0] wr_resp_desc_b_xuser_9_reg
			       ,input [31:0] wr_resp_desc_b_xuser_10_reg
			       ,input [31:0] wr_resp_desc_b_xuser_11_reg
			       ,input [31:0] wr_resp_desc_b_xuser_12_reg
			       ,input [31:0] wr_resp_desc_b_xuser_13_reg
			       ,input [31:0] wr_resp_desc_b_xuser_14_reg
			       ,input [31:0] wr_resp_desc_b_xuser_15_reg
			       ,input [31:0] sn_req_desc_b_attr_reg
			       ,input [31:0] sn_req_desc_b_acaddr_0_reg
			       ,input [31:0] sn_req_desc_b_acaddr_1_reg
			       ,input [31:0] sn_req_desc_b_acaddr_2_reg
			       ,input [31:0] sn_req_desc_b_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_b_resp_reg
			       ,input [31:0] rd_req_desc_c_txn_type_reg
			       ,input [31:0] rd_req_desc_c_size_reg
			       ,input [31:0] rd_req_desc_c_axsize_reg
			       ,input [31:0] rd_req_desc_c_attr_reg
			       ,input [31:0] rd_req_desc_c_axaddr_0_reg
			       ,input [31:0] rd_req_desc_c_axaddr_1_reg
			       ,input [31:0] rd_req_desc_c_axaddr_2_reg
			       ,input [31:0] rd_req_desc_c_axaddr_3_reg
			       ,input [31:0] rd_req_desc_c_axid_0_reg
			       ,input [31:0] rd_req_desc_c_axid_1_reg
			       ,input [31:0] rd_req_desc_c_axid_2_reg
			       ,input [31:0] rd_req_desc_c_axid_3_reg
			       ,input [31:0] rd_req_desc_c_axuser_0_reg
			       ,input [31:0] rd_req_desc_c_axuser_1_reg
			       ,input [31:0] rd_req_desc_c_axuser_2_reg
			       ,input [31:0] rd_req_desc_c_axuser_3_reg
			       ,input [31:0] rd_req_desc_c_axuser_4_reg
			       ,input [31:0] rd_req_desc_c_axuser_5_reg
			       ,input [31:0] rd_req_desc_c_axuser_6_reg
			       ,input [31:0] rd_req_desc_c_axuser_7_reg
			       ,input [31:0] rd_req_desc_c_axuser_8_reg
			       ,input [31:0] rd_req_desc_c_axuser_9_reg
			       ,input [31:0] rd_req_desc_c_axuser_10_reg
			       ,input [31:0] rd_req_desc_c_axuser_11_reg
			       ,input [31:0] rd_req_desc_c_axuser_12_reg
			       ,input [31:0] rd_req_desc_c_axuser_13_reg
			       ,input [31:0] rd_req_desc_c_axuser_14_reg
			       ,input [31:0] rd_req_desc_c_axuser_15_reg
			       ,input [31:0] rd_resp_desc_c_data_offset_reg
			       ,input [31:0] rd_resp_desc_c_data_size_reg
			       ,input [31:0] rd_resp_desc_c_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_c_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_c_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_c_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_c_resp_reg
			       ,input [31:0] rd_resp_desc_c_xid_0_reg
			       ,input [31:0] rd_resp_desc_c_xid_1_reg
			       ,input [31:0] rd_resp_desc_c_xid_2_reg
			       ,input [31:0] rd_resp_desc_c_xid_3_reg
			       ,input [31:0] rd_resp_desc_c_xuser_0_reg
			       ,input [31:0] rd_resp_desc_c_xuser_1_reg
			       ,input [31:0] rd_resp_desc_c_xuser_2_reg
			       ,input [31:0] rd_resp_desc_c_xuser_3_reg
			       ,input [31:0] rd_resp_desc_c_xuser_4_reg
			       ,input [31:0] rd_resp_desc_c_xuser_5_reg
			       ,input [31:0] rd_resp_desc_c_xuser_6_reg
			       ,input [31:0] rd_resp_desc_c_xuser_7_reg
			       ,input [31:0] rd_resp_desc_c_xuser_8_reg
			       ,input [31:0] rd_resp_desc_c_xuser_9_reg
			       ,input [31:0] rd_resp_desc_c_xuser_10_reg
			       ,input [31:0] rd_resp_desc_c_xuser_11_reg
			       ,input [31:0] rd_resp_desc_c_xuser_12_reg
			       ,input [31:0] rd_resp_desc_c_xuser_13_reg
			       ,input [31:0] rd_resp_desc_c_xuser_14_reg
			       ,input [31:0] rd_resp_desc_c_xuser_15_reg
			       ,input [31:0] wr_req_desc_c_txn_type_reg
			       ,input [31:0] wr_req_desc_c_size_reg
			       ,input [31:0] wr_req_desc_c_data_offset_reg
			       ,input [31:0] wr_req_desc_c_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_c_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_c_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_c_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_c_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_c_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_c_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_c_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_c_axsize_reg
			       ,input [31:0] wr_req_desc_c_attr_reg
			       ,input [31:0] wr_req_desc_c_axaddr_0_reg
			       ,input [31:0] wr_req_desc_c_axaddr_1_reg
			       ,input [31:0] wr_req_desc_c_axaddr_2_reg
			       ,input [31:0] wr_req_desc_c_axaddr_3_reg
			       ,input [31:0] wr_req_desc_c_axid_0_reg
			       ,input [31:0] wr_req_desc_c_axid_1_reg
			       ,input [31:0] wr_req_desc_c_axid_2_reg
			       ,input [31:0] wr_req_desc_c_axid_3_reg
			       ,input [31:0] wr_req_desc_c_axuser_0_reg
			       ,input [31:0] wr_req_desc_c_axuser_1_reg
			       ,input [31:0] wr_req_desc_c_axuser_2_reg
			       ,input [31:0] wr_req_desc_c_axuser_3_reg
			       ,input [31:0] wr_req_desc_c_axuser_4_reg
			       ,input [31:0] wr_req_desc_c_axuser_5_reg
			       ,input [31:0] wr_req_desc_c_axuser_6_reg
			       ,input [31:0] wr_req_desc_c_axuser_7_reg
			       ,input [31:0] wr_req_desc_c_axuser_8_reg
			       ,input [31:0] wr_req_desc_c_axuser_9_reg
			       ,input [31:0] wr_req_desc_c_axuser_10_reg
			       ,input [31:0] wr_req_desc_c_axuser_11_reg
			       ,input [31:0] wr_req_desc_c_axuser_12_reg
			       ,input [31:0] wr_req_desc_c_axuser_13_reg
			       ,input [31:0] wr_req_desc_c_axuser_14_reg
			       ,input [31:0] wr_req_desc_c_axuser_15_reg
			       ,input [31:0] wr_req_desc_c_wuser_0_reg
			       ,input [31:0] wr_req_desc_c_wuser_1_reg
			       ,input [31:0] wr_req_desc_c_wuser_2_reg
			       ,input [31:0] wr_req_desc_c_wuser_3_reg
			       ,input [31:0] wr_req_desc_c_wuser_4_reg
			       ,input [31:0] wr_req_desc_c_wuser_5_reg
			       ,input [31:0] wr_req_desc_c_wuser_6_reg
			       ,input [31:0] wr_req_desc_c_wuser_7_reg
			       ,input [31:0] wr_req_desc_c_wuser_8_reg
			       ,input [31:0] wr_req_desc_c_wuser_9_reg
			       ,input [31:0] wr_req_desc_c_wuser_10_reg
			       ,input [31:0] wr_req_desc_c_wuser_11_reg
			       ,input [31:0] wr_req_desc_c_wuser_12_reg
			       ,input [31:0] wr_req_desc_c_wuser_13_reg
			       ,input [31:0] wr_req_desc_c_wuser_14_reg
			       ,input [31:0] wr_req_desc_c_wuser_15_reg
			       ,input [31:0] wr_resp_desc_c_resp_reg
			       ,input [31:0] wr_resp_desc_c_xid_0_reg
			       ,input [31:0] wr_resp_desc_c_xid_1_reg
			       ,input [31:0] wr_resp_desc_c_xid_2_reg
			       ,input [31:0] wr_resp_desc_c_xid_3_reg
			       ,input [31:0] wr_resp_desc_c_xuser_0_reg
			       ,input [31:0] wr_resp_desc_c_xuser_1_reg
			       ,input [31:0] wr_resp_desc_c_xuser_2_reg
			       ,input [31:0] wr_resp_desc_c_xuser_3_reg
			       ,input [31:0] wr_resp_desc_c_xuser_4_reg
			       ,input [31:0] wr_resp_desc_c_xuser_5_reg
			       ,input [31:0] wr_resp_desc_c_xuser_6_reg
			       ,input [31:0] wr_resp_desc_c_xuser_7_reg
			       ,input [31:0] wr_resp_desc_c_xuser_8_reg
			       ,input [31:0] wr_resp_desc_c_xuser_9_reg
			       ,input [31:0] wr_resp_desc_c_xuser_10_reg
			       ,input [31:0] wr_resp_desc_c_xuser_11_reg
			       ,input [31:0] wr_resp_desc_c_xuser_12_reg
			       ,input [31:0] wr_resp_desc_c_xuser_13_reg
			       ,input [31:0] wr_resp_desc_c_xuser_14_reg
			       ,input [31:0] wr_resp_desc_c_xuser_15_reg
			       ,input [31:0] sn_req_desc_c_attr_reg
			       ,input [31:0] sn_req_desc_c_acaddr_0_reg
			       ,input [31:0] sn_req_desc_c_acaddr_1_reg
			       ,input [31:0] sn_req_desc_c_acaddr_2_reg
			       ,input [31:0] sn_req_desc_c_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_c_resp_reg
			       ,input [31:0] rd_req_desc_d_txn_type_reg
			       ,input [31:0] rd_req_desc_d_size_reg
			       ,input [31:0] rd_req_desc_d_axsize_reg
			       ,input [31:0] rd_req_desc_d_attr_reg
			       ,input [31:0] rd_req_desc_d_axaddr_0_reg
			       ,input [31:0] rd_req_desc_d_axaddr_1_reg
			       ,input [31:0] rd_req_desc_d_axaddr_2_reg
			       ,input [31:0] rd_req_desc_d_axaddr_3_reg
			       ,input [31:0] rd_req_desc_d_axid_0_reg
			       ,input [31:0] rd_req_desc_d_axid_1_reg
			       ,input [31:0] rd_req_desc_d_axid_2_reg
			       ,input [31:0] rd_req_desc_d_axid_3_reg
			       ,input [31:0] rd_req_desc_d_axuser_0_reg
			       ,input [31:0] rd_req_desc_d_axuser_1_reg
			       ,input [31:0] rd_req_desc_d_axuser_2_reg
			       ,input [31:0] rd_req_desc_d_axuser_3_reg
			       ,input [31:0] rd_req_desc_d_axuser_4_reg
			       ,input [31:0] rd_req_desc_d_axuser_5_reg
			       ,input [31:0] rd_req_desc_d_axuser_6_reg
			       ,input [31:0] rd_req_desc_d_axuser_7_reg
			       ,input [31:0] rd_req_desc_d_axuser_8_reg
			       ,input [31:0] rd_req_desc_d_axuser_9_reg
			       ,input [31:0] rd_req_desc_d_axuser_10_reg
			       ,input [31:0] rd_req_desc_d_axuser_11_reg
			       ,input [31:0] rd_req_desc_d_axuser_12_reg
			       ,input [31:0] rd_req_desc_d_axuser_13_reg
			       ,input [31:0] rd_req_desc_d_axuser_14_reg
			       ,input [31:0] rd_req_desc_d_axuser_15_reg
			       ,input [31:0] rd_resp_desc_d_data_offset_reg
			       ,input [31:0] rd_resp_desc_d_data_size_reg
			       ,input [31:0] rd_resp_desc_d_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_d_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_d_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_d_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_d_resp_reg
			       ,input [31:0] rd_resp_desc_d_xid_0_reg
			       ,input [31:0] rd_resp_desc_d_xid_1_reg
			       ,input [31:0] rd_resp_desc_d_xid_2_reg
			       ,input [31:0] rd_resp_desc_d_xid_3_reg
			       ,input [31:0] rd_resp_desc_d_xuser_0_reg
			       ,input [31:0] rd_resp_desc_d_xuser_1_reg
			       ,input [31:0] rd_resp_desc_d_xuser_2_reg
			       ,input [31:0] rd_resp_desc_d_xuser_3_reg
			       ,input [31:0] rd_resp_desc_d_xuser_4_reg
			       ,input [31:0] rd_resp_desc_d_xuser_5_reg
			       ,input [31:0] rd_resp_desc_d_xuser_6_reg
			       ,input [31:0] rd_resp_desc_d_xuser_7_reg
			       ,input [31:0] rd_resp_desc_d_xuser_8_reg
			       ,input [31:0] rd_resp_desc_d_xuser_9_reg
			       ,input [31:0] rd_resp_desc_d_xuser_10_reg
			       ,input [31:0] rd_resp_desc_d_xuser_11_reg
			       ,input [31:0] rd_resp_desc_d_xuser_12_reg
			       ,input [31:0] rd_resp_desc_d_xuser_13_reg
			       ,input [31:0] rd_resp_desc_d_xuser_14_reg
			       ,input [31:0] rd_resp_desc_d_xuser_15_reg
			       ,input [31:0] wr_req_desc_d_txn_type_reg
			       ,input [31:0] wr_req_desc_d_size_reg
			       ,input [31:0] wr_req_desc_d_data_offset_reg
			       ,input [31:0] wr_req_desc_d_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_d_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_d_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_d_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_d_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_d_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_d_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_d_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_d_axsize_reg
			       ,input [31:0] wr_req_desc_d_attr_reg
			       ,input [31:0] wr_req_desc_d_axaddr_0_reg
			       ,input [31:0] wr_req_desc_d_axaddr_1_reg
			       ,input [31:0] wr_req_desc_d_axaddr_2_reg
			       ,input [31:0] wr_req_desc_d_axaddr_3_reg
			       ,input [31:0] wr_req_desc_d_axid_0_reg
			       ,input [31:0] wr_req_desc_d_axid_1_reg
			       ,input [31:0] wr_req_desc_d_axid_2_reg
			       ,input [31:0] wr_req_desc_d_axid_3_reg
			       ,input [31:0] wr_req_desc_d_axuser_0_reg
			       ,input [31:0] wr_req_desc_d_axuser_1_reg
			       ,input [31:0] wr_req_desc_d_axuser_2_reg
			       ,input [31:0] wr_req_desc_d_axuser_3_reg
			       ,input [31:0] wr_req_desc_d_axuser_4_reg
			       ,input [31:0] wr_req_desc_d_axuser_5_reg
			       ,input [31:0] wr_req_desc_d_axuser_6_reg
			       ,input [31:0] wr_req_desc_d_axuser_7_reg
			       ,input [31:0] wr_req_desc_d_axuser_8_reg
			       ,input [31:0] wr_req_desc_d_axuser_9_reg
			       ,input [31:0] wr_req_desc_d_axuser_10_reg
			       ,input [31:0] wr_req_desc_d_axuser_11_reg
			       ,input [31:0] wr_req_desc_d_axuser_12_reg
			       ,input [31:0] wr_req_desc_d_axuser_13_reg
			       ,input [31:0] wr_req_desc_d_axuser_14_reg
			       ,input [31:0] wr_req_desc_d_axuser_15_reg
			       ,input [31:0] wr_req_desc_d_wuser_0_reg
			       ,input [31:0] wr_req_desc_d_wuser_1_reg
			       ,input [31:0] wr_req_desc_d_wuser_2_reg
			       ,input [31:0] wr_req_desc_d_wuser_3_reg
			       ,input [31:0] wr_req_desc_d_wuser_4_reg
			       ,input [31:0] wr_req_desc_d_wuser_5_reg
			       ,input [31:0] wr_req_desc_d_wuser_6_reg
			       ,input [31:0] wr_req_desc_d_wuser_7_reg
			       ,input [31:0] wr_req_desc_d_wuser_8_reg
			       ,input [31:0] wr_req_desc_d_wuser_9_reg
			       ,input [31:0] wr_req_desc_d_wuser_10_reg
			       ,input [31:0] wr_req_desc_d_wuser_11_reg
			       ,input [31:0] wr_req_desc_d_wuser_12_reg
			       ,input [31:0] wr_req_desc_d_wuser_13_reg
			       ,input [31:0] wr_req_desc_d_wuser_14_reg
			       ,input [31:0] wr_req_desc_d_wuser_15_reg
			       ,input [31:0] wr_resp_desc_d_resp_reg
			       ,input [31:0] wr_resp_desc_d_xid_0_reg
			       ,input [31:0] wr_resp_desc_d_xid_1_reg
			       ,input [31:0] wr_resp_desc_d_xid_2_reg
			       ,input [31:0] wr_resp_desc_d_xid_3_reg
			       ,input [31:0] wr_resp_desc_d_xuser_0_reg
			       ,input [31:0] wr_resp_desc_d_xuser_1_reg
			       ,input [31:0] wr_resp_desc_d_xuser_2_reg
			       ,input [31:0] wr_resp_desc_d_xuser_3_reg
			       ,input [31:0] wr_resp_desc_d_xuser_4_reg
			       ,input [31:0] wr_resp_desc_d_xuser_5_reg
			       ,input [31:0] wr_resp_desc_d_xuser_6_reg
			       ,input [31:0] wr_resp_desc_d_xuser_7_reg
			       ,input [31:0] wr_resp_desc_d_xuser_8_reg
			       ,input [31:0] wr_resp_desc_d_xuser_9_reg
			       ,input [31:0] wr_resp_desc_d_xuser_10_reg
			       ,input [31:0] wr_resp_desc_d_xuser_11_reg
			       ,input [31:0] wr_resp_desc_d_xuser_12_reg
			       ,input [31:0] wr_resp_desc_d_xuser_13_reg
			       ,input [31:0] wr_resp_desc_d_xuser_14_reg
			       ,input [31:0] wr_resp_desc_d_xuser_15_reg
			       ,input [31:0] sn_req_desc_d_attr_reg
			       ,input [31:0] sn_req_desc_d_acaddr_0_reg
			       ,input [31:0] sn_req_desc_d_acaddr_1_reg
			       ,input [31:0] sn_req_desc_d_acaddr_2_reg
			       ,input [31:0] sn_req_desc_d_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_d_resp_reg
			       ,input [31:0] rd_req_desc_e_txn_type_reg
			       ,input [31:0] rd_req_desc_e_size_reg
			       ,input [31:0] rd_req_desc_e_axsize_reg
			       ,input [31:0] rd_req_desc_e_attr_reg
			       ,input [31:0] rd_req_desc_e_axaddr_0_reg
			       ,input [31:0] rd_req_desc_e_axaddr_1_reg
			       ,input [31:0] rd_req_desc_e_axaddr_2_reg
			       ,input [31:0] rd_req_desc_e_axaddr_3_reg
			       ,input [31:0] rd_req_desc_e_axid_0_reg
			       ,input [31:0] rd_req_desc_e_axid_1_reg
			       ,input [31:0] rd_req_desc_e_axid_2_reg
			       ,input [31:0] rd_req_desc_e_axid_3_reg
			       ,input [31:0] rd_req_desc_e_axuser_0_reg
			       ,input [31:0] rd_req_desc_e_axuser_1_reg
			       ,input [31:0] rd_req_desc_e_axuser_2_reg
			       ,input [31:0] rd_req_desc_e_axuser_3_reg
			       ,input [31:0] rd_req_desc_e_axuser_4_reg
			       ,input [31:0] rd_req_desc_e_axuser_5_reg
			       ,input [31:0] rd_req_desc_e_axuser_6_reg
			       ,input [31:0] rd_req_desc_e_axuser_7_reg
			       ,input [31:0] rd_req_desc_e_axuser_8_reg
			       ,input [31:0] rd_req_desc_e_axuser_9_reg
			       ,input [31:0] rd_req_desc_e_axuser_10_reg
			       ,input [31:0] rd_req_desc_e_axuser_11_reg
			       ,input [31:0] rd_req_desc_e_axuser_12_reg
			       ,input [31:0] rd_req_desc_e_axuser_13_reg
			       ,input [31:0] rd_req_desc_e_axuser_14_reg
			       ,input [31:0] rd_req_desc_e_axuser_15_reg
			       ,input [31:0] rd_resp_desc_e_data_offset_reg
			       ,input [31:0] rd_resp_desc_e_data_size_reg
			       ,input [31:0] rd_resp_desc_e_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_e_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_e_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_e_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_e_resp_reg
			       ,input [31:0] rd_resp_desc_e_xid_0_reg
			       ,input [31:0] rd_resp_desc_e_xid_1_reg
			       ,input [31:0] rd_resp_desc_e_xid_2_reg
			       ,input [31:0] rd_resp_desc_e_xid_3_reg
			       ,input [31:0] rd_resp_desc_e_xuser_0_reg
			       ,input [31:0] rd_resp_desc_e_xuser_1_reg
			       ,input [31:0] rd_resp_desc_e_xuser_2_reg
			       ,input [31:0] rd_resp_desc_e_xuser_3_reg
			       ,input [31:0] rd_resp_desc_e_xuser_4_reg
			       ,input [31:0] rd_resp_desc_e_xuser_5_reg
			       ,input [31:0] rd_resp_desc_e_xuser_6_reg
			       ,input [31:0] rd_resp_desc_e_xuser_7_reg
			       ,input [31:0] rd_resp_desc_e_xuser_8_reg
			       ,input [31:0] rd_resp_desc_e_xuser_9_reg
			       ,input [31:0] rd_resp_desc_e_xuser_10_reg
			       ,input [31:0] rd_resp_desc_e_xuser_11_reg
			       ,input [31:0] rd_resp_desc_e_xuser_12_reg
			       ,input [31:0] rd_resp_desc_e_xuser_13_reg
			       ,input [31:0] rd_resp_desc_e_xuser_14_reg
			       ,input [31:0] rd_resp_desc_e_xuser_15_reg
			       ,input [31:0] wr_req_desc_e_txn_type_reg
			       ,input [31:0] wr_req_desc_e_size_reg
			       ,input [31:0] wr_req_desc_e_data_offset_reg
			       ,input [31:0] wr_req_desc_e_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_e_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_e_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_e_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_e_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_e_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_e_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_e_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_e_axsize_reg
			       ,input [31:0] wr_req_desc_e_attr_reg
			       ,input [31:0] wr_req_desc_e_axaddr_0_reg
			       ,input [31:0] wr_req_desc_e_axaddr_1_reg
			       ,input [31:0] wr_req_desc_e_axaddr_2_reg
			       ,input [31:0] wr_req_desc_e_axaddr_3_reg
			       ,input [31:0] wr_req_desc_e_axid_0_reg
			       ,input [31:0] wr_req_desc_e_axid_1_reg
			       ,input [31:0] wr_req_desc_e_axid_2_reg
			       ,input [31:0] wr_req_desc_e_axid_3_reg
			       ,input [31:0] wr_req_desc_e_axuser_0_reg
			       ,input [31:0] wr_req_desc_e_axuser_1_reg
			       ,input [31:0] wr_req_desc_e_axuser_2_reg
			       ,input [31:0] wr_req_desc_e_axuser_3_reg
			       ,input [31:0] wr_req_desc_e_axuser_4_reg
			       ,input [31:0] wr_req_desc_e_axuser_5_reg
			       ,input [31:0] wr_req_desc_e_axuser_6_reg
			       ,input [31:0] wr_req_desc_e_axuser_7_reg
			       ,input [31:0] wr_req_desc_e_axuser_8_reg
			       ,input [31:0] wr_req_desc_e_axuser_9_reg
			       ,input [31:0] wr_req_desc_e_axuser_10_reg
			       ,input [31:0] wr_req_desc_e_axuser_11_reg
			       ,input [31:0] wr_req_desc_e_axuser_12_reg
			       ,input [31:0] wr_req_desc_e_axuser_13_reg
			       ,input [31:0] wr_req_desc_e_axuser_14_reg
			       ,input [31:0] wr_req_desc_e_axuser_15_reg
			       ,input [31:0] wr_req_desc_e_wuser_0_reg
			       ,input [31:0] wr_req_desc_e_wuser_1_reg
			       ,input [31:0] wr_req_desc_e_wuser_2_reg
			       ,input [31:0] wr_req_desc_e_wuser_3_reg
			       ,input [31:0] wr_req_desc_e_wuser_4_reg
			       ,input [31:0] wr_req_desc_e_wuser_5_reg
			       ,input [31:0] wr_req_desc_e_wuser_6_reg
			       ,input [31:0] wr_req_desc_e_wuser_7_reg
			       ,input [31:0] wr_req_desc_e_wuser_8_reg
			       ,input [31:0] wr_req_desc_e_wuser_9_reg
			       ,input [31:0] wr_req_desc_e_wuser_10_reg
			       ,input [31:0] wr_req_desc_e_wuser_11_reg
			       ,input [31:0] wr_req_desc_e_wuser_12_reg
			       ,input [31:0] wr_req_desc_e_wuser_13_reg
			       ,input [31:0] wr_req_desc_e_wuser_14_reg
			       ,input [31:0] wr_req_desc_e_wuser_15_reg
			       ,input [31:0] wr_resp_desc_e_resp_reg
			       ,input [31:0] wr_resp_desc_e_xid_0_reg
			       ,input [31:0] wr_resp_desc_e_xid_1_reg
			       ,input [31:0] wr_resp_desc_e_xid_2_reg
			       ,input [31:0] wr_resp_desc_e_xid_3_reg
			       ,input [31:0] wr_resp_desc_e_xuser_0_reg
			       ,input [31:0] wr_resp_desc_e_xuser_1_reg
			       ,input [31:0] wr_resp_desc_e_xuser_2_reg
			       ,input [31:0] wr_resp_desc_e_xuser_3_reg
			       ,input [31:0] wr_resp_desc_e_xuser_4_reg
			       ,input [31:0] wr_resp_desc_e_xuser_5_reg
			       ,input [31:0] wr_resp_desc_e_xuser_6_reg
			       ,input [31:0] wr_resp_desc_e_xuser_7_reg
			       ,input [31:0] wr_resp_desc_e_xuser_8_reg
			       ,input [31:0] wr_resp_desc_e_xuser_9_reg
			       ,input [31:0] wr_resp_desc_e_xuser_10_reg
			       ,input [31:0] wr_resp_desc_e_xuser_11_reg
			       ,input [31:0] wr_resp_desc_e_xuser_12_reg
			       ,input [31:0] wr_resp_desc_e_xuser_13_reg
			       ,input [31:0] wr_resp_desc_e_xuser_14_reg
			       ,input [31:0] wr_resp_desc_e_xuser_15_reg
			       ,input [31:0] sn_req_desc_e_attr_reg
			       ,input [31:0] sn_req_desc_e_acaddr_0_reg
			       ,input [31:0] sn_req_desc_e_acaddr_1_reg
			       ,input [31:0] sn_req_desc_e_acaddr_2_reg
			       ,input [31:0] sn_req_desc_e_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_e_resp_reg
			       ,input [31:0] rd_req_desc_f_txn_type_reg
			       ,input [31:0] rd_req_desc_f_size_reg
			       ,input [31:0] rd_req_desc_f_axsize_reg
			       ,input [31:0] rd_req_desc_f_attr_reg
			       ,input [31:0] rd_req_desc_f_axaddr_0_reg
			       ,input [31:0] rd_req_desc_f_axaddr_1_reg
			       ,input [31:0] rd_req_desc_f_axaddr_2_reg
			       ,input [31:0] rd_req_desc_f_axaddr_3_reg
			       ,input [31:0] rd_req_desc_f_axid_0_reg
			       ,input [31:0] rd_req_desc_f_axid_1_reg
			       ,input [31:0] rd_req_desc_f_axid_2_reg
			       ,input [31:0] rd_req_desc_f_axid_3_reg
			       ,input [31:0] rd_req_desc_f_axuser_0_reg
			       ,input [31:0] rd_req_desc_f_axuser_1_reg
			       ,input [31:0] rd_req_desc_f_axuser_2_reg
			       ,input [31:0] rd_req_desc_f_axuser_3_reg
			       ,input [31:0] rd_req_desc_f_axuser_4_reg
			       ,input [31:0] rd_req_desc_f_axuser_5_reg
			       ,input [31:0] rd_req_desc_f_axuser_6_reg
			       ,input [31:0] rd_req_desc_f_axuser_7_reg
			       ,input [31:0] rd_req_desc_f_axuser_8_reg
			       ,input [31:0] rd_req_desc_f_axuser_9_reg
			       ,input [31:0] rd_req_desc_f_axuser_10_reg
			       ,input [31:0] rd_req_desc_f_axuser_11_reg
			       ,input [31:0] rd_req_desc_f_axuser_12_reg
			       ,input [31:0] rd_req_desc_f_axuser_13_reg
			       ,input [31:0] rd_req_desc_f_axuser_14_reg
			       ,input [31:0] rd_req_desc_f_axuser_15_reg
			       ,input [31:0] rd_resp_desc_f_data_offset_reg
			       ,input [31:0] rd_resp_desc_f_data_size_reg
			       ,input [31:0] rd_resp_desc_f_data_host_addr_0_reg
			       ,input [31:0] rd_resp_desc_f_data_host_addr_1_reg
			       ,input [31:0] rd_resp_desc_f_data_host_addr_2_reg
			       ,input [31:0] rd_resp_desc_f_data_host_addr_3_reg
			       ,input [31:0] rd_resp_desc_f_resp_reg
			       ,input [31:0] rd_resp_desc_f_xid_0_reg
			       ,input [31:0] rd_resp_desc_f_xid_1_reg
			       ,input [31:0] rd_resp_desc_f_xid_2_reg
			       ,input [31:0] rd_resp_desc_f_xid_3_reg
			       ,input [31:0] rd_resp_desc_f_xuser_0_reg
			       ,input [31:0] rd_resp_desc_f_xuser_1_reg
			       ,input [31:0] rd_resp_desc_f_xuser_2_reg
			       ,input [31:0] rd_resp_desc_f_xuser_3_reg
			       ,input [31:0] rd_resp_desc_f_xuser_4_reg
			       ,input [31:0] rd_resp_desc_f_xuser_5_reg
			       ,input [31:0] rd_resp_desc_f_xuser_6_reg
			       ,input [31:0] rd_resp_desc_f_xuser_7_reg
			       ,input [31:0] rd_resp_desc_f_xuser_8_reg
			       ,input [31:0] rd_resp_desc_f_xuser_9_reg
			       ,input [31:0] rd_resp_desc_f_xuser_10_reg
			       ,input [31:0] rd_resp_desc_f_xuser_11_reg
			       ,input [31:0] rd_resp_desc_f_xuser_12_reg
			       ,input [31:0] rd_resp_desc_f_xuser_13_reg
			       ,input [31:0] rd_resp_desc_f_xuser_14_reg
			       ,input [31:0] rd_resp_desc_f_xuser_15_reg
			       ,input [31:0] wr_req_desc_f_txn_type_reg
			       ,input [31:0] wr_req_desc_f_size_reg
			       ,input [31:0] wr_req_desc_f_data_offset_reg
			       ,input [31:0] wr_req_desc_f_data_host_addr_0_reg
			       ,input [31:0] wr_req_desc_f_data_host_addr_1_reg
			       ,input [31:0] wr_req_desc_f_data_host_addr_2_reg
			       ,input [31:0] wr_req_desc_f_data_host_addr_3_reg
			       ,input [31:0] wr_req_desc_f_wstrb_host_addr_0_reg
			       ,input [31:0] wr_req_desc_f_wstrb_host_addr_1_reg
			       ,input [31:0] wr_req_desc_f_wstrb_host_addr_2_reg
			       ,input [31:0] wr_req_desc_f_wstrb_host_addr_3_reg
			       ,input [31:0] wr_req_desc_f_axsize_reg
			       ,input [31:0] wr_req_desc_f_attr_reg
			       ,input [31:0] wr_req_desc_f_axaddr_0_reg
			       ,input [31:0] wr_req_desc_f_axaddr_1_reg
			       ,input [31:0] wr_req_desc_f_axaddr_2_reg
			       ,input [31:0] wr_req_desc_f_axaddr_3_reg
			       ,input [31:0] wr_req_desc_f_axid_0_reg
			       ,input [31:0] wr_req_desc_f_axid_1_reg
			       ,input [31:0] wr_req_desc_f_axid_2_reg
			       ,input [31:0] wr_req_desc_f_axid_3_reg
			       ,input [31:0] wr_req_desc_f_axuser_0_reg
			       ,input [31:0] wr_req_desc_f_axuser_1_reg
			       ,input [31:0] wr_req_desc_f_axuser_2_reg
			       ,input [31:0] wr_req_desc_f_axuser_3_reg
			       ,input [31:0] wr_req_desc_f_axuser_4_reg
			       ,input [31:0] wr_req_desc_f_axuser_5_reg
			       ,input [31:0] wr_req_desc_f_axuser_6_reg
			       ,input [31:0] wr_req_desc_f_axuser_7_reg
			       ,input [31:0] wr_req_desc_f_axuser_8_reg
			       ,input [31:0] wr_req_desc_f_axuser_9_reg
			       ,input [31:0] wr_req_desc_f_axuser_10_reg
			       ,input [31:0] wr_req_desc_f_axuser_11_reg
			       ,input [31:0] wr_req_desc_f_axuser_12_reg
			       ,input [31:0] wr_req_desc_f_axuser_13_reg
			       ,input [31:0] wr_req_desc_f_axuser_14_reg
			       ,input [31:0] wr_req_desc_f_axuser_15_reg
			       ,input [31:0] wr_req_desc_f_wuser_0_reg
			       ,input [31:0] wr_req_desc_f_wuser_1_reg
			       ,input [31:0] wr_req_desc_f_wuser_2_reg
			       ,input [31:0] wr_req_desc_f_wuser_3_reg
			       ,input [31:0] wr_req_desc_f_wuser_4_reg
			       ,input [31:0] wr_req_desc_f_wuser_5_reg
			       ,input [31:0] wr_req_desc_f_wuser_6_reg
			       ,input [31:0] wr_req_desc_f_wuser_7_reg
			       ,input [31:0] wr_req_desc_f_wuser_8_reg
			       ,input [31:0] wr_req_desc_f_wuser_9_reg
			       ,input [31:0] wr_req_desc_f_wuser_10_reg
			       ,input [31:0] wr_req_desc_f_wuser_11_reg
			       ,input [31:0] wr_req_desc_f_wuser_12_reg
			       ,input [31:0] wr_req_desc_f_wuser_13_reg
			       ,input [31:0] wr_req_desc_f_wuser_14_reg
			       ,input [31:0] wr_req_desc_f_wuser_15_reg
			       ,input [31:0] wr_resp_desc_f_resp_reg
			       ,input [31:0] wr_resp_desc_f_xid_0_reg
			       ,input [31:0] wr_resp_desc_f_xid_1_reg
			       ,input [31:0] wr_resp_desc_f_xid_2_reg
			       ,input [31:0] wr_resp_desc_f_xid_3_reg
			       ,input [31:0] wr_resp_desc_f_xuser_0_reg
			       ,input [31:0] wr_resp_desc_f_xuser_1_reg
			       ,input [31:0] wr_resp_desc_f_xuser_2_reg
			       ,input [31:0] wr_resp_desc_f_xuser_3_reg
			       ,input [31:0] wr_resp_desc_f_xuser_4_reg
			       ,input [31:0] wr_resp_desc_f_xuser_5_reg
			       ,input [31:0] wr_resp_desc_f_xuser_6_reg
			       ,input [31:0] wr_resp_desc_f_xuser_7_reg
			       ,input [31:0] wr_resp_desc_f_xuser_8_reg
			       ,input [31:0] wr_resp_desc_f_xuser_9_reg
			       ,input [31:0] wr_resp_desc_f_xuser_10_reg
			       ,input [31:0] wr_resp_desc_f_xuser_11_reg
			       ,input [31:0] wr_resp_desc_f_xuser_12_reg
			       ,input [31:0] wr_resp_desc_f_xuser_13_reg
			       ,input [31:0] wr_resp_desc_f_xuser_14_reg
			       ,input [31:0] wr_resp_desc_f_xuser_15_reg
			       ,input [31:0] sn_req_desc_f_attr_reg
			       ,input [31:0] sn_req_desc_f_acaddr_0_reg
			       ,input [31:0] sn_req_desc_f_acaddr_1_reg
			       ,input [31:0] sn_req_desc_f_acaddr_2_reg
			       ,input [31:0] sn_req_desc_f_acaddr_3_reg
			       ,input [31:0] sn_resp_desc_f_resp_reg
   
   
			       ,output [31:0] uc2rb_intr_error_status_reg
			       ,output [31:0] uc2rb_rd_req_fifo_free_level_reg
			       ,output [31:0] uc2rb_rd_req_intr_comp_status_reg
			       ,output [31:0] uc2rb_rd_resp_fifo_pop_desc_reg
			       ,output [31:0] uc2rb_rd_resp_fifo_fill_level_reg
			       ,output [31:0] uc2rb_wr_req_fifo_free_level_reg
			       ,output [31:0] uc2rb_wr_req_intr_comp_status_reg
			       ,output [31:0] uc2rb_wr_resp_fifo_pop_desc_reg
			       ,output [31:0] uc2rb_wr_resp_fifo_fill_level_reg
			       ,output [31:0] uc2rb_sn_req_fifo_pop_desc_reg
			       ,output [31:0] uc2rb_sn_req_fifo_fill_level_reg
			       ,output [31:0] uc2rb_sn_resp_fifo_free_level_reg
			       ,output [31:0] uc2rb_sn_resp_intr_comp_status_reg
			       ,output [31:0] uc2rb_sn_data_fifo_free_level_reg
			       ,output [31:0] uc2rb_sn_data_intr_comp_status_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_0_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_1_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_2_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_3_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_4_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_5_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_6_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_7_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_8_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_9_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_a_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_b_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_c_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_d_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_e_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_data_offset_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_data_size_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_resp_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_0_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_1_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_2_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_3_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_4_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_5_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_6_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_7_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_8_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_9_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_10_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_11_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_12_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_13_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_14_reg
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_15_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_resp_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_0_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_1_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_2_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_3_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_4_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_5_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_6_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_7_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_8_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_9_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_10_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_11_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_12_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_13_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_14_reg
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_15_reg
			       ,output [31:0] uc2rb_sn_req_desc_f_attr_reg
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_0_reg
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_1_reg
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_2_reg
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_3_reg
   
   
			       ,output [31:0] uc2rb_intr_error_status_reg_we
			       ,output [31:0] uc2rb_rd_req_fifo_free_level_reg_we
			       ,output [31:0] uc2rb_rd_req_intr_comp_status_reg_we
			       ,output [31:0] uc2rb_rd_resp_fifo_pop_desc_reg_we
			       ,output [31:0] uc2rb_rd_resp_fifo_fill_level_reg_we
			       ,output [31:0] uc2rb_wr_req_fifo_free_level_reg_we
			       ,output [31:0] uc2rb_wr_req_intr_comp_status_reg_we
			       ,output [31:0] uc2rb_wr_resp_fifo_pop_desc_reg_we
			       ,output [31:0] uc2rb_wr_resp_fifo_fill_level_reg_we
			       ,output [31:0] uc2rb_sn_req_fifo_pop_desc_reg_we
			       ,output [31:0] uc2rb_sn_req_fifo_fill_level_reg_we
			       ,output [31:0] uc2rb_sn_resp_fifo_free_level_reg_we
			       ,output [31:0] uc2rb_sn_resp_intr_comp_status_reg_we
			       ,output [31:0] uc2rb_sn_data_fifo_free_level_reg_we
			       ,output [31:0] uc2rb_sn_data_intr_comp_status_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_0_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_0_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_0_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_0_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_1_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_1_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_1_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_1_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_2_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_2_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_2_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_2_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_3_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_3_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_3_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_3_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_4_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_4_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_4_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_4_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_5_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_5_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_5_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_5_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_6_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_6_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_6_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_6_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_7_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_7_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_7_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_7_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_8_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_8_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_8_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_8_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_9_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_9_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_9_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_9_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_a_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_a_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_a_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_a_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_b_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_b_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_b_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_b_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_c_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_c_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_c_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_c_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_d_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_d_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_d_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_d_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_e_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_e_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_e_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_e_acaddr_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_data_offset_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_data_size_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_resp_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xid_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_0_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_1_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_2_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_3_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_4_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_5_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_6_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_7_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_8_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_9_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_10_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_11_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_12_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_13_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_14_reg_we
			       ,output [31:0] uc2rb_rd_resp_desc_f_xuser_15_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_resp_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xid_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_0_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_1_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_2_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_3_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_4_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_5_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_6_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_7_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_8_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_9_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_10_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_11_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_12_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_13_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_14_reg_we
			       ,output [31:0] uc2rb_wr_resp_desc_f_xuser_15_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_f_attr_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_0_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_1_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_2_reg_we
			       ,output [31:0] uc2rb_sn_req_desc_f_acaddr_3_reg_we
   
   
   
			       //RAM commands  
			       //RDATA_RAM
			       ,output uc2rb_wr_we 
			       ,output [(M_ACE_USR_XX_DATA_WIDTH/8)-1:0] uc2rb_wr_bwe //Generate all 1s always.     
			       ,output [(`CLOG2((XX_RAM_SIZE*8)/M_ACE_USR_XX_DATA_WIDTH))-1:0] uc2rb_wr_addr 
			       ,output [M_ACE_USR_XX_DATA_WIDTH-1:0] uc2rb_wr_data 
   
			       //WDATA_RAM and WSTRB_RAM                               
			       ,output [(`CLOG2((XX_RAM_SIZE*8)/M_ACE_USR_XX_DATA_WIDTH))-1:0] uc2rb_rd_addr 
			       ,input [M_ACE_USR_XX_DATA_WIDTH-1:0] rb2uc_rd_data 
			       ,input [(M_ACE_USR_XX_DATA_WIDTH/8)-1:0] rb2uc_rd_wstrb
   
			       //CDDATA_RAM                               
			       ,output [(`CLOG2((SN_RAM_SIZE*8)/M_ACE_USR_SN_DATA_WIDTH))-1:0] uc2rb_sn_addr 
			       ,input [M_ACE_USR_SN_DATA_WIDTH-1:0] rb2uc_sn_data 
   
			       ,output [XX_MAX_DESC-1:0] rd_uc2hm_trig 
			       ,input [XX_MAX_DESC-1:0] rd_hm2uc_done
			       ,output [XX_MAX_DESC-1:0] wr_uc2hm_trig 
			       ,input [XX_MAX_DESC-1:0] wr_hm2uc_done
   
			       //pop request to FIFO
			       ,input rd_resp_fifo_pop_desc_conn 
			       ,input wr_resp_fifo_pop_desc_conn 
			       ,input sn_req_fifo_pop_desc_conn
   
			       //output from FIFO
			       ,output [(`CLOG2(XX_MAX_DESC))-1:0] rd_resp_fifo_out
			       ,output rd_resp_fifo_out_valid //it is one clock cycle pulse
			       ,output [(`CLOG2(XX_MAX_DESC))-1:0] wr_resp_fifo_out
			       ,output wr_resp_fifo_out_valid //it is one clock cycle pulse
			       ,output [(`CLOG2(SN_MAX_DESC))-1:0] sn_req_fifo_out
			       ,output sn_req_fifo_out_valid  //it is one clock cycle pulse

			       );
   
   localparam XX_DESC_IDX_WIDTH                            = `CLOG2(XX_MAX_DESC);
   localparam XX_RAM_OFFSET_WIDTH                          = `CLOG2((XX_RAM_SIZE*8)/M_ACE_USR_XX_DATA_WIDTH);

   localparam ADDR_WIDTH                                   = M_ACE_USR_ADDR_WIDTH; 
   localparam XX_DATA_WIDTH                                = M_ACE_USR_XX_DATA_WIDTH; 
   localparam SN_DATA_WIDTH                                = M_ACE_USR_SN_DATA_WIDTH; 
   localparam ID_WIDTH                                     = M_ACE_USR_ID_WIDTH;   
   localparam AWUSER_WIDTH                                 = M_ACE_USR_AWUSER_WIDTH; 
   localparam WUSER_WIDTH                                  = M_ACE_USR_WUSER_WIDTH; 
   localparam BUSER_WIDTH                                  = M_ACE_USR_BUSER_WIDTH; 
   localparam ARUSER_WIDTH                                 = M_ACE_USR_ARUSER_WIDTH; 
   localparam RUSER_WIDTH                                  = M_ACE_USR_RUSER_WIDTH; 


   ace_usr_mst_control_field #(
			       /*AUTOINSTPARAM*/
                               // Parameters
                               .ACE_PROTOCOL       (ACE_PROTOCOL),
                               .ADDR_WIDTH         (ADDR_WIDTH),
                               .XX_DATA_WIDTH      (XX_DATA_WIDTH),
                               .SN_DATA_WIDTH      (SN_DATA_WIDTH),
                               .ID_WIDTH           (ID_WIDTH),
                               .AWUSER_WIDTH       (AWUSER_WIDTH),
                               .WUSER_WIDTH        (WUSER_WIDTH),
                               .BUSER_WIDTH        (BUSER_WIDTH),
                               .ARUSER_WIDTH       (ARUSER_WIDTH),
                               .RUSER_WIDTH        (RUSER_WIDTH),
                               .CACHE_LINE_SIZE    (CACHE_LINE_SIZE),
                               .XX_MAX_DESC        (XX_MAX_DESC),
                               .SN_MAX_DESC        (SN_MAX_DESC),
                               .XX_RAM_SIZE        (XX_RAM_SIZE),
                               .SN_RAM_SIZE        (SN_RAM_SIZE)) i_ace_usr_mst_control_field (
											       /*AUTOINST*/
                                                                                               // Outputs
                                                                                               .m_ace_usr_awid     (m_ace_usr_awid),
                                                                                               .m_ace_usr_awaddr   (m_ace_usr_awaddr),
                                                                                               .m_ace_usr_awlen    (m_ace_usr_awlen),
                                                                                               .m_ace_usr_awsize   (m_ace_usr_awsize),
                                                                                               .m_ace_usr_awburst  (m_ace_usr_awburst),
                                                                                               .m_ace_usr_awlock   (m_ace_usr_awlock),
                                                                                               .m_ace_usr_awcache  (m_ace_usr_awcache),
                                                                                               .m_ace_usr_awprot   (m_ace_usr_awprot),
                                                                                               .m_ace_usr_awqos    (m_ace_usr_awqos),
                                                                                               .m_ace_usr_awregion (m_ace_usr_awregion),
                                                                                               .m_ace_usr_awuser   (m_ace_usr_awuser),
                                                                                               .m_ace_usr_awsnoop  (m_ace_usr_awsnoop),
                                                                                               .m_ace_usr_awdomain (m_ace_usr_awdomain),
                                                                                               .m_ace_usr_awbar    (m_ace_usr_awbar),
                                                                                               .m_ace_usr_awunique (m_ace_usr_awunique),
                                                                                               .m_ace_usr_awvalid  (m_ace_usr_awvalid),
                                                                                               .m_ace_usr_wdata    (m_ace_usr_wdata),
                                                                                               .m_ace_usr_wstrb    (m_ace_usr_wstrb),
                                                                                               .m_ace_usr_wlast    (m_ace_usr_wlast),
                                                                                               .m_ace_usr_wuser    (m_ace_usr_wuser),
                                                                                               .m_ace_usr_wvalid   (m_ace_usr_wvalid),
                                                                                               .m_ace_usr_bready   (m_ace_usr_bready),
                                                                                               .m_ace_usr_wack     (m_ace_usr_wack),
                                                                                               .m_ace_usr_arid     (m_ace_usr_arid),
                                                                                               .m_ace_usr_araddr   (m_ace_usr_araddr),
                                                                                               .m_ace_usr_arlen    (m_ace_usr_arlen),
                                                                                               .m_ace_usr_arsize   (m_ace_usr_arsize),
                                                                                               .m_ace_usr_arburst  (m_ace_usr_arburst),
                                                                                               .m_ace_usr_arlock   (m_ace_usr_arlock),
                                                                                               .m_ace_usr_arcache  (m_ace_usr_arcache),
                                                                                               .m_ace_usr_arprot   (m_ace_usr_arprot),
                                                                                               .m_ace_usr_arqos    (m_ace_usr_arqos),
                                                                                               .m_ace_usr_arregion (m_ace_usr_arregion),
                                                                                               .m_ace_usr_aruser   (m_ace_usr_aruser),
                                                                                               .m_ace_usr_arsnoop  (m_ace_usr_arsnoop),
                                                                                               .m_ace_usr_ardomain (m_ace_usr_ardomain),
                                                                                               .m_ace_usr_arbar    (m_ace_usr_arbar),
                                                                                               .m_ace_usr_arvalid  (m_ace_usr_arvalid),
                                                                                               .m_ace_usr_rready   (m_ace_usr_rready),
                                                                                               .m_ace_usr_rack     (m_ace_usr_rack),
                                                                                               .m_ace_usr_acready  (m_ace_usr_acready),
                                                                                               .m_ace_usr_crresp   (m_ace_usr_crresp),
                                                                                               .m_ace_usr_crvalid  (m_ace_usr_crvalid),
                                                                                               .m_ace_usr_cddata   (m_ace_usr_cddata),
                                                                                               .m_ace_usr_cdlast   (m_ace_usr_cdlast),
                                                                                               .m_ace_usr_cdvalid  (m_ace_usr_cdvalid),
                                                                                               .uc2rb_intr_error_status_reg(uc2rb_intr_error_status_reg),
                                                                                               .uc2rb_rd_req_fifo_free_level_reg(uc2rb_rd_req_fifo_free_level_reg),
                                                                                               .uc2rb_rd_req_intr_comp_status_reg(uc2rb_rd_req_intr_comp_status_reg),
                                                                                               .uc2rb_rd_resp_fifo_pop_desc_reg(uc2rb_rd_resp_fifo_pop_desc_reg),
                                                                                               .uc2rb_rd_resp_fifo_fill_level_reg(uc2rb_rd_resp_fifo_fill_level_reg),
                                                                                               .uc2rb_wr_req_fifo_free_level_reg(uc2rb_wr_req_fifo_free_level_reg),
                                                                                               .uc2rb_wr_req_intr_comp_status_reg(uc2rb_wr_req_intr_comp_status_reg),
                                                                                               .uc2rb_wr_resp_fifo_pop_desc_reg(uc2rb_wr_resp_fifo_pop_desc_reg),
                                                                                               .uc2rb_wr_resp_fifo_fill_level_reg(uc2rb_wr_resp_fifo_fill_level_reg),
                                                                                               .uc2rb_sn_req_fifo_pop_desc_reg(uc2rb_sn_req_fifo_pop_desc_reg),
                                                                                               .uc2rb_sn_req_fifo_fill_level_reg(uc2rb_sn_req_fifo_fill_level_reg),
                                                                                               .uc2rb_sn_resp_fifo_free_level_reg(uc2rb_sn_resp_fifo_free_level_reg),
                                                                                               .uc2rb_sn_resp_intr_comp_status_reg(uc2rb_sn_resp_intr_comp_status_reg),
                                                                                               .uc2rb_sn_data_fifo_free_level_reg(uc2rb_sn_data_fifo_free_level_reg),
                                                                                               .uc2rb_sn_data_intr_comp_status_reg(uc2rb_sn_data_intr_comp_status_reg),
                                                                                               .uc2rb_rd_resp_desc_0_data_offset_reg(uc2rb_rd_resp_desc_0_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_0_data_size_reg(uc2rb_rd_resp_desc_0_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_0_resp_reg(uc2rb_rd_resp_desc_0_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xid_0_reg(uc2rb_rd_resp_desc_0_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xid_1_reg(uc2rb_rd_resp_desc_0_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xid_2_reg(uc2rb_rd_resp_desc_0_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xid_3_reg(uc2rb_rd_resp_desc_0_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_0_reg(uc2rb_rd_resp_desc_0_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_1_reg(uc2rb_rd_resp_desc_0_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_2_reg(uc2rb_rd_resp_desc_0_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_3_reg(uc2rb_rd_resp_desc_0_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_4_reg(uc2rb_rd_resp_desc_0_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_5_reg(uc2rb_rd_resp_desc_0_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_6_reg(uc2rb_rd_resp_desc_0_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_7_reg(uc2rb_rd_resp_desc_0_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_8_reg(uc2rb_rd_resp_desc_0_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_9_reg(uc2rb_rd_resp_desc_0_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_10_reg(uc2rb_rd_resp_desc_0_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_11_reg(uc2rb_rd_resp_desc_0_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_12_reg(uc2rb_rd_resp_desc_0_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_13_reg(uc2rb_rd_resp_desc_0_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_14_reg(uc2rb_rd_resp_desc_0_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_15_reg(uc2rb_rd_resp_desc_0_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_0_resp_reg(uc2rb_wr_resp_desc_0_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xid_0_reg(uc2rb_wr_resp_desc_0_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xid_1_reg(uc2rb_wr_resp_desc_0_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xid_2_reg(uc2rb_wr_resp_desc_0_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xid_3_reg(uc2rb_wr_resp_desc_0_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_0_reg(uc2rb_wr_resp_desc_0_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_1_reg(uc2rb_wr_resp_desc_0_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_2_reg(uc2rb_wr_resp_desc_0_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_3_reg(uc2rb_wr_resp_desc_0_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_4_reg(uc2rb_wr_resp_desc_0_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_5_reg(uc2rb_wr_resp_desc_0_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_6_reg(uc2rb_wr_resp_desc_0_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_7_reg(uc2rb_wr_resp_desc_0_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_8_reg(uc2rb_wr_resp_desc_0_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_9_reg(uc2rb_wr_resp_desc_0_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_10_reg(uc2rb_wr_resp_desc_0_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_11_reg(uc2rb_wr_resp_desc_0_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_12_reg(uc2rb_wr_resp_desc_0_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_13_reg(uc2rb_wr_resp_desc_0_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_14_reg(uc2rb_wr_resp_desc_0_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_15_reg(uc2rb_wr_resp_desc_0_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_0_attr_reg(uc2rb_sn_req_desc_0_attr_reg),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_0_reg(uc2rb_sn_req_desc_0_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_1_reg(uc2rb_sn_req_desc_0_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_2_reg(uc2rb_sn_req_desc_0_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_3_reg(uc2rb_sn_req_desc_0_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_1_data_offset_reg(uc2rb_rd_resp_desc_1_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_1_data_size_reg(uc2rb_rd_resp_desc_1_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_1_resp_reg(uc2rb_rd_resp_desc_1_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xid_0_reg(uc2rb_rd_resp_desc_1_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xid_1_reg(uc2rb_rd_resp_desc_1_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xid_2_reg(uc2rb_rd_resp_desc_1_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xid_3_reg(uc2rb_rd_resp_desc_1_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_0_reg(uc2rb_rd_resp_desc_1_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_1_reg(uc2rb_rd_resp_desc_1_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_2_reg(uc2rb_rd_resp_desc_1_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_3_reg(uc2rb_rd_resp_desc_1_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_4_reg(uc2rb_rd_resp_desc_1_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_5_reg(uc2rb_rd_resp_desc_1_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_6_reg(uc2rb_rd_resp_desc_1_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_7_reg(uc2rb_rd_resp_desc_1_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_8_reg(uc2rb_rd_resp_desc_1_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_9_reg(uc2rb_rd_resp_desc_1_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_10_reg(uc2rb_rd_resp_desc_1_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_11_reg(uc2rb_rd_resp_desc_1_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_12_reg(uc2rb_rd_resp_desc_1_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_13_reg(uc2rb_rd_resp_desc_1_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_14_reg(uc2rb_rd_resp_desc_1_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_15_reg(uc2rb_rd_resp_desc_1_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_1_resp_reg(uc2rb_wr_resp_desc_1_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xid_0_reg(uc2rb_wr_resp_desc_1_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xid_1_reg(uc2rb_wr_resp_desc_1_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xid_2_reg(uc2rb_wr_resp_desc_1_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xid_3_reg(uc2rb_wr_resp_desc_1_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_0_reg(uc2rb_wr_resp_desc_1_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_1_reg(uc2rb_wr_resp_desc_1_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_2_reg(uc2rb_wr_resp_desc_1_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_3_reg(uc2rb_wr_resp_desc_1_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_4_reg(uc2rb_wr_resp_desc_1_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_5_reg(uc2rb_wr_resp_desc_1_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_6_reg(uc2rb_wr_resp_desc_1_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_7_reg(uc2rb_wr_resp_desc_1_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_8_reg(uc2rb_wr_resp_desc_1_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_9_reg(uc2rb_wr_resp_desc_1_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_10_reg(uc2rb_wr_resp_desc_1_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_11_reg(uc2rb_wr_resp_desc_1_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_12_reg(uc2rb_wr_resp_desc_1_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_13_reg(uc2rb_wr_resp_desc_1_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_14_reg(uc2rb_wr_resp_desc_1_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_15_reg(uc2rb_wr_resp_desc_1_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_1_attr_reg(uc2rb_sn_req_desc_1_attr_reg),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_0_reg(uc2rb_sn_req_desc_1_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_1_reg(uc2rb_sn_req_desc_1_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_2_reg(uc2rb_sn_req_desc_1_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_3_reg(uc2rb_sn_req_desc_1_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_2_data_offset_reg(uc2rb_rd_resp_desc_2_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_2_data_size_reg(uc2rb_rd_resp_desc_2_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_2_resp_reg(uc2rb_rd_resp_desc_2_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xid_0_reg(uc2rb_rd_resp_desc_2_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xid_1_reg(uc2rb_rd_resp_desc_2_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xid_2_reg(uc2rb_rd_resp_desc_2_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xid_3_reg(uc2rb_rd_resp_desc_2_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_0_reg(uc2rb_rd_resp_desc_2_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_1_reg(uc2rb_rd_resp_desc_2_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_2_reg(uc2rb_rd_resp_desc_2_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_3_reg(uc2rb_rd_resp_desc_2_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_4_reg(uc2rb_rd_resp_desc_2_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_5_reg(uc2rb_rd_resp_desc_2_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_6_reg(uc2rb_rd_resp_desc_2_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_7_reg(uc2rb_rd_resp_desc_2_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_8_reg(uc2rb_rd_resp_desc_2_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_9_reg(uc2rb_rd_resp_desc_2_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_10_reg(uc2rb_rd_resp_desc_2_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_11_reg(uc2rb_rd_resp_desc_2_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_12_reg(uc2rb_rd_resp_desc_2_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_13_reg(uc2rb_rd_resp_desc_2_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_14_reg(uc2rb_rd_resp_desc_2_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_15_reg(uc2rb_rd_resp_desc_2_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_2_resp_reg(uc2rb_wr_resp_desc_2_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xid_0_reg(uc2rb_wr_resp_desc_2_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xid_1_reg(uc2rb_wr_resp_desc_2_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xid_2_reg(uc2rb_wr_resp_desc_2_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xid_3_reg(uc2rb_wr_resp_desc_2_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_0_reg(uc2rb_wr_resp_desc_2_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_1_reg(uc2rb_wr_resp_desc_2_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_2_reg(uc2rb_wr_resp_desc_2_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_3_reg(uc2rb_wr_resp_desc_2_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_4_reg(uc2rb_wr_resp_desc_2_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_5_reg(uc2rb_wr_resp_desc_2_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_6_reg(uc2rb_wr_resp_desc_2_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_7_reg(uc2rb_wr_resp_desc_2_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_8_reg(uc2rb_wr_resp_desc_2_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_9_reg(uc2rb_wr_resp_desc_2_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_10_reg(uc2rb_wr_resp_desc_2_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_11_reg(uc2rb_wr_resp_desc_2_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_12_reg(uc2rb_wr_resp_desc_2_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_13_reg(uc2rb_wr_resp_desc_2_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_14_reg(uc2rb_wr_resp_desc_2_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_15_reg(uc2rb_wr_resp_desc_2_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_2_attr_reg(uc2rb_sn_req_desc_2_attr_reg),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_0_reg(uc2rb_sn_req_desc_2_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_1_reg(uc2rb_sn_req_desc_2_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_2_reg(uc2rb_sn_req_desc_2_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_3_reg(uc2rb_sn_req_desc_2_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_3_data_offset_reg(uc2rb_rd_resp_desc_3_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_3_data_size_reg(uc2rb_rd_resp_desc_3_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_3_resp_reg(uc2rb_rd_resp_desc_3_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xid_0_reg(uc2rb_rd_resp_desc_3_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xid_1_reg(uc2rb_rd_resp_desc_3_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xid_2_reg(uc2rb_rd_resp_desc_3_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xid_3_reg(uc2rb_rd_resp_desc_3_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_0_reg(uc2rb_rd_resp_desc_3_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_1_reg(uc2rb_rd_resp_desc_3_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_2_reg(uc2rb_rd_resp_desc_3_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_3_reg(uc2rb_rd_resp_desc_3_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_4_reg(uc2rb_rd_resp_desc_3_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_5_reg(uc2rb_rd_resp_desc_3_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_6_reg(uc2rb_rd_resp_desc_3_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_7_reg(uc2rb_rd_resp_desc_3_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_8_reg(uc2rb_rd_resp_desc_3_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_9_reg(uc2rb_rd_resp_desc_3_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_10_reg(uc2rb_rd_resp_desc_3_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_11_reg(uc2rb_rd_resp_desc_3_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_12_reg(uc2rb_rd_resp_desc_3_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_13_reg(uc2rb_rd_resp_desc_3_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_14_reg(uc2rb_rd_resp_desc_3_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_15_reg(uc2rb_rd_resp_desc_3_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_3_resp_reg(uc2rb_wr_resp_desc_3_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xid_0_reg(uc2rb_wr_resp_desc_3_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xid_1_reg(uc2rb_wr_resp_desc_3_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xid_2_reg(uc2rb_wr_resp_desc_3_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xid_3_reg(uc2rb_wr_resp_desc_3_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_0_reg(uc2rb_wr_resp_desc_3_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_1_reg(uc2rb_wr_resp_desc_3_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_2_reg(uc2rb_wr_resp_desc_3_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_3_reg(uc2rb_wr_resp_desc_3_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_4_reg(uc2rb_wr_resp_desc_3_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_5_reg(uc2rb_wr_resp_desc_3_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_6_reg(uc2rb_wr_resp_desc_3_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_7_reg(uc2rb_wr_resp_desc_3_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_8_reg(uc2rb_wr_resp_desc_3_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_9_reg(uc2rb_wr_resp_desc_3_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_10_reg(uc2rb_wr_resp_desc_3_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_11_reg(uc2rb_wr_resp_desc_3_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_12_reg(uc2rb_wr_resp_desc_3_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_13_reg(uc2rb_wr_resp_desc_3_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_14_reg(uc2rb_wr_resp_desc_3_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_15_reg(uc2rb_wr_resp_desc_3_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_3_attr_reg(uc2rb_sn_req_desc_3_attr_reg),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_0_reg(uc2rb_sn_req_desc_3_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_1_reg(uc2rb_sn_req_desc_3_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_2_reg(uc2rb_sn_req_desc_3_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_3_reg(uc2rb_sn_req_desc_3_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_4_data_offset_reg(uc2rb_rd_resp_desc_4_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_4_data_size_reg(uc2rb_rd_resp_desc_4_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_4_resp_reg(uc2rb_rd_resp_desc_4_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xid_0_reg(uc2rb_rd_resp_desc_4_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xid_1_reg(uc2rb_rd_resp_desc_4_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xid_2_reg(uc2rb_rd_resp_desc_4_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xid_3_reg(uc2rb_rd_resp_desc_4_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_0_reg(uc2rb_rd_resp_desc_4_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_1_reg(uc2rb_rd_resp_desc_4_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_2_reg(uc2rb_rd_resp_desc_4_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_3_reg(uc2rb_rd_resp_desc_4_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_4_reg(uc2rb_rd_resp_desc_4_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_5_reg(uc2rb_rd_resp_desc_4_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_6_reg(uc2rb_rd_resp_desc_4_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_7_reg(uc2rb_rd_resp_desc_4_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_8_reg(uc2rb_rd_resp_desc_4_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_9_reg(uc2rb_rd_resp_desc_4_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_10_reg(uc2rb_rd_resp_desc_4_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_11_reg(uc2rb_rd_resp_desc_4_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_12_reg(uc2rb_rd_resp_desc_4_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_13_reg(uc2rb_rd_resp_desc_4_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_14_reg(uc2rb_rd_resp_desc_4_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_15_reg(uc2rb_rd_resp_desc_4_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_4_resp_reg(uc2rb_wr_resp_desc_4_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xid_0_reg(uc2rb_wr_resp_desc_4_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xid_1_reg(uc2rb_wr_resp_desc_4_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xid_2_reg(uc2rb_wr_resp_desc_4_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xid_3_reg(uc2rb_wr_resp_desc_4_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_0_reg(uc2rb_wr_resp_desc_4_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_1_reg(uc2rb_wr_resp_desc_4_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_2_reg(uc2rb_wr_resp_desc_4_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_3_reg(uc2rb_wr_resp_desc_4_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_4_reg(uc2rb_wr_resp_desc_4_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_5_reg(uc2rb_wr_resp_desc_4_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_6_reg(uc2rb_wr_resp_desc_4_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_7_reg(uc2rb_wr_resp_desc_4_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_8_reg(uc2rb_wr_resp_desc_4_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_9_reg(uc2rb_wr_resp_desc_4_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_10_reg(uc2rb_wr_resp_desc_4_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_11_reg(uc2rb_wr_resp_desc_4_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_12_reg(uc2rb_wr_resp_desc_4_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_13_reg(uc2rb_wr_resp_desc_4_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_14_reg(uc2rb_wr_resp_desc_4_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_15_reg(uc2rb_wr_resp_desc_4_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_4_attr_reg(uc2rb_sn_req_desc_4_attr_reg),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_0_reg(uc2rb_sn_req_desc_4_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_1_reg(uc2rb_sn_req_desc_4_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_2_reg(uc2rb_sn_req_desc_4_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_3_reg(uc2rb_sn_req_desc_4_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_5_data_offset_reg(uc2rb_rd_resp_desc_5_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_5_data_size_reg(uc2rb_rd_resp_desc_5_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_5_resp_reg(uc2rb_rd_resp_desc_5_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xid_0_reg(uc2rb_rd_resp_desc_5_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xid_1_reg(uc2rb_rd_resp_desc_5_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xid_2_reg(uc2rb_rd_resp_desc_5_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xid_3_reg(uc2rb_rd_resp_desc_5_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_0_reg(uc2rb_rd_resp_desc_5_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_1_reg(uc2rb_rd_resp_desc_5_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_2_reg(uc2rb_rd_resp_desc_5_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_3_reg(uc2rb_rd_resp_desc_5_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_4_reg(uc2rb_rd_resp_desc_5_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_5_reg(uc2rb_rd_resp_desc_5_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_6_reg(uc2rb_rd_resp_desc_5_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_7_reg(uc2rb_rd_resp_desc_5_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_8_reg(uc2rb_rd_resp_desc_5_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_9_reg(uc2rb_rd_resp_desc_5_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_10_reg(uc2rb_rd_resp_desc_5_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_11_reg(uc2rb_rd_resp_desc_5_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_12_reg(uc2rb_rd_resp_desc_5_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_13_reg(uc2rb_rd_resp_desc_5_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_14_reg(uc2rb_rd_resp_desc_5_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_15_reg(uc2rb_rd_resp_desc_5_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_5_resp_reg(uc2rb_wr_resp_desc_5_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xid_0_reg(uc2rb_wr_resp_desc_5_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xid_1_reg(uc2rb_wr_resp_desc_5_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xid_2_reg(uc2rb_wr_resp_desc_5_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xid_3_reg(uc2rb_wr_resp_desc_5_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_0_reg(uc2rb_wr_resp_desc_5_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_1_reg(uc2rb_wr_resp_desc_5_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_2_reg(uc2rb_wr_resp_desc_5_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_3_reg(uc2rb_wr_resp_desc_5_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_4_reg(uc2rb_wr_resp_desc_5_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_5_reg(uc2rb_wr_resp_desc_5_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_6_reg(uc2rb_wr_resp_desc_5_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_7_reg(uc2rb_wr_resp_desc_5_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_8_reg(uc2rb_wr_resp_desc_5_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_9_reg(uc2rb_wr_resp_desc_5_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_10_reg(uc2rb_wr_resp_desc_5_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_11_reg(uc2rb_wr_resp_desc_5_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_12_reg(uc2rb_wr_resp_desc_5_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_13_reg(uc2rb_wr_resp_desc_5_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_14_reg(uc2rb_wr_resp_desc_5_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_15_reg(uc2rb_wr_resp_desc_5_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_5_attr_reg(uc2rb_sn_req_desc_5_attr_reg),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_0_reg(uc2rb_sn_req_desc_5_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_1_reg(uc2rb_sn_req_desc_5_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_2_reg(uc2rb_sn_req_desc_5_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_3_reg(uc2rb_sn_req_desc_5_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_6_data_offset_reg(uc2rb_rd_resp_desc_6_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_6_data_size_reg(uc2rb_rd_resp_desc_6_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_6_resp_reg(uc2rb_rd_resp_desc_6_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xid_0_reg(uc2rb_rd_resp_desc_6_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xid_1_reg(uc2rb_rd_resp_desc_6_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xid_2_reg(uc2rb_rd_resp_desc_6_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xid_3_reg(uc2rb_rd_resp_desc_6_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_0_reg(uc2rb_rd_resp_desc_6_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_1_reg(uc2rb_rd_resp_desc_6_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_2_reg(uc2rb_rd_resp_desc_6_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_3_reg(uc2rb_rd_resp_desc_6_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_4_reg(uc2rb_rd_resp_desc_6_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_5_reg(uc2rb_rd_resp_desc_6_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_6_reg(uc2rb_rd_resp_desc_6_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_7_reg(uc2rb_rd_resp_desc_6_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_8_reg(uc2rb_rd_resp_desc_6_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_9_reg(uc2rb_rd_resp_desc_6_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_10_reg(uc2rb_rd_resp_desc_6_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_11_reg(uc2rb_rd_resp_desc_6_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_12_reg(uc2rb_rd_resp_desc_6_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_13_reg(uc2rb_rd_resp_desc_6_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_14_reg(uc2rb_rd_resp_desc_6_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_15_reg(uc2rb_rd_resp_desc_6_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_6_resp_reg(uc2rb_wr_resp_desc_6_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xid_0_reg(uc2rb_wr_resp_desc_6_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xid_1_reg(uc2rb_wr_resp_desc_6_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xid_2_reg(uc2rb_wr_resp_desc_6_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xid_3_reg(uc2rb_wr_resp_desc_6_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_0_reg(uc2rb_wr_resp_desc_6_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_1_reg(uc2rb_wr_resp_desc_6_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_2_reg(uc2rb_wr_resp_desc_6_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_3_reg(uc2rb_wr_resp_desc_6_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_4_reg(uc2rb_wr_resp_desc_6_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_5_reg(uc2rb_wr_resp_desc_6_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_6_reg(uc2rb_wr_resp_desc_6_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_7_reg(uc2rb_wr_resp_desc_6_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_8_reg(uc2rb_wr_resp_desc_6_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_9_reg(uc2rb_wr_resp_desc_6_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_10_reg(uc2rb_wr_resp_desc_6_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_11_reg(uc2rb_wr_resp_desc_6_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_12_reg(uc2rb_wr_resp_desc_6_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_13_reg(uc2rb_wr_resp_desc_6_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_14_reg(uc2rb_wr_resp_desc_6_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_15_reg(uc2rb_wr_resp_desc_6_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_6_attr_reg(uc2rb_sn_req_desc_6_attr_reg),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_0_reg(uc2rb_sn_req_desc_6_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_1_reg(uc2rb_sn_req_desc_6_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_2_reg(uc2rb_sn_req_desc_6_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_3_reg(uc2rb_sn_req_desc_6_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_7_data_offset_reg(uc2rb_rd_resp_desc_7_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_7_data_size_reg(uc2rb_rd_resp_desc_7_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_7_resp_reg(uc2rb_rd_resp_desc_7_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xid_0_reg(uc2rb_rd_resp_desc_7_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xid_1_reg(uc2rb_rd_resp_desc_7_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xid_2_reg(uc2rb_rd_resp_desc_7_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xid_3_reg(uc2rb_rd_resp_desc_7_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_0_reg(uc2rb_rd_resp_desc_7_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_1_reg(uc2rb_rd_resp_desc_7_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_2_reg(uc2rb_rd_resp_desc_7_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_3_reg(uc2rb_rd_resp_desc_7_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_4_reg(uc2rb_rd_resp_desc_7_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_5_reg(uc2rb_rd_resp_desc_7_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_6_reg(uc2rb_rd_resp_desc_7_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_7_reg(uc2rb_rd_resp_desc_7_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_8_reg(uc2rb_rd_resp_desc_7_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_9_reg(uc2rb_rd_resp_desc_7_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_10_reg(uc2rb_rd_resp_desc_7_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_11_reg(uc2rb_rd_resp_desc_7_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_12_reg(uc2rb_rd_resp_desc_7_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_13_reg(uc2rb_rd_resp_desc_7_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_14_reg(uc2rb_rd_resp_desc_7_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_15_reg(uc2rb_rd_resp_desc_7_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_7_resp_reg(uc2rb_wr_resp_desc_7_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xid_0_reg(uc2rb_wr_resp_desc_7_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xid_1_reg(uc2rb_wr_resp_desc_7_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xid_2_reg(uc2rb_wr_resp_desc_7_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xid_3_reg(uc2rb_wr_resp_desc_7_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_0_reg(uc2rb_wr_resp_desc_7_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_1_reg(uc2rb_wr_resp_desc_7_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_2_reg(uc2rb_wr_resp_desc_7_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_3_reg(uc2rb_wr_resp_desc_7_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_4_reg(uc2rb_wr_resp_desc_7_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_5_reg(uc2rb_wr_resp_desc_7_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_6_reg(uc2rb_wr_resp_desc_7_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_7_reg(uc2rb_wr_resp_desc_7_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_8_reg(uc2rb_wr_resp_desc_7_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_9_reg(uc2rb_wr_resp_desc_7_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_10_reg(uc2rb_wr_resp_desc_7_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_11_reg(uc2rb_wr_resp_desc_7_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_12_reg(uc2rb_wr_resp_desc_7_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_13_reg(uc2rb_wr_resp_desc_7_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_14_reg(uc2rb_wr_resp_desc_7_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_15_reg(uc2rb_wr_resp_desc_7_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_7_attr_reg(uc2rb_sn_req_desc_7_attr_reg),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_0_reg(uc2rb_sn_req_desc_7_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_1_reg(uc2rb_sn_req_desc_7_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_2_reg(uc2rb_sn_req_desc_7_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_3_reg(uc2rb_sn_req_desc_7_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_8_data_offset_reg(uc2rb_rd_resp_desc_8_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_8_data_size_reg(uc2rb_rd_resp_desc_8_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_8_resp_reg(uc2rb_rd_resp_desc_8_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xid_0_reg(uc2rb_rd_resp_desc_8_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xid_1_reg(uc2rb_rd_resp_desc_8_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xid_2_reg(uc2rb_rd_resp_desc_8_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xid_3_reg(uc2rb_rd_resp_desc_8_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_0_reg(uc2rb_rd_resp_desc_8_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_1_reg(uc2rb_rd_resp_desc_8_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_2_reg(uc2rb_rd_resp_desc_8_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_3_reg(uc2rb_rd_resp_desc_8_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_4_reg(uc2rb_rd_resp_desc_8_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_5_reg(uc2rb_rd_resp_desc_8_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_6_reg(uc2rb_rd_resp_desc_8_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_7_reg(uc2rb_rd_resp_desc_8_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_8_reg(uc2rb_rd_resp_desc_8_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_9_reg(uc2rb_rd_resp_desc_8_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_10_reg(uc2rb_rd_resp_desc_8_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_11_reg(uc2rb_rd_resp_desc_8_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_12_reg(uc2rb_rd_resp_desc_8_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_13_reg(uc2rb_rd_resp_desc_8_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_14_reg(uc2rb_rd_resp_desc_8_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_15_reg(uc2rb_rd_resp_desc_8_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_8_resp_reg(uc2rb_wr_resp_desc_8_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xid_0_reg(uc2rb_wr_resp_desc_8_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xid_1_reg(uc2rb_wr_resp_desc_8_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xid_2_reg(uc2rb_wr_resp_desc_8_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xid_3_reg(uc2rb_wr_resp_desc_8_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_0_reg(uc2rb_wr_resp_desc_8_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_1_reg(uc2rb_wr_resp_desc_8_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_2_reg(uc2rb_wr_resp_desc_8_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_3_reg(uc2rb_wr_resp_desc_8_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_4_reg(uc2rb_wr_resp_desc_8_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_5_reg(uc2rb_wr_resp_desc_8_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_6_reg(uc2rb_wr_resp_desc_8_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_7_reg(uc2rb_wr_resp_desc_8_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_8_reg(uc2rb_wr_resp_desc_8_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_9_reg(uc2rb_wr_resp_desc_8_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_10_reg(uc2rb_wr_resp_desc_8_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_11_reg(uc2rb_wr_resp_desc_8_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_12_reg(uc2rb_wr_resp_desc_8_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_13_reg(uc2rb_wr_resp_desc_8_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_14_reg(uc2rb_wr_resp_desc_8_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_15_reg(uc2rb_wr_resp_desc_8_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_8_attr_reg(uc2rb_sn_req_desc_8_attr_reg),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_0_reg(uc2rb_sn_req_desc_8_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_1_reg(uc2rb_sn_req_desc_8_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_2_reg(uc2rb_sn_req_desc_8_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_3_reg(uc2rb_sn_req_desc_8_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_9_data_offset_reg(uc2rb_rd_resp_desc_9_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_9_data_size_reg(uc2rb_rd_resp_desc_9_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_9_resp_reg(uc2rb_rd_resp_desc_9_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xid_0_reg(uc2rb_rd_resp_desc_9_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xid_1_reg(uc2rb_rd_resp_desc_9_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xid_2_reg(uc2rb_rd_resp_desc_9_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xid_3_reg(uc2rb_rd_resp_desc_9_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_0_reg(uc2rb_rd_resp_desc_9_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_1_reg(uc2rb_rd_resp_desc_9_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_2_reg(uc2rb_rd_resp_desc_9_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_3_reg(uc2rb_rd_resp_desc_9_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_4_reg(uc2rb_rd_resp_desc_9_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_5_reg(uc2rb_rd_resp_desc_9_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_6_reg(uc2rb_rd_resp_desc_9_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_7_reg(uc2rb_rd_resp_desc_9_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_8_reg(uc2rb_rd_resp_desc_9_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_9_reg(uc2rb_rd_resp_desc_9_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_10_reg(uc2rb_rd_resp_desc_9_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_11_reg(uc2rb_rd_resp_desc_9_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_12_reg(uc2rb_rd_resp_desc_9_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_13_reg(uc2rb_rd_resp_desc_9_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_14_reg(uc2rb_rd_resp_desc_9_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_15_reg(uc2rb_rd_resp_desc_9_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_9_resp_reg(uc2rb_wr_resp_desc_9_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xid_0_reg(uc2rb_wr_resp_desc_9_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xid_1_reg(uc2rb_wr_resp_desc_9_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xid_2_reg(uc2rb_wr_resp_desc_9_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xid_3_reg(uc2rb_wr_resp_desc_9_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_0_reg(uc2rb_wr_resp_desc_9_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_1_reg(uc2rb_wr_resp_desc_9_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_2_reg(uc2rb_wr_resp_desc_9_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_3_reg(uc2rb_wr_resp_desc_9_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_4_reg(uc2rb_wr_resp_desc_9_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_5_reg(uc2rb_wr_resp_desc_9_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_6_reg(uc2rb_wr_resp_desc_9_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_7_reg(uc2rb_wr_resp_desc_9_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_8_reg(uc2rb_wr_resp_desc_9_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_9_reg(uc2rb_wr_resp_desc_9_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_10_reg(uc2rb_wr_resp_desc_9_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_11_reg(uc2rb_wr_resp_desc_9_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_12_reg(uc2rb_wr_resp_desc_9_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_13_reg(uc2rb_wr_resp_desc_9_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_14_reg(uc2rb_wr_resp_desc_9_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_15_reg(uc2rb_wr_resp_desc_9_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_9_attr_reg(uc2rb_sn_req_desc_9_attr_reg),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_0_reg(uc2rb_sn_req_desc_9_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_1_reg(uc2rb_sn_req_desc_9_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_2_reg(uc2rb_sn_req_desc_9_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_3_reg(uc2rb_sn_req_desc_9_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_a_data_offset_reg(uc2rb_rd_resp_desc_a_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_a_data_size_reg(uc2rb_rd_resp_desc_a_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_a_resp_reg(uc2rb_rd_resp_desc_a_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xid_0_reg(uc2rb_rd_resp_desc_a_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xid_1_reg(uc2rb_rd_resp_desc_a_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xid_2_reg(uc2rb_rd_resp_desc_a_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xid_3_reg(uc2rb_rd_resp_desc_a_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_0_reg(uc2rb_rd_resp_desc_a_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_1_reg(uc2rb_rd_resp_desc_a_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_2_reg(uc2rb_rd_resp_desc_a_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_3_reg(uc2rb_rd_resp_desc_a_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_4_reg(uc2rb_rd_resp_desc_a_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_5_reg(uc2rb_rd_resp_desc_a_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_6_reg(uc2rb_rd_resp_desc_a_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_7_reg(uc2rb_rd_resp_desc_a_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_8_reg(uc2rb_rd_resp_desc_a_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_9_reg(uc2rb_rd_resp_desc_a_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_10_reg(uc2rb_rd_resp_desc_a_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_11_reg(uc2rb_rd_resp_desc_a_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_12_reg(uc2rb_rd_resp_desc_a_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_13_reg(uc2rb_rd_resp_desc_a_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_14_reg(uc2rb_rd_resp_desc_a_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_15_reg(uc2rb_rd_resp_desc_a_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_a_resp_reg(uc2rb_wr_resp_desc_a_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xid_0_reg(uc2rb_wr_resp_desc_a_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xid_1_reg(uc2rb_wr_resp_desc_a_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xid_2_reg(uc2rb_wr_resp_desc_a_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xid_3_reg(uc2rb_wr_resp_desc_a_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_0_reg(uc2rb_wr_resp_desc_a_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_1_reg(uc2rb_wr_resp_desc_a_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_2_reg(uc2rb_wr_resp_desc_a_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_3_reg(uc2rb_wr_resp_desc_a_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_4_reg(uc2rb_wr_resp_desc_a_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_5_reg(uc2rb_wr_resp_desc_a_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_6_reg(uc2rb_wr_resp_desc_a_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_7_reg(uc2rb_wr_resp_desc_a_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_8_reg(uc2rb_wr_resp_desc_a_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_9_reg(uc2rb_wr_resp_desc_a_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_10_reg(uc2rb_wr_resp_desc_a_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_11_reg(uc2rb_wr_resp_desc_a_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_12_reg(uc2rb_wr_resp_desc_a_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_13_reg(uc2rb_wr_resp_desc_a_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_14_reg(uc2rb_wr_resp_desc_a_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_15_reg(uc2rb_wr_resp_desc_a_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_a_attr_reg(uc2rb_sn_req_desc_a_attr_reg),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_0_reg(uc2rb_sn_req_desc_a_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_1_reg(uc2rb_sn_req_desc_a_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_2_reg(uc2rb_sn_req_desc_a_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_3_reg(uc2rb_sn_req_desc_a_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_b_data_offset_reg(uc2rb_rd_resp_desc_b_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_b_data_size_reg(uc2rb_rd_resp_desc_b_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_b_resp_reg(uc2rb_rd_resp_desc_b_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xid_0_reg(uc2rb_rd_resp_desc_b_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xid_1_reg(uc2rb_rd_resp_desc_b_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xid_2_reg(uc2rb_rd_resp_desc_b_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xid_3_reg(uc2rb_rd_resp_desc_b_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_0_reg(uc2rb_rd_resp_desc_b_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_1_reg(uc2rb_rd_resp_desc_b_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_2_reg(uc2rb_rd_resp_desc_b_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_3_reg(uc2rb_rd_resp_desc_b_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_4_reg(uc2rb_rd_resp_desc_b_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_5_reg(uc2rb_rd_resp_desc_b_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_6_reg(uc2rb_rd_resp_desc_b_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_7_reg(uc2rb_rd_resp_desc_b_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_8_reg(uc2rb_rd_resp_desc_b_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_9_reg(uc2rb_rd_resp_desc_b_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_10_reg(uc2rb_rd_resp_desc_b_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_11_reg(uc2rb_rd_resp_desc_b_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_12_reg(uc2rb_rd_resp_desc_b_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_13_reg(uc2rb_rd_resp_desc_b_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_14_reg(uc2rb_rd_resp_desc_b_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_15_reg(uc2rb_rd_resp_desc_b_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_b_resp_reg(uc2rb_wr_resp_desc_b_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xid_0_reg(uc2rb_wr_resp_desc_b_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xid_1_reg(uc2rb_wr_resp_desc_b_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xid_2_reg(uc2rb_wr_resp_desc_b_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xid_3_reg(uc2rb_wr_resp_desc_b_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_0_reg(uc2rb_wr_resp_desc_b_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_1_reg(uc2rb_wr_resp_desc_b_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_2_reg(uc2rb_wr_resp_desc_b_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_3_reg(uc2rb_wr_resp_desc_b_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_4_reg(uc2rb_wr_resp_desc_b_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_5_reg(uc2rb_wr_resp_desc_b_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_6_reg(uc2rb_wr_resp_desc_b_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_7_reg(uc2rb_wr_resp_desc_b_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_8_reg(uc2rb_wr_resp_desc_b_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_9_reg(uc2rb_wr_resp_desc_b_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_10_reg(uc2rb_wr_resp_desc_b_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_11_reg(uc2rb_wr_resp_desc_b_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_12_reg(uc2rb_wr_resp_desc_b_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_13_reg(uc2rb_wr_resp_desc_b_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_14_reg(uc2rb_wr_resp_desc_b_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_15_reg(uc2rb_wr_resp_desc_b_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_b_attr_reg(uc2rb_sn_req_desc_b_attr_reg),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_0_reg(uc2rb_sn_req_desc_b_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_1_reg(uc2rb_sn_req_desc_b_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_2_reg(uc2rb_sn_req_desc_b_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_3_reg(uc2rb_sn_req_desc_b_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_c_data_offset_reg(uc2rb_rd_resp_desc_c_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_c_data_size_reg(uc2rb_rd_resp_desc_c_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_c_resp_reg(uc2rb_rd_resp_desc_c_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xid_0_reg(uc2rb_rd_resp_desc_c_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xid_1_reg(uc2rb_rd_resp_desc_c_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xid_2_reg(uc2rb_rd_resp_desc_c_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xid_3_reg(uc2rb_rd_resp_desc_c_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_0_reg(uc2rb_rd_resp_desc_c_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_1_reg(uc2rb_rd_resp_desc_c_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_2_reg(uc2rb_rd_resp_desc_c_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_3_reg(uc2rb_rd_resp_desc_c_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_4_reg(uc2rb_rd_resp_desc_c_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_5_reg(uc2rb_rd_resp_desc_c_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_6_reg(uc2rb_rd_resp_desc_c_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_7_reg(uc2rb_rd_resp_desc_c_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_8_reg(uc2rb_rd_resp_desc_c_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_9_reg(uc2rb_rd_resp_desc_c_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_10_reg(uc2rb_rd_resp_desc_c_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_11_reg(uc2rb_rd_resp_desc_c_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_12_reg(uc2rb_rd_resp_desc_c_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_13_reg(uc2rb_rd_resp_desc_c_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_14_reg(uc2rb_rd_resp_desc_c_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_15_reg(uc2rb_rd_resp_desc_c_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_c_resp_reg(uc2rb_wr_resp_desc_c_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xid_0_reg(uc2rb_wr_resp_desc_c_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xid_1_reg(uc2rb_wr_resp_desc_c_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xid_2_reg(uc2rb_wr_resp_desc_c_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xid_3_reg(uc2rb_wr_resp_desc_c_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_0_reg(uc2rb_wr_resp_desc_c_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_1_reg(uc2rb_wr_resp_desc_c_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_2_reg(uc2rb_wr_resp_desc_c_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_3_reg(uc2rb_wr_resp_desc_c_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_4_reg(uc2rb_wr_resp_desc_c_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_5_reg(uc2rb_wr_resp_desc_c_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_6_reg(uc2rb_wr_resp_desc_c_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_7_reg(uc2rb_wr_resp_desc_c_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_8_reg(uc2rb_wr_resp_desc_c_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_9_reg(uc2rb_wr_resp_desc_c_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_10_reg(uc2rb_wr_resp_desc_c_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_11_reg(uc2rb_wr_resp_desc_c_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_12_reg(uc2rb_wr_resp_desc_c_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_13_reg(uc2rb_wr_resp_desc_c_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_14_reg(uc2rb_wr_resp_desc_c_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_15_reg(uc2rb_wr_resp_desc_c_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_c_attr_reg(uc2rb_sn_req_desc_c_attr_reg),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_0_reg(uc2rb_sn_req_desc_c_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_1_reg(uc2rb_sn_req_desc_c_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_2_reg(uc2rb_sn_req_desc_c_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_3_reg(uc2rb_sn_req_desc_c_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_d_data_offset_reg(uc2rb_rd_resp_desc_d_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_d_data_size_reg(uc2rb_rd_resp_desc_d_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_d_resp_reg(uc2rb_rd_resp_desc_d_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xid_0_reg(uc2rb_rd_resp_desc_d_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xid_1_reg(uc2rb_rd_resp_desc_d_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xid_2_reg(uc2rb_rd_resp_desc_d_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xid_3_reg(uc2rb_rd_resp_desc_d_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_0_reg(uc2rb_rd_resp_desc_d_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_1_reg(uc2rb_rd_resp_desc_d_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_2_reg(uc2rb_rd_resp_desc_d_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_3_reg(uc2rb_rd_resp_desc_d_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_4_reg(uc2rb_rd_resp_desc_d_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_5_reg(uc2rb_rd_resp_desc_d_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_6_reg(uc2rb_rd_resp_desc_d_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_7_reg(uc2rb_rd_resp_desc_d_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_8_reg(uc2rb_rd_resp_desc_d_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_9_reg(uc2rb_rd_resp_desc_d_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_10_reg(uc2rb_rd_resp_desc_d_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_11_reg(uc2rb_rd_resp_desc_d_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_12_reg(uc2rb_rd_resp_desc_d_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_13_reg(uc2rb_rd_resp_desc_d_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_14_reg(uc2rb_rd_resp_desc_d_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_15_reg(uc2rb_rd_resp_desc_d_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_d_resp_reg(uc2rb_wr_resp_desc_d_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xid_0_reg(uc2rb_wr_resp_desc_d_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xid_1_reg(uc2rb_wr_resp_desc_d_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xid_2_reg(uc2rb_wr_resp_desc_d_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xid_3_reg(uc2rb_wr_resp_desc_d_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_0_reg(uc2rb_wr_resp_desc_d_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_1_reg(uc2rb_wr_resp_desc_d_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_2_reg(uc2rb_wr_resp_desc_d_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_3_reg(uc2rb_wr_resp_desc_d_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_4_reg(uc2rb_wr_resp_desc_d_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_5_reg(uc2rb_wr_resp_desc_d_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_6_reg(uc2rb_wr_resp_desc_d_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_7_reg(uc2rb_wr_resp_desc_d_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_8_reg(uc2rb_wr_resp_desc_d_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_9_reg(uc2rb_wr_resp_desc_d_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_10_reg(uc2rb_wr_resp_desc_d_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_11_reg(uc2rb_wr_resp_desc_d_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_12_reg(uc2rb_wr_resp_desc_d_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_13_reg(uc2rb_wr_resp_desc_d_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_14_reg(uc2rb_wr_resp_desc_d_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_15_reg(uc2rb_wr_resp_desc_d_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_d_attr_reg(uc2rb_sn_req_desc_d_attr_reg),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_0_reg(uc2rb_sn_req_desc_d_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_1_reg(uc2rb_sn_req_desc_d_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_2_reg(uc2rb_sn_req_desc_d_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_3_reg(uc2rb_sn_req_desc_d_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_e_data_offset_reg(uc2rb_rd_resp_desc_e_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_e_data_size_reg(uc2rb_rd_resp_desc_e_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_e_resp_reg(uc2rb_rd_resp_desc_e_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xid_0_reg(uc2rb_rd_resp_desc_e_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xid_1_reg(uc2rb_rd_resp_desc_e_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xid_2_reg(uc2rb_rd_resp_desc_e_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xid_3_reg(uc2rb_rd_resp_desc_e_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_0_reg(uc2rb_rd_resp_desc_e_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_1_reg(uc2rb_rd_resp_desc_e_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_2_reg(uc2rb_rd_resp_desc_e_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_3_reg(uc2rb_rd_resp_desc_e_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_4_reg(uc2rb_rd_resp_desc_e_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_5_reg(uc2rb_rd_resp_desc_e_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_6_reg(uc2rb_rd_resp_desc_e_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_7_reg(uc2rb_rd_resp_desc_e_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_8_reg(uc2rb_rd_resp_desc_e_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_9_reg(uc2rb_rd_resp_desc_e_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_10_reg(uc2rb_rd_resp_desc_e_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_11_reg(uc2rb_rd_resp_desc_e_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_12_reg(uc2rb_rd_resp_desc_e_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_13_reg(uc2rb_rd_resp_desc_e_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_14_reg(uc2rb_rd_resp_desc_e_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_15_reg(uc2rb_rd_resp_desc_e_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_e_resp_reg(uc2rb_wr_resp_desc_e_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xid_0_reg(uc2rb_wr_resp_desc_e_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xid_1_reg(uc2rb_wr_resp_desc_e_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xid_2_reg(uc2rb_wr_resp_desc_e_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xid_3_reg(uc2rb_wr_resp_desc_e_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_0_reg(uc2rb_wr_resp_desc_e_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_1_reg(uc2rb_wr_resp_desc_e_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_2_reg(uc2rb_wr_resp_desc_e_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_3_reg(uc2rb_wr_resp_desc_e_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_4_reg(uc2rb_wr_resp_desc_e_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_5_reg(uc2rb_wr_resp_desc_e_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_6_reg(uc2rb_wr_resp_desc_e_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_7_reg(uc2rb_wr_resp_desc_e_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_8_reg(uc2rb_wr_resp_desc_e_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_9_reg(uc2rb_wr_resp_desc_e_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_10_reg(uc2rb_wr_resp_desc_e_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_11_reg(uc2rb_wr_resp_desc_e_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_12_reg(uc2rb_wr_resp_desc_e_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_13_reg(uc2rb_wr_resp_desc_e_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_14_reg(uc2rb_wr_resp_desc_e_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_15_reg(uc2rb_wr_resp_desc_e_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_e_attr_reg(uc2rb_sn_req_desc_e_attr_reg),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_0_reg(uc2rb_sn_req_desc_e_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_1_reg(uc2rb_sn_req_desc_e_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_2_reg(uc2rb_sn_req_desc_e_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_3_reg(uc2rb_sn_req_desc_e_acaddr_3_reg),
                                                                                               .uc2rb_rd_resp_desc_f_data_offset_reg(uc2rb_rd_resp_desc_f_data_offset_reg),
                                                                                               .uc2rb_rd_resp_desc_f_data_size_reg(uc2rb_rd_resp_desc_f_data_size_reg),
                                                                                               .uc2rb_rd_resp_desc_f_resp_reg(uc2rb_rd_resp_desc_f_resp_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xid_0_reg(uc2rb_rd_resp_desc_f_xid_0_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xid_1_reg(uc2rb_rd_resp_desc_f_xid_1_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xid_2_reg(uc2rb_rd_resp_desc_f_xid_2_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xid_3_reg(uc2rb_rd_resp_desc_f_xid_3_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_0_reg(uc2rb_rd_resp_desc_f_xuser_0_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_1_reg(uc2rb_rd_resp_desc_f_xuser_1_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_2_reg(uc2rb_rd_resp_desc_f_xuser_2_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_3_reg(uc2rb_rd_resp_desc_f_xuser_3_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_4_reg(uc2rb_rd_resp_desc_f_xuser_4_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_5_reg(uc2rb_rd_resp_desc_f_xuser_5_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_6_reg(uc2rb_rd_resp_desc_f_xuser_6_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_7_reg(uc2rb_rd_resp_desc_f_xuser_7_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_8_reg(uc2rb_rd_resp_desc_f_xuser_8_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_9_reg(uc2rb_rd_resp_desc_f_xuser_9_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_10_reg(uc2rb_rd_resp_desc_f_xuser_10_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_11_reg(uc2rb_rd_resp_desc_f_xuser_11_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_12_reg(uc2rb_rd_resp_desc_f_xuser_12_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_13_reg(uc2rb_rd_resp_desc_f_xuser_13_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_14_reg(uc2rb_rd_resp_desc_f_xuser_14_reg),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_15_reg(uc2rb_rd_resp_desc_f_xuser_15_reg),
                                                                                               .uc2rb_wr_resp_desc_f_resp_reg(uc2rb_wr_resp_desc_f_resp_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xid_0_reg(uc2rb_wr_resp_desc_f_xid_0_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xid_1_reg(uc2rb_wr_resp_desc_f_xid_1_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xid_2_reg(uc2rb_wr_resp_desc_f_xid_2_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xid_3_reg(uc2rb_wr_resp_desc_f_xid_3_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_0_reg(uc2rb_wr_resp_desc_f_xuser_0_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_1_reg(uc2rb_wr_resp_desc_f_xuser_1_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_2_reg(uc2rb_wr_resp_desc_f_xuser_2_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_3_reg(uc2rb_wr_resp_desc_f_xuser_3_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_4_reg(uc2rb_wr_resp_desc_f_xuser_4_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_5_reg(uc2rb_wr_resp_desc_f_xuser_5_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_6_reg(uc2rb_wr_resp_desc_f_xuser_6_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_7_reg(uc2rb_wr_resp_desc_f_xuser_7_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_8_reg(uc2rb_wr_resp_desc_f_xuser_8_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_9_reg(uc2rb_wr_resp_desc_f_xuser_9_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_10_reg(uc2rb_wr_resp_desc_f_xuser_10_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_11_reg(uc2rb_wr_resp_desc_f_xuser_11_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_12_reg(uc2rb_wr_resp_desc_f_xuser_12_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_13_reg(uc2rb_wr_resp_desc_f_xuser_13_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_14_reg(uc2rb_wr_resp_desc_f_xuser_14_reg),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_15_reg(uc2rb_wr_resp_desc_f_xuser_15_reg),
                                                                                               .uc2rb_sn_req_desc_f_attr_reg(uc2rb_sn_req_desc_f_attr_reg),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_0_reg(uc2rb_sn_req_desc_f_acaddr_0_reg),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_1_reg(uc2rb_sn_req_desc_f_acaddr_1_reg),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_2_reg(uc2rb_sn_req_desc_f_acaddr_2_reg),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_3_reg(uc2rb_sn_req_desc_f_acaddr_3_reg),
                                                                                               .uc2rb_intr_error_status_reg_we(uc2rb_intr_error_status_reg_we),
                                                                                               .uc2rb_rd_req_fifo_free_level_reg_we(uc2rb_rd_req_fifo_free_level_reg_we),
                                                                                               .uc2rb_rd_req_intr_comp_status_reg_we(uc2rb_rd_req_intr_comp_status_reg_we),
                                                                                               .uc2rb_rd_resp_fifo_pop_desc_reg_we(uc2rb_rd_resp_fifo_pop_desc_reg_we),
                                                                                               .uc2rb_rd_resp_fifo_fill_level_reg_we(uc2rb_rd_resp_fifo_fill_level_reg_we),
                                                                                               .uc2rb_wr_req_fifo_free_level_reg_we(uc2rb_wr_req_fifo_free_level_reg_we),
                                                                                               .uc2rb_wr_req_intr_comp_status_reg_we(uc2rb_wr_req_intr_comp_status_reg_we),
                                                                                               .uc2rb_wr_resp_fifo_pop_desc_reg_we(uc2rb_wr_resp_fifo_pop_desc_reg_we),
                                                                                               .uc2rb_wr_resp_fifo_fill_level_reg_we(uc2rb_wr_resp_fifo_fill_level_reg_we),
                                                                                               .uc2rb_sn_req_fifo_pop_desc_reg_we(uc2rb_sn_req_fifo_pop_desc_reg_we),
                                                                                               .uc2rb_sn_req_fifo_fill_level_reg_we(uc2rb_sn_req_fifo_fill_level_reg_we),
                                                                                               .uc2rb_sn_resp_fifo_free_level_reg_we(uc2rb_sn_resp_fifo_free_level_reg_we),
                                                                                               .uc2rb_sn_resp_intr_comp_status_reg_we(uc2rb_sn_resp_intr_comp_status_reg_we),
                                                                                               .uc2rb_sn_data_fifo_free_level_reg_we(uc2rb_sn_data_fifo_free_level_reg_we),
                                                                                               .uc2rb_sn_data_intr_comp_status_reg_we(uc2rb_sn_data_intr_comp_status_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_data_offset_reg_we(uc2rb_rd_resp_desc_0_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_data_size_reg_we(uc2rb_rd_resp_desc_0_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_resp_reg_we(uc2rb_rd_resp_desc_0_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xid_0_reg_we(uc2rb_rd_resp_desc_0_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xid_1_reg_we(uc2rb_rd_resp_desc_0_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xid_2_reg_we(uc2rb_rd_resp_desc_0_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xid_3_reg_we(uc2rb_rd_resp_desc_0_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_0_reg_we(uc2rb_rd_resp_desc_0_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_1_reg_we(uc2rb_rd_resp_desc_0_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_2_reg_we(uc2rb_rd_resp_desc_0_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_3_reg_we(uc2rb_rd_resp_desc_0_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_4_reg_we(uc2rb_rd_resp_desc_0_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_5_reg_we(uc2rb_rd_resp_desc_0_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_6_reg_we(uc2rb_rd_resp_desc_0_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_7_reg_we(uc2rb_rd_resp_desc_0_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_8_reg_we(uc2rb_rd_resp_desc_0_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_9_reg_we(uc2rb_rd_resp_desc_0_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_10_reg_we(uc2rb_rd_resp_desc_0_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_11_reg_we(uc2rb_rd_resp_desc_0_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_12_reg_we(uc2rb_rd_resp_desc_0_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_13_reg_we(uc2rb_rd_resp_desc_0_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_14_reg_we(uc2rb_rd_resp_desc_0_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_0_xuser_15_reg_we(uc2rb_rd_resp_desc_0_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_resp_reg_we(uc2rb_wr_resp_desc_0_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xid_0_reg_we(uc2rb_wr_resp_desc_0_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xid_1_reg_we(uc2rb_wr_resp_desc_0_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xid_2_reg_we(uc2rb_wr_resp_desc_0_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xid_3_reg_we(uc2rb_wr_resp_desc_0_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_0_reg_we(uc2rb_wr_resp_desc_0_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_1_reg_we(uc2rb_wr_resp_desc_0_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_2_reg_we(uc2rb_wr_resp_desc_0_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_3_reg_we(uc2rb_wr_resp_desc_0_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_4_reg_we(uc2rb_wr_resp_desc_0_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_5_reg_we(uc2rb_wr_resp_desc_0_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_6_reg_we(uc2rb_wr_resp_desc_0_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_7_reg_we(uc2rb_wr_resp_desc_0_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_8_reg_we(uc2rb_wr_resp_desc_0_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_9_reg_we(uc2rb_wr_resp_desc_0_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_10_reg_we(uc2rb_wr_resp_desc_0_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_11_reg_we(uc2rb_wr_resp_desc_0_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_12_reg_we(uc2rb_wr_resp_desc_0_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_13_reg_we(uc2rb_wr_resp_desc_0_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_14_reg_we(uc2rb_wr_resp_desc_0_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_0_xuser_15_reg_we(uc2rb_wr_resp_desc_0_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_0_attr_reg_we(uc2rb_sn_req_desc_0_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_0_reg_we(uc2rb_sn_req_desc_0_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_1_reg_we(uc2rb_sn_req_desc_0_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_2_reg_we(uc2rb_sn_req_desc_0_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_0_acaddr_3_reg_we(uc2rb_sn_req_desc_0_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_data_offset_reg_we(uc2rb_rd_resp_desc_1_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_data_size_reg_we(uc2rb_rd_resp_desc_1_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_resp_reg_we(uc2rb_rd_resp_desc_1_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xid_0_reg_we(uc2rb_rd_resp_desc_1_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xid_1_reg_we(uc2rb_rd_resp_desc_1_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xid_2_reg_we(uc2rb_rd_resp_desc_1_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xid_3_reg_we(uc2rb_rd_resp_desc_1_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_0_reg_we(uc2rb_rd_resp_desc_1_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_1_reg_we(uc2rb_rd_resp_desc_1_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_2_reg_we(uc2rb_rd_resp_desc_1_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_3_reg_we(uc2rb_rd_resp_desc_1_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_4_reg_we(uc2rb_rd_resp_desc_1_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_5_reg_we(uc2rb_rd_resp_desc_1_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_6_reg_we(uc2rb_rd_resp_desc_1_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_7_reg_we(uc2rb_rd_resp_desc_1_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_8_reg_we(uc2rb_rd_resp_desc_1_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_9_reg_we(uc2rb_rd_resp_desc_1_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_10_reg_we(uc2rb_rd_resp_desc_1_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_11_reg_we(uc2rb_rd_resp_desc_1_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_12_reg_we(uc2rb_rd_resp_desc_1_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_13_reg_we(uc2rb_rd_resp_desc_1_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_14_reg_we(uc2rb_rd_resp_desc_1_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_1_xuser_15_reg_we(uc2rb_rd_resp_desc_1_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_resp_reg_we(uc2rb_wr_resp_desc_1_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xid_0_reg_we(uc2rb_wr_resp_desc_1_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xid_1_reg_we(uc2rb_wr_resp_desc_1_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xid_2_reg_we(uc2rb_wr_resp_desc_1_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xid_3_reg_we(uc2rb_wr_resp_desc_1_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_0_reg_we(uc2rb_wr_resp_desc_1_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_1_reg_we(uc2rb_wr_resp_desc_1_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_2_reg_we(uc2rb_wr_resp_desc_1_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_3_reg_we(uc2rb_wr_resp_desc_1_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_4_reg_we(uc2rb_wr_resp_desc_1_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_5_reg_we(uc2rb_wr_resp_desc_1_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_6_reg_we(uc2rb_wr_resp_desc_1_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_7_reg_we(uc2rb_wr_resp_desc_1_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_8_reg_we(uc2rb_wr_resp_desc_1_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_9_reg_we(uc2rb_wr_resp_desc_1_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_10_reg_we(uc2rb_wr_resp_desc_1_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_11_reg_we(uc2rb_wr_resp_desc_1_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_12_reg_we(uc2rb_wr_resp_desc_1_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_13_reg_we(uc2rb_wr_resp_desc_1_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_14_reg_we(uc2rb_wr_resp_desc_1_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_1_xuser_15_reg_we(uc2rb_wr_resp_desc_1_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_1_attr_reg_we(uc2rb_sn_req_desc_1_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_0_reg_we(uc2rb_sn_req_desc_1_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_1_reg_we(uc2rb_sn_req_desc_1_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_2_reg_we(uc2rb_sn_req_desc_1_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_1_acaddr_3_reg_we(uc2rb_sn_req_desc_1_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_data_offset_reg_we(uc2rb_rd_resp_desc_2_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_data_size_reg_we(uc2rb_rd_resp_desc_2_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_resp_reg_we(uc2rb_rd_resp_desc_2_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xid_0_reg_we(uc2rb_rd_resp_desc_2_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xid_1_reg_we(uc2rb_rd_resp_desc_2_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xid_2_reg_we(uc2rb_rd_resp_desc_2_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xid_3_reg_we(uc2rb_rd_resp_desc_2_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_0_reg_we(uc2rb_rd_resp_desc_2_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_1_reg_we(uc2rb_rd_resp_desc_2_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_2_reg_we(uc2rb_rd_resp_desc_2_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_3_reg_we(uc2rb_rd_resp_desc_2_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_4_reg_we(uc2rb_rd_resp_desc_2_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_5_reg_we(uc2rb_rd_resp_desc_2_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_6_reg_we(uc2rb_rd_resp_desc_2_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_7_reg_we(uc2rb_rd_resp_desc_2_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_8_reg_we(uc2rb_rd_resp_desc_2_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_9_reg_we(uc2rb_rd_resp_desc_2_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_10_reg_we(uc2rb_rd_resp_desc_2_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_11_reg_we(uc2rb_rd_resp_desc_2_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_12_reg_we(uc2rb_rd_resp_desc_2_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_13_reg_we(uc2rb_rd_resp_desc_2_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_14_reg_we(uc2rb_rd_resp_desc_2_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_2_xuser_15_reg_we(uc2rb_rd_resp_desc_2_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_resp_reg_we(uc2rb_wr_resp_desc_2_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xid_0_reg_we(uc2rb_wr_resp_desc_2_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xid_1_reg_we(uc2rb_wr_resp_desc_2_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xid_2_reg_we(uc2rb_wr_resp_desc_2_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xid_3_reg_we(uc2rb_wr_resp_desc_2_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_0_reg_we(uc2rb_wr_resp_desc_2_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_1_reg_we(uc2rb_wr_resp_desc_2_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_2_reg_we(uc2rb_wr_resp_desc_2_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_3_reg_we(uc2rb_wr_resp_desc_2_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_4_reg_we(uc2rb_wr_resp_desc_2_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_5_reg_we(uc2rb_wr_resp_desc_2_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_6_reg_we(uc2rb_wr_resp_desc_2_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_7_reg_we(uc2rb_wr_resp_desc_2_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_8_reg_we(uc2rb_wr_resp_desc_2_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_9_reg_we(uc2rb_wr_resp_desc_2_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_10_reg_we(uc2rb_wr_resp_desc_2_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_11_reg_we(uc2rb_wr_resp_desc_2_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_12_reg_we(uc2rb_wr_resp_desc_2_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_13_reg_we(uc2rb_wr_resp_desc_2_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_14_reg_we(uc2rb_wr_resp_desc_2_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_2_xuser_15_reg_we(uc2rb_wr_resp_desc_2_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_2_attr_reg_we(uc2rb_sn_req_desc_2_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_0_reg_we(uc2rb_sn_req_desc_2_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_1_reg_we(uc2rb_sn_req_desc_2_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_2_reg_we(uc2rb_sn_req_desc_2_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_2_acaddr_3_reg_we(uc2rb_sn_req_desc_2_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_data_offset_reg_we(uc2rb_rd_resp_desc_3_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_data_size_reg_we(uc2rb_rd_resp_desc_3_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_resp_reg_we(uc2rb_rd_resp_desc_3_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xid_0_reg_we(uc2rb_rd_resp_desc_3_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xid_1_reg_we(uc2rb_rd_resp_desc_3_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xid_2_reg_we(uc2rb_rd_resp_desc_3_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xid_3_reg_we(uc2rb_rd_resp_desc_3_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_0_reg_we(uc2rb_rd_resp_desc_3_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_1_reg_we(uc2rb_rd_resp_desc_3_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_2_reg_we(uc2rb_rd_resp_desc_3_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_3_reg_we(uc2rb_rd_resp_desc_3_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_4_reg_we(uc2rb_rd_resp_desc_3_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_5_reg_we(uc2rb_rd_resp_desc_3_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_6_reg_we(uc2rb_rd_resp_desc_3_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_7_reg_we(uc2rb_rd_resp_desc_3_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_8_reg_we(uc2rb_rd_resp_desc_3_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_9_reg_we(uc2rb_rd_resp_desc_3_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_10_reg_we(uc2rb_rd_resp_desc_3_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_11_reg_we(uc2rb_rd_resp_desc_3_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_12_reg_we(uc2rb_rd_resp_desc_3_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_13_reg_we(uc2rb_rd_resp_desc_3_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_14_reg_we(uc2rb_rd_resp_desc_3_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_3_xuser_15_reg_we(uc2rb_rd_resp_desc_3_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_resp_reg_we(uc2rb_wr_resp_desc_3_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xid_0_reg_we(uc2rb_wr_resp_desc_3_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xid_1_reg_we(uc2rb_wr_resp_desc_3_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xid_2_reg_we(uc2rb_wr_resp_desc_3_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xid_3_reg_we(uc2rb_wr_resp_desc_3_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_0_reg_we(uc2rb_wr_resp_desc_3_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_1_reg_we(uc2rb_wr_resp_desc_3_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_2_reg_we(uc2rb_wr_resp_desc_3_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_3_reg_we(uc2rb_wr_resp_desc_3_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_4_reg_we(uc2rb_wr_resp_desc_3_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_5_reg_we(uc2rb_wr_resp_desc_3_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_6_reg_we(uc2rb_wr_resp_desc_3_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_7_reg_we(uc2rb_wr_resp_desc_3_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_8_reg_we(uc2rb_wr_resp_desc_3_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_9_reg_we(uc2rb_wr_resp_desc_3_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_10_reg_we(uc2rb_wr_resp_desc_3_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_11_reg_we(uc2rb_wr_resp_desc_3_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_12_reg_we(uc2rb_wr_resp_desc_3_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_13_reg_we(uc2rb_wr_resp_desc_3_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_14_reg_we(uc2rb_wr_resp_desc_3_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_3_xuser_15_reg_we(uc2rb_wr_resp_desc_3_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_3_attr_reg_we(uc2rb_sn_req_desc_3_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_0_reg_we(uc2rb_sn_req_desc_3_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_1_reg_we(uc2rb_sn_req_desc_3_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_2_reg_we(uc2rb_sn_req_desc_3_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_3_acaddr_3_reg_we(uc2rb_sn_req_desc_3_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_data_offset_reg_we(uc2rb_rd_resp_desc_4_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_data_size_reg_we(uc2rb_rd_resp_desc_4_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_resp_reg_we(uc2rb_rd_resp_desc_4_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xid_0_reg_we(uc2rb_rd_resp_desc_4_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xid_1_reg_we(uc2rb_rd_resp_desc_4_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xid_2_reg_we(uc2rb_rd_resp_desc_4_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xid_3_reg_we(uc2rb_rd_resp_desc_4_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_0_reg_we(uc2rb_rd_resp_desc_4_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_1_reg_we(uc2rb_rd_resp_desc_4_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_2_reg_we(uc2rb_rd_resp_desc_4_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_3_reg_we(uc2rb_rd_resp_desc_4_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_4_reg_we(uc2rb_rd_resp_desc_4_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_5_reg_we(uc2rb_rd_resp_desc_4_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_6_reg_we(uc2rb_rd_resp_desc_4_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_7_reg_we(uc2rb_rd_resp_desc_4_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_8_reg_we(uc2rb_rd_resp_desc_4_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_9_reg_we(uc2rb_rd_resp_desc_4_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_10_reg_we(uc2rb_rd_resp_desc_4_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_11_reg_we(uc2rb_rd_resp_desc_4_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_12_reg_we(uc2rb_rd_resp_desc_4_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_13_reg_we(uc2rb_rd_resp_desc_4_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_14_reg_we(uc2rb_rd_resp_desc_4_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_4_xuser_15_reg_we(uc2rb_rd_resp_desc_4_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_resp_reg_we(uc2rb_wr_resp_desc_4_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xid_0_reg_we(uc2rb_wr_resp_desc_4_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xid_1_reg_we(uc2rb_wr_resp_desc_4_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xid_2_reg_we(uc2rb_wr_resp_desc_4_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xid_3_reg_we(uc2rb_wr_resp_desc_4_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_0_reg_we(uc2rb_wr_resp_desc_4_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_1_reg_we(uc2rb_wr_resp_desc_4_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_2_reg_we(uc2rb_wr_resp_desc_4_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_3_reg_we(uc2rb_wr_resp_desc_4_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_4_reg_we(uc2rb_wr_resp_desc_4_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_5_reg_we(uc2rb_wr_resp_desc_4_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_6_reg_we(uc2rb_wr_resp_desc_4_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_7_reg_we(uc2rb_wr_resp_desc_4_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_8_reg_we(uc2rb_wr_resp_desc_4_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_9_reg_we(uc2rb_wr_resp_desc_4_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_10_reg_we(uc2rb_wr_resp_desc_4_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_11_reg_we(uc2rb_wr_resp_desc_4_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_12_reg_we(uc2rb_wr_resp_desc_4_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_13_reg_we(uc2rb_wr_resp_desc_4_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_14_reg_we(uc2rb_wr_resp_desc_4_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_4_xuser_15_reg_we(uc2rb_wr_resp_desc_4_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_4_attr_reg_we(uc2rb_sn_req_desc_4_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_0_reg_we(uc2rb_sn_req_desc_4_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_1_reg_we(uc2rb_sn_req_desc_4_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_2_reg_we(uc2rb_sn_req_desc_4_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_4_acaddr_3_reg_we(uc2rb_sn_req_desc_4_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_data_offset_reg_we(uc2rb_rd_resp_desc_5_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_data_size_reg_we(uc2rb_rd_resp_desc_5_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_resp_reg_we(uc2rb_rd_resp_desc_5_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xid_0_reg_we(uc2rb_rd_resp_desc_5_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xid_1_reg_we(uc2rb_rd_resp_desc_5_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xid_2_reg_we(uc2rb_rd_resp_desc_5_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xid_3_reg_we(uc2rb_rd_resp_desc_5_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_0_reg_we(uc2rb_rd_resp_desc_5_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_1_reg_we(uc2rb_rd_resp_desc_5_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_2_reg_we(uc2rb_rd_resp_desc_5_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_3_reg_we(uc2rb_rd_resp_desc_5_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_4_reg_we(uc2rb_rd_resp_desc_5_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_5_reg_we(uc2rb_rd_resp_desc_5_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_6_reg_we(uc2rb_rd_resp_desc_5_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_7_reg_we(uc2rb_rd_resp_desc_5_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_8_reg_we(uc2rb_rd_resp_desc_5_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_9_reg_we(uc2rb_rd_resp_desc_5_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_10_reg_we(uc2rb_rd_resp_desc_5_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_11_reg_we(uc2rb_rd_resp_desc_5_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_12_reg_we(uc2rb_rd_resp_desc_5_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_13_reg_we(uc2rb_rd_resp_desc_5_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_14_reg_we(uc2rb_rd_resp_desc_5_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_5_xuser_15_reg_we(uc2rb_rd_resp_desc_5_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_resp_reg_we(uc2rb_wr_resp_desc_5_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xid_0_reg_we(uc2rb_wr_resp_desc_5_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xid_1_reg_we(uc2rb_wr_resp_desc_5_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xid_2_reg_we(uc2rb_wr_resp_desc_5_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xid_3_reg_we(uc2rb_wr_resp_desc_5_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_0_reg_we(uc2rb_wr_resp_desc_5_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_1_reg_we(uc2rb_wr_resp_desc_5_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_2_reg_we(uc2rb_wr_resp_desc_5_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_3_reg_we(uc2rb_wr_resp_desc_5_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_4_reg_we(uc2rb_wr_resp_desc_5_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_5_reg_we(uc2rb_wr_resp_desc_5_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_6_reg_we(uc2rb_wr_resp_desc_5_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_7_reg_we(uc2rb_wr_resp_desc_5_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_8_reg_we(uc2rb_wr_resp_desc_5_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_9_reg_we(uc2rb_wr_resp_desc_5_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_10_reg_we(uc2rb_wr_resp_desc_5_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_11_reg_we(uc2rb_wr_resp_desc_5_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_12_reg_we(uc2rb_wr_resp_desc_5_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_13_reg_we(uc2rb_wr_resp_desc_5_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_14_reg_we(uc2rb_wr_resp_desc_5_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_5_xuser_15_reg_we(uc2rb_wr_resp_desc_5_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_5_attr_reg_we(uc2rb_sn_req_desc_5_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_0_reg_we(uc2rb_sn_req_desc_5_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_1_reg_we(uc2rb_sn_req_desc_5_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_2_reg_we(uc2rb_sn_req_desc_5_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_5_acaddr_3_reg_we(uc2rb_sn_req_desc_5_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_data_offset_reg_we(uc2rb_rd_resp_desc_6_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_data_size_reg_we(uc2rb_rd_resp_desc_6_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_resp_reg_we(uc2rb_rd_resp_desc_6_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xid_0_reg_we(uc2rb_rd_resp_desc_6_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xid_1_reg_we(uc2rb_rd_resp_desc_6_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xid_2_reg_we(uc2rb_rd_resp_desc_6_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xid_3_reg_we(uc2rb_rd_resp_desc_6_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_0_reg_we(uc2rb_rd_resp_desc_6_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_1_reg_we(uc2rb_rd_resp_desc_6_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_2_reg_we(uc2rb_rd_resp_desc_6_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_3_reg_we(uc2rb_rd_resp_desc_6_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_4_reg_we(uc2rb_rd_resp_desc_6_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_5_reg_we(uc2rb_rd_resp_desc_6_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_6_reg_we(uc2rb_rd_resp_desc_6_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_7_reg_we(uc2rb_rd_resp_desc_6_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_8_reg_we(uc2rb_rd_resp_desc_6_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_9_reg_we(uc2rb_rd_resp_desc_6_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_10_reg_we(uc2rb_rd_resp_desc_6_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_11_reg_we(uc2rb_rd_resp_desc_6_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_12_reg_we(uc2rb_rd_resp_desc_6_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_13_reg_we(uc2rb_rd_resp_desc_6_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_14_reg_we(uc2rb_rd_resp_desc_6_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_6_xuser_15_reg_we(uc2rb_rd_resp_desc_6_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_resp_reg_we(uc2rb_wr_resp_desc_6_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xid_0_reg_we(uc2rb_wr_resp_desc_6_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xid_1_reg_we(uc2rb_wr_resp_desc_6_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xid_2_reg_we(uc2rb_wr_resp_desc_6_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xid_3_reg_we(uc2rb_wr_resp_desc_6_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_0_reg_we(uc2rb_wr_resp_desc_6_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_1_reg_we(uc2rb_wr_resp_desc_6_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_2_reg_we(uc2rb_wr_resp_desc_6_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_3_reg_we(uc2rb_wr_resp_desc_6_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_4_reg_we(uc2rb_wr_resp_desc_6_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_5_reg_we(uc2rb_wr_resp_desc_6_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_6_reg_we(uc2rb_wr_resp_desc_6_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_7_reg_we(uc2rb_wr_resp_desc_6_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_8_reg_we(uc2rb_wr_resp_desc_6_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_9_reg_we(uc2rb_wr_resp_desc_6_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_10_reg_we(uc2rb_wr_resp_desc_6_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_11_reg_we(uc2rb_wr_resp_desc_6_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_12_reg_we(uc2rb_wr_resp_desc_6_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_13_reg_we(uc2rb_wr_resp_desc_6_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_14_reg_we(uc2rb_wr_resp_desc_6_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_6_xuser_15_reg_we(uc2rb_wr_resp_desc_6_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_6_attr_reg_we(uc2rb_sn_req_desc_6_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_0_reg_we(uc2rb_sn_req_desc_6_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_1_reg_we(uc2rb_sn_req_desc_6_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_2_reg_we(uc2rb_sn_req_desc_6_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_6_acaddr_3_reg_we(uc2rb_sn_req_desc_6_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_data_offset_reg_we(uc2rb_rd_resp_desc_7_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_data_size_reg_we(uc2rb_rd_resp_desc_7_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_resp_reg_we(uc2rb_rd_resp_desc_7_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xid_0_reg_we(uc2rb_rd_resp_desc_7_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xid_1_reg_we(uc2rb_rd_resp_desc_7_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xid_2_reg_we(uc2rb_rd_resp_desc_7_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xid_3_reg_we(uc2rb_rd_resp_desc_7_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_0_reg_we(uc2rb_rd_resp_desc_7_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_1_reg_we(uc2rb_rd_resp_desc_7_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_2_reg_we(uc2rb_rd_resp_desc_7_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_3_reg_we(uc2rb_rd_resp_desc_7_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_4_reg_we(uc2rb_rd_resp_desc_7_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_5_reg_we(uc2rb_rd_resp_desc_7_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_6_reg_we(uc2rb_rd_resp_desc_7_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_7_reg_we(uc2rb_rd_resp_desc_7_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_8_reg_we(uc2rb_rd_resp_desc_7_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_9_reg_we(uc2rb_rd_resp_desc_7_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_10_reg_we(uc2rb_rd_resp_desc_7_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_11_reg_we(uc2rb_rd_resp_desc_7_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_12_reg_we(uc2rb_rd_resp_desc_7_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_13_reg_we(uc2rb_rd_resp_desc_7_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_14_reg_we(uc2rb_rd_resp_desc_7_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_7_xuser_15_reg_we(uc2rb_rd_resp_desc_7_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_resp_reg_we(uc2rb_wr_resp_desc_7_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xid_0_reg_we(uc2rb_wr_resp_desc_7_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xid_1_reg_we(uc2rb_wr_resp_desc_7_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xid_2_reg_we(uc2rb_wr_resp_desc_7_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xid_3_reg_we(uc2rb_wr_resp_desc_7_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_0_reg_we(uc2rb_wr_resp_desc_7_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_1_reg_we(uc2rb_wr_resp_desc_7_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_2_reg_we(uc2rb_wr_resp_desc_7_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_3_reg_we(uc2rb_wr_resp_desc_7_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_4_reg_we(uc2rb_wr_resp_desc_7_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_5_reg_we(uc2rb_wr_resp_desc_7_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_6_reg_we(uc2rb_wr_resp_desc_7_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_7_reg_we(uc2rb_wr_resp_desc_7_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_8_reg_we(uc2rb_wr_resp_desc_7_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_9_reg_we(uc2rb_wr_resp_desc_7_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_10_reg_we(uc2rb_wr_resp_desc_7_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_11_reg_we(uc2rb_wr_resp_desc_7_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_12_reg_we(uc2rb_wr_resp_desc_7_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_13_reg_we(uc2rb_wr_resp_desc_7_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_14_reg_we(uc2rb_wr_resp_desc_7_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_7_xuser_15_reg_we(uc2rb_wr_resp_desc_7_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_7_attr_reg_we(uc2rb_sn_req_desc_7_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_0_reg_we(uc2rb_sn_req_desc_7_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_1_reg_we(uc2rb_sn_req_desc_7_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_2_reg_we(uc2rb_sn_req_desc_7_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_7_acaddr_3_reg_we(uc2rb_sn_req_desc_7_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_data_offset_reg_we(uc2rb_rd_resp_desc_8_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_data_size_reg_we(uc2rb_rd_resp_desc_8_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_resp_reg_we(uc2rb_rd_resp_desc_8_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xid_0_reg_we(uc2rb_rd_resp_desc_8_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xid_1_reg_we(uc2rb_rd_resp_desc_8_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xid_2_reg_we(uc2rb_rd_resp_desc_8_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xid_3_reg_we(uc2rb_rd_resp_desc_8_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_0_reg_we(uc2rb_rd_resp_desc_8_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_1_reg_we(uc2rb_rd_resp_desc_8_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_2_reg_we(uc2rb_rd_resp_desc_8_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_3_reg_we(uc2rb_rd_resp_desc_8_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_4_reg_we(uc2rb_rd_resp_desc_8_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_5_reg_we(uc2rb_rd_resp_desc_8_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_6_reg_we(uc2rb_rd_resp_desc_8_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_7_reg_we(uc2rb_rd_resp_desc_8_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_8_reg_we(uc2rb_rd_resp_desc_8_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_9_reg_we(uc2rb_rd_resp_desc_8_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_10_reg_we(uc2rb_rd_resp_desc_8_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_11_reg_we(uc2rb_rd_resp_desc_8_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_12_reg_we(uc2rb_rd_resp_desc_8_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_13_reg_we(uc2rb_rd_resp_desc_8_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_14_reg_we(uc2rb_rd_resp_desc_8_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_8_xuser_15_reg_we(uc2rb_rd_resp_desc_8_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_resp_reg_we(uc2rb_wr_resp_desc_8_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xid_0_reg_we(uc2rb_wr_resp_desc_8_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xid_1_reg_we(uc2rb_wr_resp_desc_8_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xid_2_reg_we(uc2rb_wr_resp_desc_8_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xid_3_reg_we(uc2rb_wr_resp_desc_8_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_0_reg_we(uc2rb_wr_resp_desc_8_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_1_reg_we(uc2rb_wr_resp_desc_8_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_2_reg_we(uc2rb_wr_resp_desc_8_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_3_reg_we(uc2rb_wr_resp_desc_8_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_4_reg_we(uc2rb_wr_resp_desc_8_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_5_reg_we(uc2rb_wr_resp_desc_8_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_6_reg_we(uc2rb_wr_resp_desc_8_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_7_reg_we(uc2rb_wr_resp_desc_8_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_8_reg_we(uc2rb_wr_resp_desc_8_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_9_reg_we(uc2rb_wr_resp_desc_8_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_10_reg_we(uc2rb_wr_resp_desc_8_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_11_reg_we(uc2rb_wr_resp_desc_8_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_12_reg_we(uc2rb_wr_resp_desc_8_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_13_reg_we(uc2rb_wr_resp_desc_8_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_14_reg_we(uc2rb_wr_resp_desc_8_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_8_xuser_15_reg_we(uc2rb_wr_resp_desc_8_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_8_attr_reg_we(uc2rb_sn_req_desc_8_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_0_reg_we(uc2rb_sn_req_desc_8_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_1_reg_we(uc2rb_sn_req_desc_8_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_2_reg_we(uc2rb_sn_req_desc_8_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_8_acaddr_3_reg_we(uc2rb_sn_req_desc_8_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_data_offset_reg_we(uc2rb_rd_resp_desc_9_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_data_size_reg_we(uc2rb_rd_resp_desc_9_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_resp_reg_we(uc2rb_rd_resp_desc_9_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xid_0_reg_we(uc2rb_rd_resp_desc_9_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xid_1_reg_we(uc2rb_rd_resp_desc_9_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xid_2_reg_we(uc2rb_rd_resp_desc_9_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xid_3_reg_we(uc2rb_rd_resp_desc_9_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_0_reg_we(uc2rb_rd_resp_desc_9_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_1_reg_we(uc2rb_rd_resp_desc_9_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_2_reg_we(uc2rb_rd_resp_desc_9_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_3_reg_we(uc2rb_rd_resp_desc_9_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_4_reg_we(uc2rb_rd_resp_desc_9_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_5_reg_we(uc2rb_rd_resp_desc_9_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_6_reg_we(uc2rb_rd_resp_desc_9_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_7_reg_we(uc2rb_rd_resp_desc_9_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_8_reg_we(uc2rb_rd_resp_desc_9_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_9_reg_we(uc2rb_rd_resp_desc_9_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_10_reg_we(uc2rb_rd_resp_desc_9_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_11_reg_we(uc2rb_rd_resp_desc_9_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_12_reg_we(uc2rb_rd_resp_desc_9_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_13_reg_we(uc2rb_rd_resp_desc_9_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_14_reg_we(uc2rb_rd_resp_desc_9_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_9_xuser_15_reg_we(uc2rb_rd_resp_desc_9_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_resp_reg_we(uc2rb_wr_resp_desc_9_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xid_0_reg_we(uc2rb_wr_resp_desc_9_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xid_1_reg_we(uc2rb_wr_resp_desc_9_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xid_2_reg_we(uc2rb_wr_resp_desc_9_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xid_3_reg_we(uc2rb_wr_resp_desc_9_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_0_reg_we(uc2rb_wr_resp_desc_9_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_1_reg_we(uc2rb_wr_resp_desc_9_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_2_reg_we(uc2rb_wr_resp_desc_9_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_3_reg_we(uc2rb_wr_resp_desc_9_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_4_reg_we(uc2rb_wr_resp_desc_9_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_5_reg_we(uc2rb_wr_resp_desc_9_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_6_reg_we(uc2rb_wr_resp_desc_9_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_7_reg_we(uc2rb_wr_resp_desc_9_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_8_reg_we(uc2rb_wr_resp_desc_9_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_9_reg_we(uc2rb_wr_resp_desc_9_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_10_reg_we(uc2rb_wr_resp_desc_9_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_11_reg_we(uc2rb_wr_resp_desc_9_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_12_reg_we(uc2rb_wr_resp_desc_9_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_13_reg_we(uc2rb_wr_resp_desc_9_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_14_reg_we(uc2rb_wr_resp_desc_9_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_9_xuser_15_reg_we(uc2rb_wr_resp_desc_9_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_9_attr_reg_we(uc2rb_sn_req_desc_9_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_0_reg_we(uc2rb_sn_req_desc_9_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_1_reg_we(uc2rb_sn_req_desc_9_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_2_reg_we(uc2rb_sn_req_desc_9_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_9_acaddr_3_reg_we(uc2rb_sn_req_desc_9_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_data_offset_reg_we(uc2rb_rd_resp_desc_a_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_data_size_reg_we(uc2rb_rd_resp_desc_a_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_resp_reg_we(uc2rb_rd_resp_desc_a_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xid_0_reg_we(uc2rb_rd_resp_desc_a_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xid_1_reg_we(uc2rb_rd_resp_desc_a_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xid_2_reg_we(uc2rb_rd_resp_desc_a_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xid_3_reg_we(uc2rb_rd_resp_desc_a_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_0_reg_we(uc2rb_rd_resp_desc_a_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_1_reg_we(uc2rb_rd_resp_desc_a_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_2_reg_we(uc2rb_rd_resp_desc_a_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_3_reg_we(uc2rb_rd_resp_desc_a_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_4_reg_we(uc2rb_rd_resp_desc_a_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_5_reg_we(uc2rb_rd_resp_desc_a_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_6_reg_we(uc2rb_rd_resp_desc_a_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_7_reg_we(uc2rb_rd_resp_desc_a_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_8_reg_we(uc2rb_rd_resp_desc_a_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_9_reg_we(uc2rb_rd_resp_desc_a_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_10_reg_we(uc2rb_rd_resp_desc_a_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_11_reg_we(uc2rb_rd_resp_desc_a_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_12_reg_we(uc2rb_rd_resp_desc_a_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_13_reg_we(uc2rb_rd_resp_desc_a_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_14_reg_we(uc2rb_rd_resp_desc_a_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_a_xuser_15_reg_we(uc2rb_rd_resp_desc_a_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_resp_reg_we(uc2rb_wr_resp_desc_a_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xid_0_reg_we(uc2rb_wr_resp_desc_a_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xid_1_reg_we(uc2rb_wr_resp_desc_a_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xid_2_reg_we(uc2rb_wr_resp_desc_a_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xid_3_reg_we(uc2rb_wr_resp_desc_a_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_0_reg_we(uc2rb_wr_resp_desc_a_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_1_reg_we(uc2rb_wr_resp_desc_a_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_2_reg_we(uc2rb_wr_resp_desc_a_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_3_reg_we(uc2rb_wr_resp_desc_a_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_4_reg_we(uc2rb_wr_resp_desc_a_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_5_reg_we(uc2rb_wr_resp_desc_a_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_6_reg_we(uc2rb_wr_resp_desc_a_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_7_reg_we(uc2rb_wr_resp_desc_a_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_8_reg_we(uc2rb_wr_resp_desc_a_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_9_reg_we(uc2rb_wr_resp_desc_a_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_10_reg_we(uc2rb_wr_resp_desc_a_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_11_reg_we(uc2rb_wr_resp_desc_a_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_12_reg_we(uc2rb_wr_resp_desc_a_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_13_reg_we(uc2rb_wr_resp_desc_a_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_14_reg_we(uc2rb_wr_resp_desc_a_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_a_xuser_15_reg_we(uc2rb_wr_resp_desc_a_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_a_attr_reg_we(uc2rb_sn_req_desc_a_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_0_reg_we(uc2rb_sn_req_desc_a_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_1_reg_we(uc2rb_sn_req_desc_a_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_2_reg_we(uc2rb_sn_req_desc_a_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_a_acaddr_3_reg_we(uc2rb_sn_req_desc_a_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_data_offset_reg_we(uc2rb_rd_resp_desc_b_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_data_size_reg_we(uc2rb_rd_resp_desc_b_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_resp_reg_we(uc2rb_rd_resp_desc_b_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xid_0_reg_we(uc2rb_rd_resp_desc_b_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xid_1_reg_we(uc2rb_rd_resp_desc_b_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xid_2_reg_we(uc2rb_rd_resp_desc_b_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xid_3_reg_we(uc2rb_rd_resp_desc_b_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_0_reg_we(uc2rb_rd_resp_desc_b_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_1_reg_we(uc2rb_rd_resp_desc_b_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_2_reg_we(uc2rb_rd_resp_desc_b_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_3_reg_we(uc2rb_rd_resp_desc_b_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_4_reg_we(uc2rb_rd_resp_desc_b_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_5_reg_we(uc2rb_rd_resp_desc_b_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_6_reg_we(uc2rb_rd_resp_desc_b_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_7_reg_we(uc2rb_rd_resp_desc_b_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_8_reg_we(uc2rb_rd_resp_desc_b_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_9_reg_we(uc2rb_rd_resp_desc_b_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_10_reg_we(uc2rb_rd_resp_desc_b_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_11_reg_we(uc2rb_rd_resp_desc_b_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_12_reg_we(uc2rb_rd_resp_desc_b_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_13_reg_we(uc2rb_rd_resp_desc_b_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_14_reg_we(uc2rb_rd_resp_desc_b_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_b_xuser_15_reg_we(uc2rb_rd_resp_desc_b_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_resp_reg_we(uc2rb_wr_resp_desc_b_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xid_0_reg_we(uc2rb_wr_resp_desc_b_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xid_1_reg_we(uc2rb_wr_resp_desc_b_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xid_2_reg_we(uc2rb_wr_resp_desc_b_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xid_3_reg_we(uc2rb_wr_resp_desc_b_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_0_reg_we(uc2rb_wr_resp_desc_b_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_1_reg_we(uc2rb_wr_resp_desc_b_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_2_reg_we(uc2rb_wr_resp_desc_b_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_3_reg_we(uc2rb_wr_resp_desc_b_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_4_reg_we(uc2rb_wr_resp_desc_b_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_5_reg_we(uc2rb_wr_resp_desc_b_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_6_reg_we(uc2rb_wr_resp_desc_b_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_7_reg_we(uc2rb_wr_resp_desc_b_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_8_reg_we(uc2rb_wr_resp_desc_b_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_9_reg_we(uc2rb_wr_resp_desc_b_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_10_reg_we(uc2rb_wr_resp_desc_b_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_11_reg_we(uc2rb_wr_resp_desc_b_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_12_reg_we(uc2rb_wr_resp_desc_b_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_13_reg_we(uc2rb_wr_resp_desc_b_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_14_reg_we(uc2rb_wr_resp_desc_b_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_b_xuser_15_reg_we(uc2rb_wr_resp_desc_b_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_b_attr_reg_we(uc2rb_sn_req_desc_b_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_0_reg_we(uc2rb_sn_req_desc_b_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_1_reg_we(uc2rb_sn_req_desc_b_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_2_reg_we(uc2rb_sn_req_desc_b_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_b_acaddr_3_reg_we(uc2rb_sn_req_desc_b_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_data_offset_reg_we(uc2rb_rd_resp_desc_c_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_data_size_reg_we(uc2rb_rd_resp_desc_c_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_resp_reg_we(uc2rb_rd_resp_desc_c_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xid_0_reg_we(uc2rb_rd_resp_desc_c_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xid_1_reg_we(uc2rb_rd_resp_desc_c_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xid_2_reg_we(uc2rb_rd_resp_desc_c_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xid_3_reg_we(uc2rb_rd_resp_desc_c_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_0_reg_we(uc2rb_rd_resp_desc_c_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_1_reg_we(uc2rb_rd_resp_desc_c_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_2_reg_we(uc2rb_rd_resp_desc_c_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_3_reg_we(uc2rb_rd_resp_desc_c_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_4_reg_we(uc2rb_rd_resp_desc_c_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_5_reg_we(uc2rb_rd_resp_desc_c_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_6_reg_we(uc2rb_rd_resp_desc_c_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_7_reg_we(uc2rb_rd_resp_desc_c_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_8_reg_we(uc2rb_rd_resp_desc_c_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_9_reg_we(uc2rb_rd_resp_desc_c_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_10_reg_we(uc2rb_rd_resp_desc_c_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_11_reg_we(uc2rb_rd_resp_desc_c_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_12_reg_we(uc2rb_rd_resp_desc_c_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_13_reg_we(uc2rb_rd_resp_desc_c_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_14_reg_we(uc2rb_rd_resp_desc_c_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_c_xuser_15_reg_we(uc2rb_rd_resp_desc_c_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_resp_reg_we(uc2rb_wr_resp_desc_c_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xid_0_reg_we(uc2rb_wr_resp_desc_c_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xid_1_reg_we(uc2rb_wr_resp_desc_c_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xid_2_reg_we(uc2rb_wr_resp_desc_c_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xid_3_reg_we(uc2rb_wr_resp_desc_c_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_0_reg_we(uc2rb_wr_resp_desc_c_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_1_reg_we(uc2rb_wr_resp_desc_c_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_2_reg_we(uc2rb_wr_resp_desc_c_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_3_reg_we(uc2rb_wr_resp_desc_c_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_4_reg_we(uc2rb_wr_resp_desc_c_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_5_reg_we(uc2rb_wr_resp_desc_c_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_6_reg_we(uc2rb_wr_resp_desc_c_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_7_reg_we(uc2rb_wr_resp_desc_c_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_8_reg_we(uc2rb_wr_resp_desc_c_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_9_reg_we(uc2rb_wr_resp_desc_c_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_10_reg_we(uc2rb_wr_resp_desc_c_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_11_reg_we(uc2rb_wr_resp_desc_c_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_12_reg_we(uc2rb_wr_resp_desc_c_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_13_reg_we(uc2rb_wr_resp_desc_c_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_14_reg_we(uc2rb_wr_resp_desc_c_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_c_xuser_15_reg_we(uc2rb_wr_resp_desc_c_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_c_attr_reg_we(uc2rb_sn_req_desc_c_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_0_reg_we(uc2rb_sn_req_desc_c_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_1_reg_we(uc2rb_sn_req_desc_c_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_2_reg_we(uc2rb_sn_req_desc_c_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_c_acaddr_3_reg_we(uc2rb_sn_req_desc_c_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_data_offset_reg_we(uc2rb_rd_resp_desc_d_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_data_size_reg_we(uc2rb_rd_resp_desc_d_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_resp_reg_we(uc2rb_rd_resp_desc_d_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xid_0_reg_we(uc2rb_rd_resp_desc_d_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xid_1_reg_we(uc2rb_rd_resp_desc_d_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xid_2_reg_we(uc2rb_rd_resp_desc_d_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xid_3_reg_we(uc2rb_rd_resp_desc_d_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_0_reg_we(uc2rb_rd_resp_desc_d_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_1_reg_we(uc2rb_rd_resp_desc_d_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_2_reg_we(uc2rb_rd_resp_desc_d_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_3_reg_we(uc2rb_rd_resp_desc_d_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_4_reg_we(uc2rb_rd_resp_desc_d_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_5_reg_we(uc2rb_rd_resp_desc_d_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_6_reg_we(uc2rb_rd_resp_desc_d_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_7_reg_we(uc2rb_rd_resp_desc_d_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_8_reg_we(uc2rb_rd_resp_desc_d_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_9_reg_we(uc2rb_rd_resp_desc_d_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_10_reg_we(uc2rb_rd_resp_desc_d_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_11_reg_we(uc2rb_rd_resp_desc_d_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_12_reg_we(uc2rb_rd_resp_desc_d_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_13_reg_we(uc2rb_rd_resp_desc_d_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_14_reg_we(uc2rb_rd_resp_desc_d_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_d_xuser_15_reg_we(uc2rb_rd_resp_desc_d_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_resp_reg_we(uc2rb_wr_resp_desc_d_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xid_0_reg_we(uc2rb_wr_resp_desc_d_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xid_1_reg_we(uc2rb_wr_resp_desc_d_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xid_2_reg_we(uc2rb_wr_resp_desc_d_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xid_3_reg_we(uc2rb_wr_resp_desc_d_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_0_reg_we(uc2rb_wr_resp_desc_d_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_1_reg_we(uc2rb_wr_resp_desc_d_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_2_reg_we(uc2rb_wr_resp_desc_d_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_3_reg_we(uc2rb_wr_resp_desc_d_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_4_reg_we(uc2rb_wr_resp_desc_d_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_5_reg_we(uc2rb_wr_resp_desc_d_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_6_reg_we(uc2rb_wr_resp_desc_d_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_7_reg_we(uc2rb_wr_resp_desc_d_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_8_reg_we(uc2rb_wr_resp_desc_d_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_9_reg_we(uc2rb_wr_resp_desc_d_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_10_reg_we(uc2rb_wr_resp_desc_d_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_11_reg_we(uc2rb_wr_resp_desc_d_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_12_reg_we(uc2rb_wr_resp_desc_d_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_13_reg_we(uc2rb_wr_resp_desc_d_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_14_reg_we(uc2rb_wr_resp_desc_d_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_d_xuser_15_reg_we(uc2rb_wr_resp_desc_d_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_d_attr_reg_we(uc2rb_sn_req_desc_d_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_0_reg_we(uc2rb_sn_req_desc_d_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_1_reg_we(uc2rb_sn_req_desc_d_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_2_reg_we(uc2rb_sn_req_desc_d_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_d_acaddr_3_reg_we(uc2rb_sn_req_desc_d_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_data_offset_reg_we(uc2rb_rd_resp_desc_e_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_data_size_reg_we(uc2rb_rd_resp_desc_e_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_resp_reg_we(uc2rb_rd_resp_desc_e_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xid_0_reg_we(uc2rb_rd_resp_desc_e_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xid_1_reg_we(uc2rb_rd_resp_desc_e_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xid_2_reg_we(uc2rb_rd_resp_desc_e_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xid_3_reg_we(uc2rb_rd_resp_desc_e_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_0_reg_we(uc2rb_rd_resp_desc_e_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_1_reg_we(uc2rb_rd_resp_desc_e_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_2_reg_we(uc2rb_rd_resp_desc_e_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_3_reg_we(uc2rb_rd_resp_desc_e_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_4_reg_we(uc2rb_rd_resp_desc_e_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_5_reg_we(uc2rb_rd_resp_desc_e_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_6_reg_we(uc2rb_rd_resp_desc_e_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_7_reg_we(uc2rb_rd_resp_desc_e_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_8_reg_we(uc2rb_rd_resp_desc_e_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_9_reg_we(uc2rb_rd_resp_desc_e_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_10_reg_we(uc2rb_rd_resp_desc_e_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_11_reg_we(uc2rb_rd_resp_desc_e_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_12_reg_we(uc2rb_rd_resp_desc_e_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_13_reg_we(uc2rb_rd_resp_desc_e_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_14_reg_we(uc2rb_rd_resp_desc_e_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_e_xuser_15_reg_we(uc2rb_rd_resp_desc_e_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_resp_reg_we(uc2rb_wr_resp_desc_e_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xid_0_reg_we(uc2rb_wr_resp_desc_e_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xid_1_reg_we(uc2rb_wr_resp_desc_e_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xid_2_reg_we(uc2rb_wr_resp_desc_e_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xid_3_reg_we(uc2rb_wr_resp_desc_e_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_0_reg_we(uc2rb_wr_resp_desc_e_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_1_reg_we(uc2rb_wr_resp_desc_e_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_2_reg_we(uc2rb_wr_resp_desc_e_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_3_reg_we(uc2rb_wr_resp_desc_e_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_4_reg_we(uc2rb_wr_resp_desc_e_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_5_reg_we(uc2rb_wr_resp_desc_e_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_6_reg_we(uc2rb_wr_resp_desc_e_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_7_reg_we(uc2rb_wr_resp_desc_e_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_8_reg_we(uc2rb_wr_resp_desc_e_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_9_reg_we(uc2rb_wr_resp_desc_e_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_10_reg_we(uc2rb_wr_resp_desc_e_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_11_reg_we(uc2rb_wr_resp_desc_e_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_12_reg_we(uc2rb_wr_resp_desc_e_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_13_reg_we(uc2rb_wr_resp_desc_e_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_14_reg_we(uc2rb_wr_resp_desc_e_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_e_xuser_15_reg_we(uc2rb_wr_resp_desc_e_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_e_attr_reg_we(uc2rb_sn_req_desc_e_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_0_reg_we(uc2rb_sn_req_desc_e_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_1_reg_we(uc2rb_sn_req_desc_e_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_2_reg_we(uc2rb_sn_req_desc_e_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_e_acaddr_3_reg_we(uc2rb_sn_req_desc_e_acaddr_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_data_offset_reg_we(uc2rb_rd_resp_desc_f_data_offset_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_data_size_reg_we(uc2rb_rd_resp_desc_f_data_size_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_resp_reg_we(uc2rb_rd_resp_desc_f_resp_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xid_0_reg_we(uc2rb_rd_resp_desc_f_xid_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xid_1_reg_we(uc2rb_rd_resp_desc_f_xid_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xid_2_reg_we(uc2rb_rd_resp_desc_f_xid_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xid_3_reg_we(uc2rb_rd_resp_desc_f_xid_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_0_reg_we(uc2rb_rd_resp_desc_f_xuser_0_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_1_reg_we(uc2rb_rd_resp_desc_f_xuser_1_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_2_reg_we(uc2rb_rd_resp_desc_f_xuser_2_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_3_reg_we(uc2rb_rd_resp_desc_f_xuser_3_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_4_reg_we(uc2rb_rd_resp_desc_f_xuser_4_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_5_reg_we(uc2rb_rd_resp_desc_f_xuser_5_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_6_reg_we(uc2rb_rd_resp_desc_f_xuser_6_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_7_reg_we(uc2rb_rd_resp_desc_f_xuser_7_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_8_reg_we(uc2rb_rd_resp_desc_f_xuser_8_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_9_reg_we(uc2rb_rd_resp_desc_f_xuser_9_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_10_reg_we(uc2rb_rd_resp_desc_f_xuser_10_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_11_reg_we(uc2rb_rd_resp_desc_f_xuser_11_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_12_reg_we(uc2rb_rd_resp_desc_f_xuser_12_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_13_reg_we(uc2rb_rd_resp_desc_f_xuser_13_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_14_reg_we(uc2rb_rd_resp_desc_f_xuser_14_reg_we),
                                                                                               .uc2rb_rd_resp_desc_f_xuser_15_reg_we(uc2rb_rd_resp_desc_f_xuser_15_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_resp_reg_we(uc2rb_wr_resp_desc_f_resp_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xid_0_reg_we(uc2rb_wr_resp_desc_f_xid_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xid_1_reg_we(uc2rb_wr_resp_desc_f_xid_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xid_2_reg_we(uc2rb_wr_resp_desc_f_xid_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xid_3_reg_we(uc2rb_wr_resp_desc_f_xid_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_0_reg_we(uc2rb_wr_resp_desc_f_xuser_0_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_1_reg_we(uc2rb_wr_resp_desc_f_xuser_1_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_2_reg_we(uc2rb_wr_resp_desc_f_xuser_2_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_3_reg_we(uc2rb_wr_resp_desc_f_xuser_3_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_4_reg_we(uc2rb_wr_resp_desc_f_xuser_4_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_5_reg_we(uc2rb_wr_resp_desc_f_xuser_5_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_6_reg_we(uc2rb_wr_resp_desc_f_xuser_6_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_7_reg_we(uc2rb_wr_resp_desc_f_xuser_7_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_8_reg_we(uc2rb_wr_resp_desc_f_xuser_8_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_9_reg_we(uc2rb_wr_resp_desc_f_xuser_9_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_10_reg_we(uc2rb_wr_resp_desc_f_xuser_10_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_11_reg_we(uc2rb_wr_resp_desc_f_xuser_11_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_12_reg_we(uc2rb_wr_resp_desc_f_xuser_12_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_13_reg_we(uc2rb_wr_resp_desc_f_xuser_13_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_14_reg_we(uc2rb_wr_resp_desc_f_xuser_14_reg_we),
                                                                                               .uc2rb_wr_resp_desc_f_xuser_15_reg_we(uc2rb_wr_resp_desc_f_xuser_15_reg_we),
                                                                                               .uc2rb_sn_req_desc_f_attr_reg_we(uc2rb_sn_req_desc_f_attr_reg_we),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_0_reg_we(uc2rb_sn_req_desc_f_acaddr_0_reg_we),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_1_reg_we(uc2rb_sn_req_desc_f_acaddr_1_reg_we),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_2_reg_we(uc2rb_sn_req_desc_f_acaddr_2_reg_we),
                                                                                               .uc2rb_sn_req_desc_f_acaddr_3_reg_we(uc2rb_sn_req_desc_f_acaddr_3_reg_we),
                                                                                               .uc2rb_wr_we        (uc2rb_wr_we),
                                                                                               .uc2rb_wr_bwe       (uc2rb_wr_bwe),
                                                                                               .uc2rb_wr_addr      (uc2rb_wr_addr),
                                                                                               .uc2rb_wr_data      (uc2rb_wr_data),
                                                                                               .uc2rb_rd_addr      (uc2rb_rd_addr),
                                                                                               .uc2rb_sn_addr      (uc2rb_sn_addr),
                                                                                               .rd_uc2hm_trig      (rd_uc2hm_trig),
                                                                                               .wr_uc2hm_trig      (wr_uc2hm_trig),
                                                                                               .rd_resp_fifo_out   (rd_resp_fifo_out),
                                                                                               .rd_resp_fifo_out_valid(rd_resp_fifo_out_valid),
                                                                                               .wr_resp_fifo_out   (wr_resp_fifo_out),
                                                                                               .wr_resp_fifo_out_valid(wr_resp_fifo_out_valid),
                                                                                               .sn_req_fifo_out    (sn_req_fifo_out),
                                                                                               .sn_req_fifo_out_valid(sn_req_fifo_out_valid),
                                                                                               // Inputs
                                                                                               .clk                (clk),
                                                                                               .resetn             (resetn),
                                                                                               .m_ace_usr_awready  (m_ace_usr_awready),
                                                                                               .m_ace_usr_wready   (m_ace_usr_wready),
                                                                                               .m_ace_usr_bid      (m_ace_usr_bid),
                                                                                               .m_ace_usr_bresp    (m_ace_usr_bresp),
                                                                                               .m_ace_usr_buser    (m_ace_usr_buser),
                                                                                               .m_ace_usr_bvalid   (m_ace_usr_bvalid),
                                                                                               .m_ace_usr_arready  (m_ace_usr_arready),
                                                                                               .m_ace_usr_rid      (m_ace_usr_rid),
                                                                                               .m_ace_usr_rdata    (m_ace_usr_rdata),
                                                                                               .m_ace_usr_rresp    (m_ace_usr_rresp),
                                                                                               .m_ace_usr_rlast    (m_ace_usr_rlast),
                                                                                               .m_ace_usr_ruser    (m_ace_usr_ruser),
                                                                                               .m_ace_usr_rvalid   (m_ace_usr_rvalid),
                                                                                               .m_ace_usr_acaddr   (m_ace_usr_acaddr),
                                                                                               .m_ace_usr_acsnoop  (m_ace_usr_acsnoop),
                                                                                               .m_ace_usr_acprot   (m_ace_usr_acprot),
                                                                                               .m_ace_usr_acvalid  (m_ace_usr_acvalid),
                                                                                               .m_ace_usr_crready  (m_ace_usr_crready),
                                                                                               .m_ace_usr_cdready  (m_ace_usr_cdready),
                                                                                               .bridge_identification_reg(bridge_identification_reg),
                                                                                               .last_bridge_reg    (last_bridge_reg),
                                                                                               .version_reg        (version_reg),
                                                                                               .bridge_type_reg    (bridge_type_reg),
                                                                                               .mode_select_reg    (mode_select_reg),
                                                                                               .reset_reg          (reset_reg),
                                                                                               .h2c_intr_0_reg     (h2c_intr_0_reg),
                                                                                               .h2c_intr_1_reg     (h2c_intr_1_reg),
                                                                                               .h2c_intr_2_reg     (h2c_intr_2_reg),
                                                                                               .h2c_intr_3_reg     (h2c_intr_3_reg),
                                                                                               .c2h_intr_status_0_reg(c2h_intr_status_0_reg),
                                                                                               .intr_c2h_toggle_status_0_reg(intr_c2h_toggle_status_0_reg),
                                                                                               .intr_c2h_toggle_clear_0_reg(intr_c2h_toggle_clear_0_reg),
                                                                                               .intr_c2h_toggle_enable_0_reg(intr_c2h_toggle_enable_0_reg),
                                                                                               .c2h_intr_status_1_reg(c2h_intr_status_1_reg),
                                                                                               .intr_c2h_toggle_status_1_reg(intr_c2h_toggle_status_1_reg),
                                                                                               .intr_c2h_toggle_clear_1_reg(intr_c2h_toggle_clear_1_reg),
                                                                                               .intr_c2h_toggle_enable_1_reg(intr_c2h_toggle_enable_1_reg),
                                                                                               .c2h_gpio_0_reg     (c2h_gpio_0_reg),
                                                                                               .c2h_gpio_1_reg     (c2h_gpio_1_reg),
                                                                                               .c2h_gpio_2_reg     (c2h_gpio_2_reg),
                                                                                               .c2h_gpio_3_reg     (c2h_gpio_3_reg),
                                                                                               .c2h_gpio_4_reg     (c2h_gpio_4_reg),
                                                                                               .c2h_gpio_5_reg     (c2h_gpio_5_reg),
                                                                                               .c2h_gpio_6_reg     (c2h_gpio_6_reg),
                                                                                               .c2h_gpio_7_reg     (c2h_gpio_7_reg),
                                                                                               .c2h_gpio_8_reg     (c2h_gpio_8_reg),
                                                                                               .c2h_gpio_9_reg     (c2h_gpio_9_reg),
                                                                                               .c2h_gpio_10_reg    (c2h_gpio_10_reg),
                                                                                               .c2h_gpio_11_reg    (c2h_gpio_11_reg),
                                                                                               .c2h_gpio_12_reg    (c2h_gpio_12_reg),
                                                                                               .c2h_gpio_13_reg    (c2h_gpio_13_reg),
                                                                                               .c2h_gpio_14_reg    (c2h_gpio_14_reg),
                                                                                               .c2h_gpio_15_reg    (c2h_gpio_15_reg),
                                                                                               .h2c_gpio_0_reg     (h2c_gpio_0_reg),
                                                                                               .h2c_gpio_1_reg     (h2c_gpio_1_reg),
                                                                                               .h2c_gpio_2_reg     (h2c_gpio_2_reg),
                                                                                               .h2c_gpio_3_reg     (h2c_gpio_3_reg),
                                                                                               .h2c_gpio_4_reg     (h2c_gpio_4_reg),
                                                                                               .h2c_gpio_5_reg     (h2c_gpio_5_reg),
                                                                                               .h2c_gpio_6_reg     (h2c_gpio_6_reg),
                                                                                               .h2c_gpio_7_reg     (h2c_gpio_7_reg),
                                                                                               .h2c_gpio_8_reg     (h2c_gpio_8_reg),
                                                                                               .h2c_gpio_9_reg     (h2c_gpio_9_reg),
                                                                                               .h2c_gpio_10_reg    (h2c_gpio_10_reg),
                                                                                               .h2c_gpio_11_reg    (h2c_gpio_11_reg),
                                                                                               .h2c_gpio_12_reg    (h2c_gpio_12_reg),
                                                                                               .h2c_gpio_13_reg    (h2c_gpio_13_reg),
                                                                                               .h2c_gpio_14_reg    (h2c_gpio_14_reg),
                                                                                               .h2c_gpio_15_reg    (h2c_gpio_15_reg),
                                                                                               .bridge_config_reg  (bridge_config_reg),
                                                                                               .intr_status_reg    (intr_status_reg),
                                                                                               .intr_error_status_reg(intr_error_status_reg),
                                                                                               .intr_error_clear_reg(intr_error_clear_reg),
                                                                                               .intr_error_enable_reg(intr_error_enable_reg),
                                                                                               .bridge_rd_user_config_reg(bridge_rd_user_config_reg),
                                                                                               .bridge_wr_user_config_reg(bridge_wr_user_config_reg),
                                                                                               .rd_max_desc_reg    (rd_max_desc_reg),
                                                                                               .wr_max_desc_reg    (wr_max_desc_reg),
                                                                                               .sn_max_desc_reg    (sn_max_desc_reg),
                                                                                               .rd_req_fifo_push_desc_reg(rd_req_fifo_push_desc_reg),
                                                                                               .rd_req_fifo_free_level_reg(rd_req_fifo_free_level_reg),
                                                                                               .rd_req_intr_comp_status_reg(rd_req_intr_comp_status_reg),
                                                                                               .rd_req_intr_comp_clear_reg(rd_req_intr_comp_clear_reg),
                                                                                               .rd_req_intr_comp_enable_reg(rd_req_intr_comp_enable_reg),
                                                                                               .rd_resp_free_desc_reg(rd_resp_free_desc_reg),
                                                                                               .rd_resp_fifo_pop_desc_reg(rd_resp_fifo_pop_desc_reg),
                                                                                               .rd_resp_fifo_fill_level_reg(rd_resp_fifo_fill_level_reg),
                                                                                               .wr_req_fifo_push_desc_reg(wr_req_fifo_push_desc_reg),
                                                                                               .wr_req_fifo_free_level_reg(wr_req_fifo_free_level_reg),
                                                                                               .wr_req_intr_comp_status_reg(wr_req_intr_comp_status_reg),
                                                                                               .wr_req_intr_comp_clear_reg(wr_req_intr_comp_clear_reg),
                                                                                               .wr_req_intr_comp_enable_reg(wr_req_intr_comp_enable_reg),
                                                                                               .wr_resp_free_desc_reg(wr_resp_free_desc_reg),
                                                                                               .wr_resp_fifo_pop_desc_reg(wr_resp_fifo_pop_desc_reg),
                                                                                               .wr_resp_fifo_fill_level_reg(wr_resp_fifo_fill_level_reg),
                                                                                               .sn_req_free_desc_reg(sn_req_free_desc_reg),
                                                                                               .sn_req_fifo_pop_desc_reg(sn_req_fifo_pop_desc_reg),
                                                                                               .sn_req_fifo_fill_level_reg(sn_req_fifo_fill_level_reg),
                                                                                               .sn_resp_fifo_push_desc_reg(sn_resp_fifo_push_desc_reg),
                                                                                               .sn_resp_fifo_free_level_reg(sn_resp_fifo_free_level_reg),
                                                                                               .sn_resp_intr_comp_status_reg(sn_resp_intr_comp_status_reg),
                                                                                               .sn_resp_intr_comp_clear_reg(sn_resp_intr_comp_clear_reg),
                                                                                               .sn_resp_intr_comp_enable_reg(sn_resp_intr_comp_enable_reg),
                                                                                               .sn_data_fifo_push_desc_reg(sn_data_fifo_push_desc_reg),
                                                                                               .sn_data_fifo_free_level_reg(sn_data_fifo_free_level_reg),
                                                                                               .sn_data_intr_comp_status_reg(sn_data_intr_comp_status_reg),
                                                                                               .sn_data_intr_comp_clear_reg(sn_data_intr_comp_clear_reg),
                                                                                               .sn_data_intr_comp_enable_reg(sn_data_intr_comp_enable_reg),
                                                                                               .intr_fifo_enable_reg(intr_fifo_enable_reg),
                                                                                               .rd_req_desc_0_txn_type_reg(rd_req_desc_0_txn_type_reg),
                                                                                               .rd_req_desc_0_size_reg(rd_req_desc_0_size_reg),
                                                                                               .rd_req_desc_0_axsize_reg(rd_req_desc_0_axsize_reg),
                                                                                               .rd_req_desc_0_attr_reg(rd_req_desc_0_attr_reg),
                                                                                               .rd_req_desc_0_axaddr_0_reg(rd_req_desc_0_axaddr_0_reg),
                                                                                               .rd_req_desc_0_axaddr_1_reg(rd_req_desc_0_axaddr_1_reg),
                                                                                               .rd_req_desc_0_axaddr_2_reg(rd_req_desc_0_axaddr_2_reg),
                                                                                               .rd_req_desc_0_axaddr_3_reg(rd_req_desc_0_axaddr_3_reg),
                                                                                               .rd_req_desc_0_axid_0_reg(rd_req_desc_0_axid_0_reg),
                                                                                               .rd_req_desc_0_axid_1_reg(rd_req_desc_0_axid_1_reg),
                                                                                               .rd_req_desc_0_axid_2_reg(rd_req_desc_0_axid_2_reg),
                                                                                               .rd_req_desc_0_axid_3_reg(rd_req_desc_0_axid_3_reg),
                                                                                               .rd_req_desc_0_axuser_0_reg(rd_req_desc_0_axuser_0_reg),
                                                                                               .rd_req_desc_0_axuser_1_reg(rd_req_desc_0_axuser_1_reg),
                                                                                               .rd_req_desc_0_axuser_2_reg(rd_req_desc_0_axuser_2_reg),
                                                                                               .rd_req_desc_0_axuser_3_reg(rd_req_desc_0_axuser_3_reg),
                                                                                               .rd_req_desc_0_axuser_4_reg(rd_req_desc_0_axuser_4_reg),
                                                                                               .rd_req_desc_0_axuser_5_reg(rd_req_desc_0_axuser_5_reg),
                                                                                               .rd_req_desc_0_axuser_6_reg(rd_req_desc_0_axuser_6_reg),
                                                                                               .rd_req_desc_0_axuser_7_reg(rd_req_desc_0_axuser_7_reg),
                                                                                               .rd_req_desc_0_axuser_8_reg(rd_req_desc_0_axuser_8_reg),
                                                                                               .rd_req_desc_0_axuser_9_reg(rd_req_desc_0_axuser_9_reg),
                                                                                               .rd_req_desc_0_axuser_10_reg(rd_req_desc_0_axuser_10_reg),
                                                                                               .rd_req_desc_0_axuser_11_reg(rd_req_desc_0_axuser_11_reg),
                                                                                               .rd_req_desc_0_axuser_12_reg(rd_req_desc_0_axuser_12_reg),
                                                                                               .rd_req_desc_0_axuser_13_reg(rd_req_desc_0_axuser_13_reg),
                                                                                               .rd_req_desc_0_axuser_14_reg(rd_req_desc_0_axuser_14_reg),
                                                                                               .rd_req_desc_0_axuser_15_reg(rd_req_desc_0_axuser_15_reg),
                                                                                               .rd_resp_desc_0_data_offset_reg(rd_resp_desc_0_data_offset_reg),
                                                                                               .rd_resp_desc_0_data_size_reg(rd_resp_desc_0_data_size_reg),
                                                                                               .rd_resp_desc_0_data_host_addr_0_reg(rd_resp_desc_0_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_0_data_host_addr_1_reg(rd_resp_desc_0_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_0_data_host_addr_2_reg(rd_resp_desc_0_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_0_data_host_addr_3_reg(rd_resp_desc_0_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_0_resp_reg(rd_resp_desc_0_resp_reg),
                                                                                               .rd_resp_desc_0_xid_0_reg(rd_resp_desc_0_xid_0_reg),
                                                                                               .rd_resp_desc_0_xid_1_reg(rd_resp_desc_0_xid_1_reg),
                                                                                               .rd_resp_desc_0_xid_2_reg(rd_resp_desc_0_xid_2_reg),
                                                                                               .rd_resp_desc_0_xid_3_reg(rd_resp_desc_0_xid_3_reg),
                                                                                               .rd_resp_desc_0_xuser_0_reg(rd_resp_desc_0_xuser_0_reg),
                                                                                               .rd_resp_desc_0_xuser_1_reg(rd_resp_desc_0_xuser_1_reg),
                                                                                               .rd_resp_desc_0_xuser_2_reg(rd_resp_desc_0_xuser_2_reg),
                                                                                               .rd_resp_desc_0_xuser_3_reg(rd_resp_desc_0_xuser_3_reg),
                                                                                               .rd_resp_desc_0_xuser_4_reg(rd_resp_desc_0_xuser_4_reg),
                                                                                               .rd_resp_desc_0_xuser_5_reg(rd_resp_desc_0_xuser_5_reg),
                                                                                               .rd_resp_desc_0_xuser_6_reg(rd_resp_desc_0_xuser_6_reg),
                                                                                               .rd_resp_desc_0_xuser_7_reg(rd_resp_desc_0_xuser_7_reg),
                                                                                               .rd_resp_desc_0_xuser_8_reg(rd_resp_desc_0_xuser_8_reg),
                                                                                               .rd_resp_desc_0_xuser_9_reg(rd_resp_desc_0_xuser_9_reg),
                                                                                               .rd_resp_desc_0_xuser_10_reg(rd_resp_desc_0_xuser_10_reg),
                                                                                               .rd_resp_desc_0_xuser_11_reg(rd_resp_desc_0_xuser_11_reg),
                                                                                               .rd_resp_desc_0_xuser_12_reg(rd_resp_desc_0_xuser_12_reg),
                                                                                               .rd_resp_desc_0_xuser_13_reg(rd_resp_desc_0_xuser_13_reg),
                                                                                               .rd_resp_desc_0_xuser_14_reg(rd_resp_desc_0_xuser_14_reg),
                                                                                               .rd_resp_desc_0_xuser_15_reg(rd_resp_desc_0_xuser_15_reg),
                                                                                               .wr_req_desc_0_txn_type_reg(wr_req_desc_0_txn_type_reg),
                                                                                               .wr_req_desc_0_size_reg(wr_req_desc_0_size_reg),
                                                                                               .wr_req_desc_0_data_offset_reg(wr_req_desc_0_data_offset_reg),
                                                                                               .wr_req_desc_0_data_host_addr_0_reg(wr_req_desc_0_data_host_addr_0_reg),
                                                                                               .wr_req_desc_0_data_host_addr_1_reg(wr_req_desc_0_data_host_addr_1_reg),
                                                                                               .wr_req_desc_0_data_host_addr_2_reg(wr_req_desc_0_data_host_addr_2_reg),
                                                                                               .wr_req_desc_0_data_host_addr_3_reg(wr_req_desc_0_data_host_addr_3_reg),
                                                                                               .wr_req_desc_0_wstrb_host_addr_0_reg(wr_req_desc_0_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_0_wstrb_host_addr_1_reg(wr_req_desc_0_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_0_wstrb_host_addr_2_reg(wr_req_desc_0_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_0_wstrb_host_addr_3_reg(wr_req_desc_0_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_0_axsize_reg(wr_req_desc_0_axsize_reg),
                                                                                               .wr_req_desc_0_attr_reg(wr_req_desc_0_attr_reg),
                                                                                               .wr_req_desc_0_axaddr_0_reg(wr_req_desc_0_axaddr_0_reg),
                                                                                               .wr_req_desc_0_axaddr_1_reg(wr_req_desc_0_axaddr_1_reg),
                                                                                               .wr_req_desc_0_axaddr_2_reg(wr_req_desc_0_axaddr_2_reg),
                                                                                               .wr_req_desc_0_axaddr_3_reg(wr_req_desc_0_axaddr_3_reg),
                                                                                               .wr_req_desc_0_axid_0_reg(wr_req_desc_0_axid_0_reg),
                                                                                               .wr_req_desc_0_axid_1_reg(wr_req_desc_0_axid_1_reg),
                                                                                               .wr_req_desc_0_axid_2_reg(wr_req_desc_0_axid_2_reg),
                                                                                               .wr_req_desc_0_axid_3_reg(wr_req_desc_0_axid_3_reg),
                                                                                               .wr_req_desc_0_axuser_0_reg(wr_req_desc_0_axuser_0_reg),
                                                                                               .wr_req_desc_0_axuser_1_reg(wr_req_desc_0_axuser_1_reg),
                                                                                               .wr_req_desc_0_axuser_2_reg(wr_req_desc_0_axuser_2_reg),
                                                                                               .wr_req_desc_0_axuser_3_reg(wr_req_desc_0_axuser_3_reg),
                                                                                               .wr_req_desc_0_axuser_4_reg(wr_req_desc_0_axuser_4_reg),
                                                                                               .wr_req_desc_0_axuser_5_reg(wr_req_desc_0_axuser_5_reg),
                                                                                               .wr_req_desc_0_axuser_6_reg(wr_req_desc_0_axuser_6_reg),
                                                                                               .wr_req_desc_0_axuser_7_reg(wr_req_desc_0_axuser_7_reg),
                                                                                               .wr_req_desc_0_axuser_8_reg(wr_req_desc_0_axuser_8_reg),
                                                                                               .wr_req_desc_0_axuser_9_reg(wr_req_desc_0_axuser_9_reg),
                                                                                               .wr_req_desc_0_axuser_10_reg(wr_req_desc_0_axuser_10_reg),
                                                                                               .wr_req_desc_0_axuser_11_reg(wr_req_desc_0_axuser_11_reg),
                                                                                               .wr_req_desc_0_axuser_12_reg(wr_req_desc_0_axuser_12_reg),
                                                                                               .wr_req_desc_0_axuser_13_reg(wr_req_desc_0_axuser_13_reg),
                                                                                               .wr_req_desc_0_axuser_14_reg(wr_req_desc_0_axuser_14_reg),
                                                                                               .wr_req_desc_0_axuser_15_reg(wr_req_desc_0_axuser_15_reg),
                                                                                               .wr_req_desc_0_wuser_0_reg(wr_req_desc_0_wuser_0_reg),
                                                                                               .wr_req_desc_0_wuser_1_reg(wr_req_desc_0_wuser_1_reg),
                                                                                               .wr_req_desc_0_wuser_2_reg(wr_req_desc_0_wuser_2_reg),
                                                                                               .wr_req_desc_0_wuser_3_reg(wr_req_desc_0_wuser_3_reg),
                                                                                               .wr_req_desc_0_wuser_4_reg(wr_req_desc_0_wuser_4_reg),
                                                                                               .wr_req_desc_0_wuser_5_reg(wr_req_desc_0_wuser_5_reg),
                                                                                               .wr_req_desc_0_wuser_6_reg(wr_req_desc_0_wuser_6_reg),
                                                                                               .wr_req_desc_0_wuser_7_reg(wr_req_desc_0_wuser_7_reg),
                                                                                               .wr_req_desc_0_wuser_8_reg(wr_req_desc_0_wuser_8_reg),
                                                                                               .wr_req_desc_0_wuser_9_reg(wr_req_desc_0_wuser_9_reg),
                                                                                               .wr_req_desc_0_wuser_10_reg(wr_req_desc_0_wuser_10_reg),
                                                                                               .wr_req_desc_0_wuser_11_reg(wr_req_desc_0_wuser_11_reg),
                                                                                               .wr_req_desc_0_wuser_12_reg(wr_req_desc_0_wuser_12_reg),
                                                                                               .wr_req_desc_0_wuser_13_reg(wr_req_desc_0_wuser_13_reg),
                                                                                               .wr_req_desc_0_wuser_14_reg(wr_req_desc_0_wuser_14_reg),
                                                                                               .wr_req_desc_0_wuser_15_reg(wr_req_desc_0_wuser_15_reg),
                                                                                               .wr_resp_desc_0_resp_reg(wr_resp_desc_0_resp_reg),
                                                                                               .wr_resp_desc_0_xid_0_reg(wr_resp_desc_0_xid_0_reg),
                                                                                               .wr_resp_desc_0_xid_1_reg(wr_resp_desc_0_xid_1_reg),
                                                                                               .wr_resp_desc_0_xid_2_reg(wr_resp_desc_0_xid_2_reg),
                                                                                               .wr_resp_desc_0_xid_3_reg(wr_resp_desc_0_xid_3_reg),
                                                                                               .wr_resp_desc_0_xuser_0_reg(wr_resp_desc_0_xuser_0_reg),
                                                                                               .wr_resp_desc_0_xuser_1_reg(wr_resp_desc_0_xuser_1_reg),
                                                                                               .wr_resp_desc_0_xuser_2_reg(wr_resp_desc_0_xuser_2_reg),
                                                                                               .wr_resp_desc_0_xuser_3_reg(wr_resp_desc_0_xuser_3_reg),
                                                                                               .wr_resp_desc_0_xuser_4_reg(wr_resp_desc_0_xuser_4_reg),
                                                                                               .wr_resp_desc_0_xuser_5_reg(wr_resp_desc_0_xuser_5_reg),
                                                                                               .wr_resp_desc_0_xuser_6_reg(wr_resp_desc_0_xuser_6_reg),
                                                                                               .wr_resp_desc_0_xuser_7_reg(wr_resp_desc_0_xuser_7_reg),
                                                                                               .wr_resp_desc_0_xuser_8_reg(wr_resp_desc_0_xuser_8_reg),
                                                                                               .wr_resp_desc_0_xuser_9_reg(wr_resp_desc_0_xuser_9_reg),
                                                                                               .wr_resp_desc_0_xuser_10_reg(wr_resp_desc_0_xuser_10_reg),
                                                                                               .wr_resp_desc_0_xuser_11_reg(wr_resp_desc_0_xuser_11_reg),
                                                                                               .wr_resp_desc_0_xuser_12_reg(wr_resp_desc_0_xuser_12_reg),
                                                                                               .wr_resp_desc_0_xuser_13_reg(wr_resp_desc_0_xuser_13_reg),
                                                                                               .wr_resp_desc_0_xuser_14_reg(wr_resp_desc_0_xuser_14_reg),
                                                                                               .wr_resp_desc_0_xuser_15_reg(wr_resp_desc_0_xuser_15_reg),
                                                                                               .sn_req_desc_0_attr_reg(sn_req_desc_0_attr_reg),
                                                                                               .sn_req_desc_0_acaddr_0_reg(sn_req_desc_0_acaddr_0_reg),
                                                                                               .sn_req_desc_0_acaddr_1_reg(sn_req_desc_0_acaddr_1_reg),
                                                                                               .sn_req_desc_0_acaddr_2_reg(sn_req_desc_0_acaddr_2_reg),
                                                                                               .sn_req_desc_0_acaddr_3_reg(sn_req_desc_0_acaddr_3_reg),
                                                                                               .sn_resp_desc_0_resp_reg(sn_resp_desc_0_resp_reg),
                                                                                               .rd_req_desc_1_txn_type_reg(rd_req_desc_1_txn_type_reg),
                                                                                               .rd_req_desc_1_size_reg(rd_req_desc_1_size_reg),
                                                                                               .rd_req_desc_1_axsize_reg(rd_req_desc_1_axsize_reg),
                                                                                               .rd_req_desc_1_attr_reg(rd_req_desc_1_attr_reg),
                                                                                               .rd_req_desc_1_axaddr_0_reg(rd_req_desc_1_axaddr_0_reg),
                                                                                               .rd_req_desc_1_axaddr_1_reg(rd_req_desc_1_axaddr_1_reg),
                                                                                               .rd_req_desc_1_axaddr_2_reg(rd_req_desc_1_axaddr_2_reg),
                                                                                               .rd_req_desc_1_axaddr_3_reg(rd_req_desc_1_axaddr_3_reg),
                                                                                               .rd_req_desc_1_axid_0_reg(rd_req_desc_1_axid_0_reg),
                                                                                               .rd_req_desc_1_axid_1_reg(rd_req_desc_1_axid_1_reg),
                                                                                               .rd_req_desc_1_axid_2_reg(rd_req_desc_1_axid_2_reg),
                                                                                               .rd_req_desc_1_axid_3_reg(rd_req_desc_1_axid_3_reg),
                                                                                               .rd_req_desc_1_axuser_0_reg(rd_req_desc_1_axuser_0_reg),
                                                                                               .rd_req_desc_1_axuser_1_reg(rd_req_desc_1_axuser_1_reg),
                                                                                               .rd_req_desc_1_axuser_2_reg(rd_req_desc_1_axuser_2_reg),
                                                                                               .rd_req_desc_1_axuser_3_reg(rd_req_desc_1_axuser_3_reg),
                                                                                               .rd_req_desc_1_axuser_4_reg(rd_req_desc_1_axuser_4_reg),
                                                                                               .rd_req_desc_1_axuser_5_reg(rd_req_desc_1_axuser_5_reg),
                                                                                               .rd_req_desc_1_axuser_6_reg(rd_req_desc_1_axuser_6_reg),
                                                                                               .rd_req_desc_1_axuser_7_reg(rd_req_desc_1_axuser_7_reg),
                                                                                               .rd_req_desc_1_axuser_8_reg(rd_req_desc_1_axuser_8_reg),
                                                                                               .rd_req_desc_1_axuser_9_reg(rd_req_desc_1_axuser_9_reg),
                                                                                               .rd_req_desc_1_axuser_10_reg(rd_req_desc_1_axuser_10_reg),
                                                                                               .rd_req_desc_1_axuser_11_reg(rd_req_desc_1_axuser_11_reg),
                                                                                               .rd_req_desc_1_axuser_12_reg(rd_req_desc_1_axuser_12_reg),
                                                                                               .rd_req_desc_1_axuser_13_reg(rd_req_desc_1_axuser_13_reg),
                                                                                               .rd_req_desc_1_axuser_14_reg(rd_req_desc_1_axuser_14_reg),
                                                                                               .rd_req_desc_1_axuser_15_reg(rd_req_desc_1_axuser_15_reg),
                                                                                               .rd_resp_desc_1_data_offset_reg(rd_resp_desc_1_data_offset_reg),
                                                                                               .rd_resp_desc_1_data_size_reg(rd_resp_desc_1_data_size_reg),
                                                                                               .rd_resp_desc_1_data_host_addr_0_reg(rd_resp_desc_1_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_1_data_host_addr_1_reg(rd_resp_desc_1_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_1_data_host_addr_2_reg(rd_resp_desc_1_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_1_data_host_addr_3_reg(rd_resp_desc_1_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_1_resp_reg(rd_resp_desc_1_resp_reg),
                                                                                               .rd_resp_desc_1_xid_0_reg(rd_resp_desc_1_xid_0_reg),
                                                                                               .rd_resp_desc_1_xid_1_reg(rd_resp_desc_1_xid_1_reg),
                                                                                               .rd_resp_desc_1_xid_2_reg(rd_resp_desc_1_xid_2_reg),
                                                                                               .rd_resp_desc_1_xid_3_reg(rd_resp_desc_1_xid_3_reg),
                                                                                               .rd_resp_desc_1_xuser_0_reg(rd_resp_desc_1_xuser_0_reg),
                                                                                               .rd_resp_desc_1_xuser_1_reg(rd_resp_desc_1_xuser_1_reg),
                                                                                               .rd_resp_desc_1_xuser_2_reg(rd_resp_desc_1_xuser_2_reg),
                                                                                               .rd_resp_desc_1_xuser_3_reg(rd_resp_desc_1_xuser_3_reg),
                                                                                               .rd_resp_desc_1_xuser_4_reg(rd_resp_desc_1_xuser_4_reg),
                                                                                               .rd_resp_desc_1_xuser_5_reg(rd_resp_desc_1_xuser_5_reg),
                                                                                               .rd_resp_desc_1_xuser_6_reg(rd_resp_desc_1_xuser_6_reg),
                                                                                               .rd_resp_desc_1_xuser_7_reg(rd_resp_desc_1_xuser_7_reg),
                                                                                               .rd_resp_desc_1_xuser_8_reg(rd_resp_desc_1_xuser_8_reg),
                                                                                               .rd_resp_desc_1_xuser_9_reg(rd_resp_desc_1_xuser_9_reg),
                                                                                               .rd_resp_desc_1_xuser_10_reg(rd_resp_desc_1_xuser_10_reg),
                                                                                               .rd_resp_desc_1_xuser_11_reg(rd_resp_desc_1_xuser_11_reg),
                                                                                               .rd_resp_desc_1_xuser_12_reg(rd_resp_desc_1_xuser_12_reg),
                                                                                               .rd_resp_desc_1_xuser_13_reg(rd_resp_desc_1_xuser_13_reg),
                                                                                               .rd_resp_desc_1_xuser_14_reg(rd_resp_desc_1_xuser_14_reg),
                                                                                               .rd_resp_desc_1_xuser_15_reg(rd_resp_desc_1_xuser_15_reg),
                                                                                               .wr_req_desc_1_txn_type_reg(wr_req_desc_1_txn_type_reg),
                                                                                               .wr_req_desc_1_size_reg(wr_req_desc_1_size_reg),
                                                                                               .wr_req_desc_1_data_offset_reg(wr_req_desc_1_data_offset_reg),
                                                                                               .wr_req_desc_1_data_host_addr_0_reg(wr_req_desc_1_data_host_addr_0_reg),
                                                                                               .wr_req_desc_1_data_host_addr_1_reg(wr_req_desc_1_data_host_addr_1_reg),
                                                                                               .wr_req_desc_1_data_host_addr_2_reg(wr_req_desc_1_data_host_addr_2_reg),
                                                                                               .wr_req_desc_1_data_host_addr_3_reg(wr_req_desc_1_data_host_addr_3_reg),
                                                                                               .wr_req_desc_1_wstrb_host_addr_0_reg(wr_req_desc_1_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_1_wstrb_host_addr_1_reg(wr_req_desc_1_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_1_wstrb_host_addr_2_reg(wr_req_desc_1_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_1_wstrb_host_addr_3_reg(wr_req_desc_1_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_1_axsize_reg(wr_req_desc_1_axsize_reg),
                                                                                               .wr_req_desc_1_attr_reg(wr_req_desc_1_attr_reg),
                                                                                               .wr_req_desc_1_axaddr_0_reg(wr_req_desc_1_axaddr_0_reg),
                                                                                               .wr_req_desc_1_axaddr_1_reg(wr_req_desc_1_axaddr_1_reg),
                                                                                               .wr_req_desc_1_axaddr_2_reg(wr_req_desc_1_axaddr_2_reg),
                                                                                               .wr_req_desc_1_axaddr_3_reg(wr_req_desc_1_axaddr_3_reg),
                                                                                               .wr_req_desc_1_axid_0_reg(wr_req_desc_1_axid_0_reg),
                                                                                               .wr_req_desc_1_axid_1_reg(wr_req_desc_1_axid_1_reg),
                                                                                               .wr_req_desc_1_axid_2_reg(wr_req_desc_1_axid_2_reg),
                                                                                               .wr_req_desc_1_axid_3_reg(wr_req_desc_1_axid_3_reg),
                                                                                               .wr_req_desc_1_axuser_0_reg(wr_req_desc_1_axuser_0_reg),
                                                                                               .wr_req_desc_1_axuser_1_reg(wr_req_desc_1_axuser_1_reg),
                                                                                               .wr_req_desc_1_axuser_2_reg(wr_req_desc_1_axuser_2_reg),
                                                                                               .wr_req_desc_1_axuser_3_reg(wr_req_desc_1_axuser_3_reg),
                                                                                               .wr_req_desc_1_axuser_4_reg(wr_req_desc_1_axuser_4_reg),
                                                                                               .wr_req_desc_1_axuser_5_reg(wr_req_desc_1_axuser_5_reg),
                                                                                               .wr_req_desc_1_axuser_6_reg(wr_req_desc_1_axuser_6_reg),
                                                                                               .wr_req_desc_1_axuser_7_reg(wr_req_desc_1_axuser_7_reg),
                                                                                               .wr_req_desc_1_axuser_8_reg(wr_req_desc_1_axuser_8_reg),
                                                                                               .wr_req_desc_1_axuser_9_reg(wr_req_desc_1_axuser_9_reg),
                                                                                               .wr_req_desc_1_axuser_10_reg(wr_req_desc_1_axuser_10_reg),
                                                                                               .wr_req_desc_1_axuser_11_reg(wr_req_desc_1_axuser_11_reg),
                                                                                               .wr_req_desc_1_axuser_12_reg(wr_req_desc_1_axuser_12_reg),
                                                                                               .wr_req_desc_1_axuser_13_reg(wr_req_desc_1_axuser_13_reg),
                                                                                               .wr_req_desc_1_axuser_14_reg(wr_req_desc_1_axuser_14_reg),
                                                                                               .wr_req_desc_1_axuser_15_reg(wr_req_desc_1_axuser_15_reg),
                                                                                               .wr_req_desc_1_wuser_0_reg(wr_req_desc_1_wuser_0_reg),
                                                                                               .wr_req_desc_1_wuser_1_reg(wr_req_desc_1_wuser_1_reg),
                                                                                               .wr_req_desc_1_wuser_2_reg(wr_req_desc_1_wuser_2_reg),
                                                                                               .wr_req_desc_1_wuser_3_reg(wr_req_desc_1_wuser_3_reg),
                                                                                               .wr_req_desc_1_wuser_4_reg(wr_req_desc_1_wuser_4_reg),
                                                                                               .wr_req_desc_1_wuser_5_reg(wr_req_desc_1_wuser_5_reg),
                                                                                               .wr_req_desc_1_wuser_6_reg(wr_req_desc_1_wuser_6_reg),
                                                                                               .wr_req_desc_1_wuser_7_reg(wr_req_desc_1_wuser_7_reg),
                                                                                               .wr_req_desc_1_wuser_8_reg(wr_req_desc_1_wuser_8_reg),
                                                                                               .wr_req_desc_1_wuser_9_reg(wr_req_desc_1_wuser_9_reg),
                                                                                               .wr_req_desc_1_wuser_10_reg(wr_req_desc_1_wuser_10_reg),
                                                                                               .wr_req_desc_1_wuser_11_reg(wr_req_desc_1_wuser_11_reg),
                                                                                               .wr_req_desc_1_wuser_12_reg(wr_req_desc_1_wuser_12_reg),
                                                                                               .wr_req_desc_1_wuser_13_reg(wr_req_desc_1_wuser_13_reg),
                                                                                               .wr_req_desc_1_wuser_14_reg(wr_req_desc_1_wuser_14_reg),
                                                                                               .wr_req_desc_1_wuser_15_reg(wr_req_desc_1_wuser_15_reg),
                                                                                               .wr_resp_desc_1_resp_reg(wr_resp_desc_1_resp_reg),
                                                                                               .wr_resp_desc_1_xid_0_reg(wr_resp_desc_1_xid_0_reg),
                                                                                               .wr_resp_desc_1_xid_1_reg(wr_resp_desc_1_xid_1_reg),
                                                                                               .wr_resp_desc_1_xid_2_reg(wr_resp_desc_1_xid_2_reg),
                                                                                               .wr_resp_desc_1_xid_3_reg(wr_resp_desc_1_xid_3_reg),
                                                                                               .wr_resp_desc_1_xuser_0_reg(wr_resp_desc_1_xuser_0_reg),
                                                                                               .wr_resp_desc_1_xuser_1_reg(wr_resp_desc_1_xuser_1_reg),
                                                                                               .wr_resp_desc_1_xuser_2_reg(wr_resp_desc_1_xuser_2_reg),
                                                                                               .wr_resp_desc_1_xuser_3_reg(wr_resp_desc_1_xuser_3_reg),
                                                                                               .wr_resp_desc_1_xuser_4_reg(wr_resp_desc_1_xuser_4_reg),
                                                                                               .wr_resp_desc_1_xuser_5_reg(wr_resp_desc_1_xuser_5_reg),
                                                                                               .wr_resp_desc_1_xuser_6_reg(wr_resp_desc_1_xuser_6_reg),
                                                                                               .wr_resp_desc_1_xuser_7_reg(wr_resp_desc_1_xuser_7_reg),
                                                                                               .wr_resp_desc_1_xuser_8_reg(wr_resp_desc_1_xuser_8_reg),
                                                                                               .wr_resp_desc_1_xuser_9_reg(wr_resp_desc_1_xuser_9_reg),
                                                                                               .wr_resp_desc_1_xuser_10_reg(wr_resp_desc_1_xuser_10_reg),
                                                                                               .wr_resp_desc_1_xuser_11_reg(wr_resp_desc_1_xuser_11_reg),
                                                                                               .wr_resp_desc_1_xuser_12_reg(wr_resp_desc_1_xuser_12_reg),
                                                                                               .wr_resp_desc_1_xuser_13_reg(wr_resp_desc_1_xuser_13_reg),
                                                                                               .wr_resp_desc_1_xuser_14_reg(wr_resp_desc_1_xuser_14_reg),
                                                                                               .wr_resp_desc_1_xuser_15_reg(wr_resp_desc_1_xuser_15_reg),
                                                                                               .sn_req_desc_1_attr_reg(sn_req_desc_1_attr_reg),
                                                                                               .sn_req_desc_1_acaddr_0_reg(sn_req_desc_1_acaddr_0_reg),
                                                                                               .sn_req_desc_1_acaddr_1_reg(sn_req_desc_1_acaddr_1_reg),
                                                                                               .sn_req_desc_1_acaddr_2_reg(sn_req_desc_1_acaddr_2_reg),
                                                                                               .sn_req_desc_1_acaddr_3_reg(sn_req_desc_1_acaddr_3_reg),
                                                                                               .sn_resp_desc_1_resp_reg(sn_resp_desc_1_resp_reg),
                                                                                               .rd_req_desc_2_txn_type_reg(rd_req_desc_2_txn_type_reg),
                                                                                               .rd_req_desc_2_size_reg(rd_req_desc_2_size_reg),
                                                                                               .rd_req_desc_2_axsize_reg(rd_req_desc_2_axsize_reg),
                                                                                               .rd_req_desc_2_attr_reg(rd_req_desc_2_attr_reg),
                                                                                               .rd_req_desc_2_axaddr_0_reg(rd_req_desc_2_axaddr_0_reg),
                                                                                               .rd_req_desc_2_axaddr_1_reg(rd_req_desc_2_axaddr_1_reg),
                                                                                               .rd_req_desc_2_axaddr_2_reg(rd_req_desc_2_axaddr_2_reg),
                                                                                               .rd_req_desc_2_axaddr_3_reg(rd_req_desc_2_axaddr_3_reg),
                                                                                               .rd_req_desc_2_axid_0_reg(rd_req_desc_2_axid_0_reg),
                                                                                               .rd_req_desc_2_axid_1_reg(rd_req_desc_2_axid_1_reg),
                                                                                               .rd_req_desc_2_axid_2_reg(rd_req_desc_2_axid_2_reg),
                                                                                               .rd_req_desc_2_axid_3_reg(rd_req_desc_2_axid_3_reg),
                                                                                               .rd_req_desc_2_axuser_0_reg(rd_req_desc_2_axuser_0_reg),
                                                                                               .rd_req_desc_2_axuser_1_reg(rd_req_desc_2_axuser_1_reg),
                                                                                               .rd_req_desc_2_axuser_2_reg(rd_req_desc_2_axuser_2_reg),
                                                                                               .rd_req_desc_2_axuser_3_reg(rd_req_desc_2_axuser_3_reg),
                                                                                               .rd_req_desc_2_axuser_4_reg(rd_req_desc_2_axuser_4_reg),
                                                                                               .rd_req_desc_2_axuser_5_reg(rd_req_desc_2_axuser_5_reg),
                                                                                               .rd_req_desc_2_axuser_6_reg(rd_req_desc_2_axuser_6_reg),
                                                                                               .rd_req_desc_2_axuser_7_reg(rd_req_desc_2_axuser_7_reg),
                                                                                               .rd_req_desc_2_axuser_8_reg(rd_req_desc_2_axuser_8_reg),
                                                                                               .rd_req_desc_2_axuser_9_reg(rd_req_desc_2_axuser_9_reg),
                                                                                               .rd_req_desc_2_axuser_10_reg(rd_req_desc_2_axuser_10_reg),
                                                                                               .rd_req_desc_2_axuser_11_reg(rd_req_desc_2_axuser_11_reg),
                                                                                               .rd_req_desc_2_axuser_12_reg(rd_req_desc_2_axuser_12_reg),
                                                                                               .rd_req_desc_2_axuser_13_reg(rd_req_desc_2_axuser_13_reg),
                                                                                               .rd_req_desc_2_axuser_14_reg(rd_req_desc_2_axuser_14_reg),
                                                                                               .rd_req_desc_2_axuser_15_reg(rd_req_desc_2_axuser_15_reg),
                                                                                               .rd_resp_desc_2_data_offset_reg(rd_resp_desc_2_data_offset_reg),
                                                                                               .rd_resp_desc_2_data_size_reg(rd_resp_desc_2_data_size_reg),
                                                                                               .rd_resp_desc_2_data_host_addr_0_reg(rd_resp_desc_2_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_2_data_host_addr_1_reg(rd_resp_desc_2_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_2_data_host_addr_2_reg(rd_resp_desc_2_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_2_data_host_addr_3_reg(rd_resp_desc_2_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_2_resp_reg(rd_resp_desc_2_resp_reg),
                                                                                               .rd_resp_desc_2_xid_0_reg(rd_resp_desc_2_xid_0_reg),
                                                                                               .rd_resp_desc_2_xid_1_reg(rd_resp_desc_2_xid_1_reg),
                                                                                               .rd_resp_desc_2_xid_2_reg(rd_resp_desc_2_xid_2_reg),
                                                                                               .rd_resp_desc_2_xid_3_reg(rd_resp_desc_2_xid_3_reg),
                                                                                               .rd_resp_desc_2_xuser_0_reg(rd_resp_desc_2_xuser_0_reg),
                                                                                               .rd_resp_desc_2_xuser_1_reg(rd_resp_desc_2_xuser_1_reg),
                                                                                               .rd_resp_desc_2_xuser_2_reg(rd_resp_desc_2_xuser_2_reg),
                                                                                               .rd_resp_desc_2_xuser_3_reg(rd_resp_desc_2_xuser_3_reg),
                                                                                               .rd_resp_desc_2_xuser_4_reg(rd_resp_desc_2_xuser_4_reg),
                                                                                               .rd_resp_desc_2_xuser_5_reg(rd_resp_desc_2_xuser_5_reg),
                                                                                               .rd_resp_desc_2_xuser_6_reg(rd_resp_desc_2_xuser_6_reg),
                                                                                               .rd_resp_desc_2_xuser_7_reg(rd_resp_desc_2_xuser_7_reg),
                                                                                               .rd_resp_desc_2_xuser_8_reg(rd_resp_desc_2_xuser_8_reg),
                                                                                               .rd_resp_desc_2_xuser_9_reg(rd_resp_desc_2_xuser_9_reg),
                                                                                               .rd_resp_desc_2_xuser_10_reg(rd_resp_desc_2_xuser_10_reg),
                                                                                               .rd_resp_desc_2_xuser_11_reg(rd_resp_desc_2_xuser_11_reg),
                                                                                               .rd_resp_desc_2_xuser_12_reg(rd_resp_desc_2_xuser_12_reg),
                                                                                               .rd_resp_desc_2_xuser_13_reg(rd_resp_desc_2_xuser_13_reg),
                                                                                               .rd_resp_desc_2_xuser_14_reg(rd_resp_desc_2_xuser_14_reg),
                                                                                               .rd_resp_desc_2_xuser_15_reg(rd_resp_desc_2_xuser_15_reg),
                                                                                               .wr_req_desc_2_txn_type_reg(wr_req_desc_2_txn_type_reg),
                                                                                               .wr_req_desc_2_size_reg(wr_req_desc_2_size_reg),
                                                                                               .wr_req_desc_2_data_offset_reg(wr_req_desc_2_data_offset_reg),
                                                                                               .wr_req_desc_2_data_host_addr_0_reg(wr_req_desc_2_data_host_addr_0_reg),
                                                                                               .wr_req_desc_2_data_host_addr_1_reg(wr_req_desc_2_data_host_addr_1_reg),
                                                                                               .wr_req_desc_2_data_host_addr_2_reg(wr_req_desc_2_data_host_addr_2_reg),
                                                                                               .wr_req_desc_2_data_host_addr_3_reg(wr_req_desc_2_data_host_addr_3_reg),
                                                                                               .wr_req_desc_2_wstrb_host_addr_0_reg(wr_req_desc_2_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_2_wstrb_host_addr_1_reg(wr_req_desc_2_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_2_wstrb_host_addr_2_reg(wr_req_desc_2_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_2_wstrb_host_addr_3_reg(wr_req_desc_2_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_2_axsize_reg(wr_req_desc_2_axsize_reg),
                                                                                               .wr_req_desc_2_attr_reg(wr_req_desc_2_attr_reg),
                                                                                               .wr_req_desc_2_axaddr_0_reg(wr_req_desc_2_axaddr_0_reg),
                                                                                               .wr_req_desc_2_axaddr_1_reg(wr_req_desc_2_axaddr_1_reg),
                                                                                               .wr_req_desc_2_axaddr_2_reg(wr_req_desc_2_axaddr_2_reg),
                                                                                               .wr_req_desc_2_axaddr_3_reg(wr_req_desc_2_axaddr_3_reg),
                                                                                               .wr_req_desc_2_axid_0_reg(wr_req_desc_2_axid_0_reg),
                                                                                               .wr_req_desc_2_axid_1_reg(wr_req_desc_2_axid_1_reg),
                                                                                               .wr_req_desc_2_axid_2_reg(wr_req_desc_2_axid_2_reg),
                                                                                               .wr_req_desc_2_axid_3_reg(wr_req_desc_2_axid_3_reg),
                                                                                               .wr_req_desc_2_axuser_0_reg(wr_req_desc_2_axuser_0_reg),
                                                                                               .wr_req_desc_2_axuser_1_reg(wr_req_desc_2_axuser_1_reg),
                                                                                               .wr_req_desc_2_axuser_2_reg(wr_req_desc_2_axuser_2_reg),
                                                                                               .wr_req_desc_2_axuser_3_reg(wr_req_desc_2_axuser_3_reg),
                                                                                               .wr_req_desc_2_axuser_4_reg(wr_req_desc_2_axuser_4_reg),
                                                                                               .wr_req_desc_2_axuser_5_reg(wr_req_desc_2_axuser_5_reg),
                                                                                               .wr_req_desc_2_axuser_6_reg(wr_req_desc_2_axuser_6_reg),
                                                                                               .wr_req_desc_2_axuser_7_reg(wr_req_desc_2_axuser_7_reg),
                                                                                               .wr_req_desc_2_axuser_8_reg(wr_req_desc_2_axuser_8_reg),
                                                                                               .wr_req_desc_2_axuser_9_reg(wr_req_desc_2_axuser_9_reg),
                                                                                               .wr_req_desc_2_axuser_10_reg(wr_req_desc_2_axuser_10_reg),
                                                                                               .wr_req_desc_2_axuser_11_reg(wr_req_desc_2_axuser_11_reg),
                                                                                               .wr_req_desc_2_axuser_12_reg(wr_req_desc_2_axuser_12_reg),
                                                                                               .wr_req_desc_2_axuser_13_reg(wr_req_desc_2_axuser_13_reg),
                                                                                               .wr_req_desc_2_axuser_14_reg(wr_req_desc_2_axuser_14_reg),
                                                                                               .wr_req_desc_2_axuser_15_reg(wr_req_desc_2_axuser_15_reg),
                                                                                               .wr_req_desc_2_wuser_0_reg(wr_req_desc_2_wuser_0_reg),
                                                                                               .wr_req_desc_2_wuser_1_reg(wr_req_desc_2_wuser_1_reg),
                                                                                               .wr_req_desc_2_wuser_2_reg(wr_req_desc_2_wuser_2_reg),
                                                                                               .wr_req_desc_2_wuser_3_reg(wr_req_desc_2_wuser_3_reg),
                                                                                               .wr_req_desc_2_wuser_4_reg(wr_req_desc_2_wuser_4_reg),
                                                                                               .wr_req_desc_2_wuser_5_reg(wr_req_desc_2_wuser_5_reg),
                                                                                               .wr_req_desc_2_wuser_6_reg(wr_req_desc_2_wuser_6_reg),
                                                                                               .wr_req_desc_2_wuser_7_reg(wr_req_desc_2_wuser_7_reg),
                                                                                               .wr_req_desc_2_wuser_8_reg(wr_req_desc_2_wuser_8_reg),
                                                                                               .wr_req_desc_2_wuser_9_reg(wr_req_desc_2_wuser_9_reg),
                                                                                               .wr_req_desc_2_wuser_10_reg(wr_req_desc_2_wuser_10_reg),
                                                                                               .wr_req_desc_2_wuser_11_reg(wr_req_desc_2_wuser_11_reg),
                                                                                               .wr_req_desc_2_wuser_12_reg(wr_req_desc_2_wuser_12_reg),
                                                                                               .wr_req_desc_2_wuser_13_reg(wr_req_desc_2_wuser_13_reg),
                                                                                               .wr_req_desc_2_wuser_14_reg(wr_req_desc_2_wuser_14_reg),
                                                                                               .wr_req_desc_2_wuser_15_reg(wr_req_desc_2_wuser_15_reg),
                                                                                               .wr_resp_desc_2_resp_reg(wr_resp_desc_2_resp_reg),
                                                                                               .wr_resp_desc_2_xid_0_reg(wr_resp_desc_2_xid_0_reg),
                                                                                               .wr_resp_desc_2_xid_1_reg(wr_resp_desc_2_xid_1_reg),
                                                                                               .wr_resp_desc_2_xid_2_reg(wr_resp_desc_2_xid_2_reg),
                                                                                               .wr_resp_desc_2_xid_3_reg(wr_resp_desc_2_xid_3_reg),
                                                                                               .wr_resp_desc_2_xuser_0_reg(wr_resp_desc_2_xuser_0_reg),
                                                                                               .wr_resp_desc_2_xuser_1_reg(wr_resp_desc_2_xuser_1_reg),
                                                                                               .wr_resp_desc_2_xuser_2_reg(wr_resp_desc_2_xuser_2_reg),
                                                                                               .wr_resp_desc_2_xuser_3_reg(wr_resp_desc_2_xuser_3_reg),
                                                                                               .wr_resp_desc_2_xuser_4_reg(wr_resp_desc_2_xuser_4_reg),
                                                                                               .wr_resp_desc_2_xuser_5_reg(wr_resp_desc_2_xuser_5_reg),
                                                                                               .wr_resp_desc_2_xuser_6_reg(wr_resp_desc_2_xuser_6_reg),
                                                                                               .wr_resp_desc_2_xuser_7_reg(wr_resp_desc_2_xuser_7_reg),
                                                                                               .wr_resp_desc_2_xuser_8_reg(wr_resp_desc_2_xuser_8_reg),
                                                                                               .wr_resp_desc_2_xuser_9_reg(wr_resp_desc_2_xuser_9_reg),
                                                                                               .wr_resp_desc_2_xuser_10_reg(wr_resp_desc_2_xuser_10_reg),
                                                                                               .wr_resp_desc_2_xuser_11_reg(wr_resp_desc_2_xuser_11_reg),
                                                                                               .wr_resp_desc_2_xuser_12_reg(wr_resp_desc_2_xuser_12_reg),
                                                                                               .wr_resp_desc_2_xuser_13_reg(wr_resp_desc_2_xuser_13_reg),
                                                                                               .wr_resp_desc_2_xuser_14_reg(wr_resp_desc_2_xuser_14_reg),
                                                                                               .wr_resp_desc_2_xuser_15_reg(wr_resp_desc_2_xuser_15_reg),
                                                                                               .sn_req_desc_2_attr_reg(sn_req_desc_2_attr_reg),
                                                                                               .sn_req_desc_2_acaddr_0_reg(sn_req_desc_2_acaddr_0_reg),
                                                                                               .sn_req_desc_2_acaddr_1_reg(sn_req_desc_2_acaddr_1_reg),
                                                                                               .sn_req_desc_2_acaddr_2_reg(sn_req_desc_2_acaddr_2_reg),
                                                                                               .sn_req_desc_2_acaddr_3_reg(sn_req_desc_2_acaddr_3_reg),
                                                                                               .sn_resp_desc_2_resp_reg(sn_resp_desc_2_resp_reg),
                                                                                               .rd_req_desc_3_txn_type_reg(rd_req_desc_3_txn_type_reg),
                                                                                               .rd_req_desc_3_size_reg(rd_req_desc_3_size_reg),
                                                                                               .rd_req_desc_3_axsize_reg(rd_req_desc_3_axsize_reg),
                                                                                               .rd_req_desc_3_attr_reg(rd_req_desc_3_attr_reg),
                                                                                               .rd_req_desc_3_axaddr_0_reg(rd_req_desc_3_axaddr_0_reg),
                                                                                               .rd_req_desc_3_axaddr_1_reg(rd_req_desc_3_axaddr_1_reg),
                                                                                               .rd_req_desc_3_axaddr_2_reg(rd_req_desc_3_axaddr_2_reg),
                                                                                               .rd_req_desc_3_axaddr_3_reg(rd_req_desc_3_axaddr_3_reg),
                                                                                               .rd_req_desc_3_axid_0_reg(rd_req_desc_3_axid_0_reg),
                                                                                               .rd_req_desc_3_axid_1_reg(rd_req_desc_3_axid_1_reg),
                                                                                               .rd_req_desc_3_axid_2_reg(rd_req_desc_3_axid_2_reg),
                                                                                               .rd_req_desc_3_axid_3_reg(rd_req_desc_3_axid_3_reg),
                                                                                               .rd_req_desc_3_axuser_0_reg(rd_req_desc_3_axuser_0_reg),
                                                                                               .rd_req_desc_3_axuser_1_reg(rd_req_desc_3_axuser_1_reg),
                                                                                               .rd_req_desc_3_axuser_2_reg(rd_req_desc_3_axuser_2_reg),
                                                                                               .rd_req_desc_3_axuser_3_reg(rd_req_desc_3_axuser_3_reg),
                                                                                               .rd_req_desc_3_axuser_4_reg(rd_req_desc_3_axuser_4_reg),
                                                                                               .rd_req_desc_3_axuser_5_reg(rd_req_desc_3_axuser_5_reg),
                                                                                               .rd_req_desc_3_axuser_6_reg(rd_req_desc_3_axuser_6_reg),
                                                                                               .rd_req_desc_3_axuser_7_reg(rd_req_desc_3_axuser_7_reg),
                                                                                               .rd_req_desc_3_axuser_8_reg(rd_req_desc_3_axuser_8_reg),
                                                                                               .rd_req_desc_3_axuser_9_reg(rd_req_desc_3_axuser_9_reg),
                                                                                               .rd_req_desc_3_axuser_10_reg(rd_req_desc_3_axuser_10_reg),
                                                                                               .rd_req_desc_3_axuser_11_reg(rd_req_desc_3_axuser_11_reg),
                                                                                               .rd_req_desc_3_axuser_12_reg(rd_req_desc_3_axuser_12_reg),
                                                                                               .rd_req_desc_3_axuser_13_reg(rd_req_desc_3_axuser_13_reg),
                                                                                               .rd_req_desc_3_axuser_14_reg(rd_req_desc_3_axuser_14_reg),
                                                                                               .rd_req_desc_3_axuser_15_reg(rd_req_desc_3_axuser_15_reg),
                                                                                               .rd_resp_desc_3_data_offset_reg(rd_resp_desc_3_data_offset_reg),
                                                                                               .rd_resp_desc_3_data_size_reg(rd_resp_desc_3_data_size_reg),
                                                                                               .rd_resp_desc_3_data_host_addr_0_reg(rd_resp_desc_3_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_3_data_host_addr_1_reg(rd_resp_desc_3_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_3_data_host_addr_2_reg(rd_resp_desc_3_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_3_data_host_addr_3_reg(rd_resp_desc_3_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_3_resp_reg(rd_resp_desc_3_resp_reg),
                                                                                               .rd_resp_desc_3_xid_0_reg(rd_resp_desc_3_xid_0_reg),
                                                                                               .rd_resp_desc_3_xid_1_reg(rd_resp_desc_3_xid_1_reg),
                                                                                               .rd_resp_desc_3_xid_2_reg(rd_resp_desc_3_xid_2_reg),
                                                                                               .rd_resp_desc_3_xid_3_reg(rd_resp_desc_3_xid_3_reg),
                                                                                               .rd_resp_desc_3_xuser_0_reg(rd_resp_desc_3_xuser_0_reg),
                                                                                               .rd_resp_desc_3_xuser_1_reg(rd_resp_desc_3_xuser_1_reg),
                                                                                               .rd_resp_desc_3_xuser_2_reg(rd_resp_desc_3_xuser_2_reg),
                                                                                               .rd_resp_desc_3_xuser_3_reg(rd_resp_desc_3_xuser_3_reg),
                                                                                               .rd_resp_desc_3_xuser_4_reg(rd_resp_desc_3_xuser_4_reg),
                                                                                               .rd_resp_desc_3_xuser_5_reg(rd_resp_desc_3_xuser_5_reg),
                                                                                               .rd_resp_desc_3_xuser_6_reg(rd_resp_desc_3_xuser_6_reg),
                                                                                               .rd_resp_desc_3_xuser_7_reg(rd_resp_desc_3_xuser_7_reg),
                                                                                               .rd_resp_desc_3_xuser_8_reg(rd_resp_desc_3_xuser_8_reg),
                                                                                               .rd_resp_desc_3_xuser_9_reg(rd_resp_desc_3_xuser_9_reg),
                                                                                               .rd_resp_desc_3_xuser_10_reg(rd_resp_desc_3_xuser_10_reg),
                                                                                               .rd_resp_desc_3_xuser_11_reg(rd_resp_desc_3_xuser_11_reg),
                                                                                               .rd_resp_desc_3_xuser_12_reg(rd_resp_desc_3_xuser_12_reg),
                                                                                               .rd_resp_desc_3_xuser_13_reg(rd_resp_desc_3_xuser_13_reg),
                                                                                               .rd_resp_desc_3_xuser_14_reg(rd_resp_desc_3_xuser_14_reg),
                                                                                               .rd_resp_desc_3_xuser_15_reg(rd_resp_desc_3_xuser_15_reg),
                                                                                               .wr_req_desc_3_txn_type_reg(wr_req_desc_3_txn_type_reg),
                                                                                               .wr_req_desc_3_size_reg(wr_req_desc_3_size_reg),
                                                                                               .wr_req_desc_3_data_offset_reg(wr_req_desc_3_data_offset_reg),
                                                                                               .wr_req_desc_3_data_host_addr_0_reg(wr_req_desc_3_data_host_addr_0_reg),
                                                                                               .wr_req_desc_3_data_host_addr_1_reg(wr_req_desc_3_data_host_addr_1_reg),
                                                                                               .wr_req_desc_3_data_host_addr_2_reg(wr_req_desc_3_data_host_addr_2_reg),
                                                                                               .wr_req_desc_3_data_host_addr_3_reg(wr_req_desc_3_data_host_addr_3_reg),
                                                                                               .wr_req_desc_3_wstrb_host_addr_0_reg(wr_req_desc_3_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_3_wstrb_host_addr_1_reg(wr_req_desc_3_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_3_wstrb_host_addr_2_reg(wr_req_desc_3_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_3_wstrb_host_addr_3_reg(wr_req_desc_3_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_3_axsize_reg(wr_req_desc_3_axsize_reg),
                                                                                               .wr_req_desc_3_attr_reg(wr_req_desc_3_attr_reg),
                                                                                               .wr_req_desc_3_axaddr_0_reg(wr_req_desc_3_axaddr_0_reg),
                                                                                               .wr_req_desc_3_axaddr_1_reg(wr_req_desc_3_axaddr_1_reg),
                                                                                               .wr_req_desc_3_axaddr_2_reg(wr_req_desc_3_axaddr_2_reg),
                                                                                               .wr_req_desc_3_axaddr_3_reg(wr_req_desc_3_axaddr_3_reg),
                                                                                               .wr_req_desc_3_axid_0_reg(wr_req_desc_3_axid_0_reg),
                                                                                               .wr_req_desc_3_axid_1_reg(wr_req_desc_3_axid_1_reg),
                                                                                               .wr_req_desc_3_axid_2_reg(wr_req_desc_3_axid_2_reg),
                                                                                               .wr_req_desc_3_axid_3_reg(wr_req_desc_3_axid_3_reg),
                                                                                               .wr_req_desc_3_axuser_0_reg(wr_req_desc_3_axuser_0_reg),
                                                                                               .wr_req_desc_3_axuser_1_reg(wr_req_desc_3_axuser_1_reg),
                                                                                               .wr_req_desc_3_axuser_2_reg(wr_req_desc_3_axuser_2_reg),
                                                                                               .wr_req_desc_3_axuser_3_reg(wr_req_desc_3_axuser_3_reg),
                                                                                               .wr_req_desc_3_axuser_4_reg(wr_req_desc_3_axuser_4_reg),
                                                                                               .wr_req_desc_3_axuser_5_reg(wr_req_desc_3_axuser_5_reg),
                                                                                               .wr_req_desc_3_axuser_6_reg(wr_req_desc_3_axuser_6_reg),
                                                                                               .wr_req_desc_3_axuser_7_reg(wr_req_desc_3_axuser_7_reg),
                                                                                               .wr_req_desc_3_axuser_8_reg(wr_req_desc_3_axuser_8_reg),
                                                                                               .wr_req_desc_3_axuser_9_reg(wr_req_desc_3_axuser_9_reg),
                                                                                               .wr_req_desc_3_axuser_10_reg(wr_req_desc_3_axuser_10_reg),
                                                                                               .wr_req_desc_3_axuser_11_reg(wr_req_desc_3_axuser_11_reg),
                                                                                               .wr_req_desc_3_axuser_12_reg(wr_req_desc_3_axuser_12_reg),
                                                                                               .wr_req_desc_3_axuser_13_reg(wr_req_desc_3_axuser_13_reg),
                                                                                               .wr_req_desc_3_axuser_14_reg(wr_req_desc_3_axuser_14_reg),
                                                                                               .wr_req_desc_3_axuser_15_reg(wr_req_desc_3_axuser_15_reg),
                                                                                               .wr_req_desc_3_wuser_0_reg(wr_req_desc_3_wuser_0_reg),
                                                                                               .wr_req_desc_3_wuser_1_reg(wr_req_desc_3_wuser_1_reg),
                                                                                               .wr_req_desc_3_wuser_2_reg(wr_req_desc_3_wuser_2_reg),
                                                                                               .wr_req_desc_3_wuser_3_reg(wr_req_desc_3_wuser_3_reg),
                                                                                               .wr_req_desc_3_wuser_4_reg(wr_req_desc_3_wuser_4_reg),
                                                                                               .wr_req_desc_3_wuser_5_reg(wr_req_desc_3_wuser_5_reg),
                                                                                               .wr_req_desc_3_wuser_6_reg(wr_req_desc_3_wuser_6_reg),
                                                                                               .wr_req_desc_3_wuser_7_reg(wr_req_desc_3_wuser_7_reg),
                                                                                               .wr_req_desc_3_wuser_8_reg(wr_req_desc_3_wuser_8_reg),
                                                                                               .wr_req_desc_3_wuser_9_reg(wr_req_desc_3_wuser_9_reg),
                                                                                               .wr_req_desc_3_wuser_10_reg(wr_req_desc_3_wuser_10_reg),
                                                                                               .wr_req_desc_3_wuser_11_reg(wr_req_desc_3_wuser_11_reg),
                                                                                               .wr_req_desc_3_wuser_12_reg(wr_req_desc_3_wuser_12_reg),
                                                                                               .wr_req_desc_3_wuser_13_reg(wr_req_desc_3_wuser_13_reg),
                                                                                               .wr_req_desc_3_wuser_14_reg(wr_req_desc_3_wuser_14_reg),
                                                                                               .wr_req_desc_3_wuser_15_reg(wr_req_desc_3_wuser_15_reg),
                                                                                               .wr_resp_desc_3_resp_reg(wr_resp_desc_3_resp_reg),
                                                                                               .wr_resp_desc_3_xid_0_reg(wr_resp_desc_3_xid_0_reg),
                                                                                               .wr_resp_desc_3_xid_1_reg(wr_resp_desc_3_xid_1_reg),
                                                                                               .wr_resp_desc_3_xid_2_reg(wr_resp_desc_3_xid_2_reg),
                                                                                               .wr_resp_desc_3_xid_3_reg(wr_resp_desc_3_xid_3_reg),
                                                                                               .wr_resp_desc_3_xuser_0_reg(wr_resp_desc_3_xuser_0_reg),
                                                                                               .wr_resp_desc_3_xuser_1_reg(wr_resp_desc_3_xuser_1_reg),
                                                                                               .wr_resp_desc_3_xuser_2_reg(wr_resp_desc_3_xuser_2_reg),
                                                                                               .wr_resp_desc_3_xuser_3_reg(wr_resp_desc_3_xuser_3_reg),
                                                                                               .wr_resp_desc_3_xuser_4_reg(wr_resp_desc_3_xuser_4_reg),
                                                                                               .wr_resp_desc_3_xuser_5_reg(wr_resp_desc_3_xuser_5_reg),
                                                                                               .wr_resp_desc_3_xuser_6_reg(wr_resp_desc_3_xuser_6_reg),
                                                                                               .wr_resp_desc_3_xuser_7_reg(wr_resp_desc_3_xuser_7_reg),
                                                                                               .wr_resp_desc_3_xuser_8_reg(wr_resp_desc_3_xuser_8_reg),
                                                                                               .wr_resp_desc_3_xuser_9_reg(wr_resp_desc_3_xuser_9_reg),
                                                                                               .wr_resp_desc_3_xuser_10_reg(wr_resp_desc_3_xuser_10_reg),
                                                                                               .wr_resp_desc_3_xuser_11_reg(wr_resp_desc_3_xuser_11_reg),
                                                                                               .wr_resp_desc_3_xuser_12_reg(wr_resp_desc_3_xuser_12_reg),
                                                                                               .wr_resp_desc_3_xuser_13_reg(wr_resp_desc_3_xuser_13_reg),
                                                                                               .wr_resp_desc_3_xuser_14_reg(wr_resp_desc_3_xuser_14_reg),
                                                                                               .wr_resp_desc_3_xuser_15_reg(wr_resp_desc_3_xuser_15_reg),
                                                                                               .sn_req_desc_3_attr_reg(sn_req_desc_3_attr_reg),
                                                                                               .sn_req_desc_3_acaddr_0_reg(sn_req_desc_3_acaddr_0_reg),
                                                                                               .sn_req_desc_3_acaddr_1_reg(sn_req_desc_3_acaddr_1_reg),
                                                                                               .sn_req_desc_3_acaddr_2_reg(sn_req_desc_3_acaddr_2_reg),
                                                                                               .sn_req_desc_3_acaddr_3_reg(sn_req_desc_3_acaddr_3_reg),
                                                                                               .sn_resp_desc_3_resp_reg(sn_resp_desc_3_resp_reg),
                                                                                               .rd_req_desc_4_txn_type_reg(rd_req_desc_4_txn_type_reg),
                                                                                               .rd_req_desc_4_size_reg(rd_req_desc_4_size_reg),
                                                                                               .rd_req_desc_4_axsize_reg(rd_req_desc_4_axsize_reg),
                                                                                               .rd_req_desc_4_attr_reg(rd_req_desc_4_attr_reg),
                                                                                               .rd_req_desc_4_axaddr_0_reg(rd_req_desc_4_axaddr_0_reg),
                                                                                               .rd_req_desc_4_axaddr_1_reg(rd_req_desc_4_axaddr_1_reg),
                                                                                               .rd_req_desc_4_axaddr_2_reg(rd_req_desc_4_axaddr_2_reg),
                                                                                               .rd_req_desc_4_axaddr_3_reg(rd_req_desc_4_axaddr_3_reg),
                                                                                               .rd_req_desc_4_axid_0_reg(rd_req_desc_4_axid_0_reg),
                                                                                               .rd_req_desc_4_axid_1_reg(rd_req_desc_4_axid_1_reg),
                                                                                               .rd_req_desc_4_axid_2_reg(rd_req_desc_4_axid_2_reg),
                                                                                               .rd_req_desc_4_axid_3_reg(rd_req_desc_4_axid_3_reg),
                                                                                               .rd_req_desc_4_axuser_0_reg(rd_req_desc_4_axuser_0_reg),
                                                                                               .rd_req_desc_4_axuser_1_reg(rd_req_desc_4_axuser_1_reg),
                                                                                               .rd_req_desc_4_axuser_2_reg(rd_req_desc_4_axuser_2_reg),
                                                                                               .rd_req_desc_4_axuser_3_reg(rd_req_desc_4_axuser_3_reg),
                                                                                               .rd_req_desc_4_axuser_4_reg(rd_req_desc_4_axuser_4_reg),
                                                                                               .rd_req_desc_4_axuser_5_reg(rd_req_desc_4_axuser_5_reg),
                                                                                               .rd_req_desc_4_axuser_6_reg(rd_req_desc_4_axuser_6_reg),
                                                                                               .rd_req_desc_4_axuser_7_reg(rd_req_desc_4_axuser_7_reg),
                                                                                               .rd_req_desc_4_axuser_8_reg(rd_req_desc_4_axuser_8_reg),
                                                                                               .rd_req_desc_4_axuser_9_reg(rd_req_desc_4_axuser_9_reg),
                                                                                               .rd_req_desc_4_axuser_10_reg(rd_req_desc_4_axuser_10_reg),
                                                                                               .rd_req_desc_4_axuser_11_reg(rd_req_desc_4_axuser_11_reg),
                                                                                               .rd_req_desc_4_axuser_12_reg(rd_req_desc_4_axuser_12_reg),
                                                                                               .rd_req_desc_4_axuser_13_reg(rd_req_desc_4_axuser_13_reg),
                                                                                               .rd_req_desc_4_axuser_14_reg(rd_req_desc_4_axuser_14_reg),
                                                                                               .rd_req_desc_4_axuser_15_reg(rd_req_desc_4_axuser_15_reg),
                                                                                               .rd_resp_desc_4_data_offset_reg(rd_resp_desc_4_data_offset_reg),
                                                                                               .rd_resp_desc_4_data_size_reg(rd_resp_desc_4_data_size_reg),
                                                                                               .rd_resp_desc_4_data_host_addr_0_reg(rd_resp_desc_4_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_4_data_host_addr_1_reg(rd_resp_desc_4_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_4_data_host_addr_2_reg(rd_resp_desc_4_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_4_data_host_addr_3_reg(rd_resp_desc_4_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_4_resp_reg(rd_resp_desc_4_resp_reg),
                                                                                               .rd_resp_desc_4_xid_0_reg(rd_resp_desc_4_xid_0_reg),
                                                                                               .rd_resp_desc_4_xid_1_reg(rd_resp_desc_4_xid_1_reg),
                                                                                               .rd_resp_desc_4_xid_2_reg(rd_resp_desc_4_xid_2_reg),
                                                                                               .rd_resp_desc_4_xid_3_reg(rd_resp_desc_4_xid_3_reg),
                                                                                               .rd_resp_desc_4_xuser_0_reg(rd_resp_desc_4_xuser_0_reg),
                                                                                               .rd_resp_desc_4_xuser_1_reg(rd_resp_desc_4_xuser_1_reg),
                                                                                               .rd_resp_desc_4_xuser_2_reg(rd_resp_desc_4_xuser_2_reg),
                                                                                               .rd_resp_desc_4_xuser_3_reg(rd_resp_desc_4_xuser_3_reg),
                                                                                               .rd_resp_desc_4_xuser_4_reg(rd_resp_desc_4_xuser_4_reg),
                                                                                               .rd_resp_desc_4_xuser_5_reg(rd_resp_desc_4_xuser_5_reg),
                                                                                               .rd_resp_desc_4_xuser_6_reg(rd_resp_desc_4_xuser_6_reg),
                                                                                               .rd_resp_desc_4_xuser_7_reg(rd_resp_desc_4_xuser_7_reg),
                                                                                               .rd_resp_desc_4_xuser_8_reg(rd_resp_desc_4_xuser_8_reg),
                                                                                               .rd_resp_desc_4_xuser_9_reg(rd_resp_desc_4_xuser_9_reg),
                                                                                               .rd_resp_desc_4_xuser_10_reg(rd_resp_desc_4_xuser_10_reg),
                                                                                               .rd_resp_desc_4_xuser_11_reg(rd_resp_desc_4_xuser_11_reg),
                                                                                               .rd_resp_desc_4_xuser_12_reg(rd_resp_desc_4_xuser_12_reg),
                                                                                               .rd_resp_desc_4_xuser_13_reg(rd_resp_desc_4_xuser_13_reg),
                                                                                               .rd_resp_desc_4_xuser_14_reg(rd_resp_desc_4_xuser_14_reg),
                                                                                               .rd_resp_desc_4_xuser_15_reg(rd_resp_desc_4_xuser_15_reg),
                                                                                               .wr_req_desc_4_txn_type_reg(wr_req_desc_4_txn_type_reg),
                                                                                               .wr_req_desc_4_size_reg(wr_req_desc_4_size_reg),
                                                                                               .wr_req_desc_4_data_offset_reg(wr_req_desc_4_data_offset_reg),
                                                                                               .wr_req_desc_4_data_host_addr_0_reg(wr_req_desc_4_data_host_addr_0_reg),
                                                                                               .wr_req_desc_4_data_host_addr_1_reg(wr_req_desc_4_data_host_addr_1_reg),
                                                                                               .wr_req_desc_4_data_host_addr_2_reg(wr_req_desc_4_data_host_addr_2_reg),
                                                                                               .wr_req_desc_4_data_host_addr_3_reg(wr_req_desc_4_data_host_addr_3_reg),
                                                                                               .wr_req_desc_4_wstrb_host_addr_0_reg(wr_req_desc_4_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_4_wstrb_host_addr_1_reg(wr_req_desc_4_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_4_wstrb_host_addr_2_reg(wr_req_desc_4_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_4_wstrb_host_addr_3_reg(wr_req_desc_4_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_4_axsize_reg(wr_req_desc_4_axsize_reg),
                                                                                               .wr_req_desc_4_attr_reg(wr_req_desc_4_attr_reg),
                                                                                               .wr_req_desc_4_axaddr_0_reg(wr_req_desc_4_axaddr_0_reg),
                                                                                               .wr_req_desc_4_axaddr_1_reg(wr_req_desc_4_axaddr_1_reg),
                                                                                               .wr_req_desc_4_axaddr_2_reg(wr_req_desc_4_axaddr_2_reg),
                                                                                               .wr_req_desc_4_axaddr_3_reg(wr_req_desc_4_axaddr_3_reg),
                                                                                               .wr_req_desc_4_axid_0_reg(wr_req_desc_4_axid_0_reg),
                                                                                               .wr_req_desc_4_axid_1_reg(wr_req_desc_4_axid_1_reg),
                                                                                               .wr_req_desc_4_axid_2_reg(wr_req_desc_4_axid_2_reg),
                                                                                               .wr_req_desc_4_axid_3_reg(wr_req_desc_4_axid_3_reg),
                                                                                               .wr_req_desc_4_axuser_0_reg(wr_req_desc_4_axuser_0_reg),
                                                                                               .wr_req_desc_4_axuser_1_reg(wr_req_desc_4_axuser_1_reg),
                                                                                               .wr_req_desc_4_axuser_2_reg(wr_req_desc_4_axuser_2_reg),
                                                                                               .wr_req_desc_4_axuser_3_reg(wr_req_desc_4_axuser_3_reg),
                                                                                               .wr_req_desc_4_axuser_4_reg(wr_req_desc_4_axuser_4_reg),
                                                                                               .wr_req_desc_4_axuser_5_reg(wr_req_desc_4_axuser_5_reg),
                                                                                               .wr_req_desc_4_axuser_6_reg(wr_req_desc_4_axuser_6_reg),
                                                                                               .wr_req_desc_4_axuser_7_reg(wr_req_desc_4_axuser_7_reg),
                                                                                               .wr_req_desc_4_axuser_8_reg(wr_req_desc_4_axuser_8_reg),
                                                                                               .wr_req_desc_4_axuser_9_reg(wr_req_desc_4_axuser_9_reg),
                                                                                               .wr_req_desc_4_axuser_10_reg(wr_req_desc_4_axuser_10_reg),
                                                                                               .wr_req_desc_4_axuser_11_reg(wr_req_desc_4_axuser_11_reg),
                                                                                               .wr_req_desc_4_axuser_12_reg(wr_req_desc_4_axuser_12_reg),
                                                                                               .wr_req_desc_4_axuser_13_reg(wr_req_desc_4_axuser_13_reg),
                                                                                               .wr_req_desc_4_axuser_14_reg(wr_req_desc_4_axuser_14_reg),
                                                                                               .wr_req_desc_4_axuser_15_reg(wr_req_desc_4_axuser_15_reg),
                                                                                               .wr_req_desc_4_wuser_0_reg(wr_req_desc_4_wuser_0_reg),
                                                                                               .wr_req_desc_4_wuser_1_reg(wr_req_desc_4_wuser_1_reg),
                                                                                               .wr_req_desc_4_wuser_2_reg(wr_req_desc_4_wuser_2_reg),
                                                                                               .wr_req_desc_4_wuser_3_reg(wr_req_desc_4_wuser_3_reg),
                                                                                               .wr_req_desc_4_wuser_4_reg(wr_req_desc_4_wuser_4_reg),
                                                                                               .wr_req_desc_4_wuser_5_reg(wr_req_desc_4_wuser_5_reg),
                                                                                               .wr_req_desc_4_wuser_6_reg(wr_req_desc_4_wuser_6_reg),
                                                                                               .wr_req_desc_4_wuser_7_reg(wr_req_desc_4_wuser_7_reg),
                                                                                               .wr_req_desc_4_wuser_8_reg(wr_req_desc_4_wuser_8_reg),
                                                                                               .wr_req_desc_4_wuser_9_reg(wr_req_desc_4_wuser_9_reg),
                                                                                               .wr_req_desc_4_wuser_10_reg(wr_req_desc_4_wuser_10_reg),
                                                                                               .wr_req_desc_4_wuser_11_reg(wr_req_desc_4_wuser_11_reg),
                                                                                               .wr_req_desc_4_wuser_12_reg(wr_req_desc_4_wuser_12_reg),
                                                                                               .wr_req_desc_4_wuser_13_reg(wr_req_desc_4_wuser_13_reg),
                                                                                               .wr_req_desc_4_wuser_14_reg(wr_req_desc_4_wuser_14_reg),
                                                                                               .wr_req_desc_4_wuser_15_reg(wr_req_desc_4_wuser_15_reg),
                                                                                               .wr_resp_desc_4_resp_reg(wr_resp_desc_4_resp_reg),
                                                                                               .wr_resp_desc_4_xid_0_reg(wr_resp_desc_4_xid_0_reg),
                                                                                               .wr_resp_desc_4_xid_1_reg(wr_resp_desc_4_xid_1_reg),
                                                                                               .wr_resp_desc_4_xid_2_reg(wr_resp_desc_4_xid_2_reg),
                                                                                               .wr_resp_desc_4_xid_3_reg(wr_resp_desc_4_xid_3_reg),
                                                                                               .wr_resp_desc_4_xuser_0_reg(wr_resp_desc_4_xuser_0_reg),
                                                                                               .wr_resp_desc_4_xuser_1_reg(wr_resp_desc_4_xuser_1_reg),
                                                                                               .wr_resp_desc_4_xuser_2_reg(wr_resp_desc_4_xuser_2_reg),
                                                                                               .wr_resp_desc_4_xuser_3_reg(wr_resp_desc_4_xuser_3_reg),
                                                                                               .wr_resp_desc_4_xuser_4_reg(wr_resp_desc_4_xuser_4_reg),
                                                                                               .wr_resp_desc_4_xuser_5_reg(wr_resp_desc_4_xuser_5_reg),
                                                                                               .wr_resp_desc_4_xuser_6_reg(wr_resp_desc_4_xuser_6_reg),
                                                                                               .wr_resp_desc_4_xuser_7_reg(wr_resp_desc_4_xuser_7_reg),
                                                                                               .wr_resp_desc_4_xuser_8_reg(wr_resp_desc_4_xuser_8_reg),
                                                                                               .wr_resp_desc_4_xuser_9_reg(wr_resp_desc_4_xuser_9_reg),
                                                                                               .wr_resp_desc_4_xuser_10_reg(wr_resp_desc_4_xuser_10_reg),
                                                                                               .wr_resp_desc_4_xuser_11_reg(wr_resp_desc_4_xuser_11_reg),
                                                                                               .wr_resp_desc_4_xuser_12_reg(wr_resp_desc_4_xuser_12_reg),
                                                                                               .wr_resp_desc_4_xuser_13_reg(wr_resp_desc_4_xuser_13_reg),
                                                                                               .wr_resp_desc_4_xuser_14_reg(wr_resp_desc_4_xuser_14_reg),
                                                                                               .wr_resp_desc_4_xuser_15_reg(wr_resp_desc_4_xuser_15_reg),
                                                                                               .sn_req_desc_4_attr_reg(sn_req_desc_4_attr_reg),
                                                                                               .sn_req_desc_4_acaddr_0_reg(sn_req_desc_4_acaddr_0_reg),
                                                                                               .sn_req_desc_4_acaddr_1_reg(sn_req_desc_4_acaddr_1_reg),
                                                                                               .sn_req_desc_4_acaddr_2_reg(sn_req_desc_4_acaddr_2_reg),
                                                                                               .sn_req_desc_4_acaddr_3_reg(sn_req_desc_4_acaddr_3_reg),
                                                                                               .sn_resp_desc_4_resp_reg(sn_resp_desc_4_resp_reg),
                                                                                               .rd_req_desc_5_txn_type_reg(rd_req_desc_5_txn_type_reg),
                                                                                               .rd_req_desc_5_size_reg(rd_req_desc_5_size_reg),
                                                                                               .rd_req_desc_5_axsize_reg(rd_req_desc_5_axsize_reg),
                                                                                               .rd_req_desc_5_attr_reg(rd_req_desc_5_attr_reg),
                                                                                               .rd_req_desc_5_axaddr_0_reg(rd_req_desc_5_axaddr_0_reg),
                                                                                               .rd_req_desc_5_axaddr_1_reg(rd_req_desc_5_axaddr_1_reg),
                                                                                               .rd_req_desc_5_axaddr_2_reg(rd_req_desc_5_axaddr_2_reg),
                                                                                               .rd_req_desc_5_axaddr_3_reg(rd_req_desc_5_axaddr_3_reg),
                                                                                               .rd_req_desc_5_axid_0_reg(rd_req_desc_5_axid_0_reg),
                                                                                               .rd_req_desc_5_axid_1_reg(rd_req_desc_5_axid_1_reg),
                                                                                               .rd_req_desc_5_axid_2_reg(rd_req_desc_5_axid_2_reg),
                                                                                               .rd_req_desc_5_axid_3_reg(rd_req_desc_5_axid_3_reg),
                                                                                               .rd_req_desc_5_axuser_0_reg(rd_req_desc_5_axuser_0_reg),
                                                                                               .rd_req_desc_5_axuser_1_reg(rd_req_desc_5_axuser_1_reg),
                                                                                               .rd_req_desc_5_axuser_2_reg(rd_req_desc_5_axuser_2_reg),
                                                                                               .rd_req_desc_5_axuser_3_reg(rd_req_desc_5_axuser_3_reg),
                                                                                               .rd_req_desc_5_axuser_4_reg(rd_req_desc_5_axuser_4_reg),
                                                                                               .rd_req_desc_5_axuser_5_reg(rd_req_desc_5_axuser_5_reg),
                                                                                               .rd_req_desc_5_axuser_6_reg(rd_req_desc_5_axuser_6_reg),
                                                                                               .rd_req_desc_5_axuser_7_reg(rd_req_desc_5_axuser_7_reg),
                                                                                               .rd_req_desc_5_axuser_8_reg(rd_req_desc_5_axuser_8_reg),
                                                                                               .rd_req_desc_5_axuser_9_reg(rd_req_desc_5_axuser_9_reg),
                                                                                               .rd_req_desc_5_axuser_10_reg(rd_req_desc_5_axuser_10_reg),
                                                                                               .rd_req_desc_5_axuser_11_reg(rd_req_desc_5_axuser_11_reg),
                                                                                               .rd_req_desc_5_axuser_12_reg(rd_req_desc_5_axuser_12_reg),
                                                                                               .rd_req_desc_5_axuser_13_reg(rd_req_desc_5_axuser_13_reg),
                                                                                               .rd_req_desc_5_axuser_14_reg(rd_req_desc_5_axuser_14_reg),
                                                                                               .rd_req_desc_5_axuser_15_reg(rd_req_desc_5_axuser_15_reg),
                                                                                               .rd_resp_desc_5_data_offset_reg(rd_resp_desc_5_data_offset_reg),
                                                                                               .rd_resp_desc_5_data_size_reg(rd_resp_desc_5_data_size_reg),
                                                                                               .rd_resp_desc_5_data_host_addr_0_reg(rd_resp_desc_5_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_5_data_host_addr_1_reg(rd_resp_desc_5_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_5_data_host_addr_2_reg(rd_resp_desc_5_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_5_data_host_addr_3_reg(rd_resp_desc_5_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_5_resp_reg(rd_resp_desc_5_resp_reg),
                                                                                               .rd_resp_desc_5_xid_0_reg(rd_resp_desc_5_xid_0_reg),
                                                                                               .rd_resp_desc_5_xid_1_reg(rd_resp_desc_5_xid_1_reg),
                                                                                               .rd_resp_desc_5_xid_2_reg(rd_resp_desc_5_xid_2_reg),
                                                                                               .rd_resp_desc_5_xid_3_reg(rd_resp_desc_5_xid_3_reg),
                                                                                               .rd_resp_desc_5_xuser_0_reg(rd_resp_desc_5_xuser_0_reg),
                                                                                               .rd_resp_desc_5_xuser_1_reg(rd_resp_desc_5_xuser_1_reg),
                                                                                               .rd_resp_desc_5_xuser_2_reg(rd_resp_desc_5_xuser_2_reg),
                                                                                               .rd_resp_desc_5_xuser_3_reg(rd_resp_desc_5_xuser_3_reg),
                                                                                               .rd_resp_desc_5_xuser_4_reg(rd_resp_desc_5_xuser_4_reg),
                                                                                               .rd_resp_desc_5_xuser_5_reg(rd_resp_desc_5_xuser_5_reg),
                                                                                               .rd_resp_desc_5_xuser_6_reg(rd_resp_desc_5_xuser_6_reg),
                                                                                               .rd_resp_desc_5_xuser_7_reg(rd_resp_desc_5_xuser_7_reg),
                                                                                               .rd_resp_desc_5_xuser_8_reg(rd_resp_desc_5_xuser_8_reg),
                                                                                               .rd_resp_desc_5_xuser_9_reg(rd_resp_desc_5_xuser_9_reg),
                                                                                               .rd_resp_desc_5_xuser_10_reg(rd_resp_desc_5_xuser_10_reg),
                                                                                               .rd_resp_desc_5_xuser_11_reg(rd_resp_desc_5_xuser_11_reg),
                                                                                               .rd_resp_desc_5_xuser_12_reg(rd_resp_desc_5_xuser_12_reg),
                                                                                               .rd_resp_desc_5_xuser_13_reg(rd_resp_desc_5_xuser_13_reg),
                                                                                               .rd_resp_desc_5_xuser_14_reg(rd_resp_desc_5_xuser_14_reg),
                                                                                               .rd_resp_desc_5_xuser_15_reg(rd_resp_desc_5_xuser_15_reg),
                                                                                               .wr_req_desc_5_txn_type_reg(wr_req_desc_5_txn_type_reg),
                                                                                               .wr_req_desc_5_size_reg(wr_req_desc_5_size_reg),
                                                                                               .wr_req_desc_5_data_offset_reg(wr_req_desc_5_data_offset_reg),
                                                                                               .wr_req_desc_5_data_host_addr_0_reg(wr_req_desc_5_data_host_addr_0_reg),
                                                                                               .wr_req_desc_5_data_host_addr_1_reg(wr_req_desc_5_data_host_addr_1_reg),
                                                                                               .wr_req_desc_5_data_host_addr_2_reg(wr_req_desc_5_data_host_addr_2_reg),
                                                                                               .wr_req_desc_5_data_host_addr_3_reg(wr_req_desc_5_data_host_addr_3_reg),
                                                                                               .wr_req_desc_5_wstrb_host_addr_0_reg(wr_req_desc_5_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_5_wstrb_host_addr_1_reg(wr_req_desc_5_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_5_wstrb_host_addr_2_reg(wr_req_desc_5_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_5_wstrb_host_addr_3_reg(wr_req_desc_5_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_5_axsize_reg(wr_req_desc_5_axsize_reg),
                                                                                               .wr_req_desc_5_attr_reg(wr_req_desc_5_attr_reg),
                                                                                               .wr_req_desc_5_axaddr_0_reg(wr_req_desc_5_axaddr_0_reg),
                                                                                               .wr_req_desc_5_axaddr_1_reg(wr_req_desc_5_axaddr_1_reg),
                                                                                               .wr_req_desc_5_axaddr_2_reg(wr_req_desc_5_axaddr_2_reg),
                                                                                               .wr_req_desc_5_axaddr_3_reg(wr_req_desc_5_axaddr_3_reg),
                                                                                               .wr_req_desc_5_axid_0_reg(wr_req_desc_5_axid_0_reg),
                                                                                               .wr_req_desc_5_axid_1_reg(wr_req_desc_5_axid_1_reg),
                                                                                               .wr_req_desc_5_axid_2_reg(wr_req_desc_5_axid_2_reg),
                                                                                               .wr_req_desc_5_axid_3_reg(wr_req_desc_5_axid_3_reg),
                                                                                               .wr_req_desc_5_axuser_0_reg(wr_req_desc_5_axuser_0_reg),
                                                                                               .wr_req_desc_5_axuser_1_reg(wr_req_desc_5_axuser_1_reg),
                                                                                               .wr_req_desc_5_axuser_2_reg(wr_req_desc_5_axuser_2_reg),
                                                                                               .wr_req_desc_5_axuser_3_reg(wr_req_desc_5_axuser_3_reg),
                                                                                               .wr_req_desc_5_axuser_4_reg(wr_req_desc_5_axuser_4_reg),
                                                                                               .wr_req_desc_5_axuser_5_reg(wr_req_desc_5_axuser_5_reg),
                                                                                               .wr_req_desc_5_axuser_6_reg(wr_req_desc_5_axuser_6_reg),
                                                                                               .wr_req_desc_5_axuser_7_reg(wr_req_desc_5_axuser_7_reg),
                                                                                               .wr_req_desc_5_axuser_8_reg(wr_req_desc_5_axuser_8_reg),
                                                                                               .wr_req_desc_5_axuser_9_reg(wr_req_desc_5_axuser_9_reg),
                                                                                               .wr_req_desc_5_axuser_10_reg(wr_req_desc_5_axuser_10_reg),
                                                                                               .wr_req_desc_5_axuser_11_reg(wr_req_desc_5_axuser_11_reg),
                                                                                               .wr_req_desc_5_axuser_12_reg(wr_req_desc_5_axuser_12_reg),
                                                                                               .wr_req_desc_5_axuser_13_reg(wr_req_desc_5_axuser_13_reg),
                                                                                               .wr_req_desc_5_axuser_14_reg(wr_req_desc_5_axuser_14_reg),
                                                                                               .wr_req_desc_5_axuser_15_reg(wr_req_desc_5_axuser_15_reg),
                                                                                               .wr_req_desc_5_wuser_0_reg(wr_req_desc_5_wuser_0_reg),
                                                                                               .wr_req_desc_5_wuser_1_reg(wr_req_desc_5_wuser_1_reg),
                                                                                               .wr_req_desc_5_wuser_2_reg(wr_req_desc_5_wuser_2_reg),
                                                                                               .wr_req_desc_5_wuser_3_reg(wr_req_desc_5_wuser_3_reg),
                                                                                               .wr_req_desc_5_wuser_4_reg(wr_req_desc_5_wuser_4_reg),
                                                                                               .wr_req_desc_5_wuser_5_reg(wr_req_desc_5_wuser_5_reg),
                                                                                               .wr_req_desc_5_wuser_6_reg(wr_req_desc_5_wuser_6_reg),
                                                                                               .wr_req_desc_5_wuser_7_reg(wr_req_desc_5_wuser_7_reg),
                                                                                               .wr_req_desc_5_wuser_8_reg(wr_req_desc_5_wuser_8_reg),
                                                                                               .wr_req_desc_5_wuser_9_reg(wr_req_desc_5_wuser_9_reg),
                                                                                               .wr_req_desc_5_wuser_10_reg(wr_req_desc_5_wuser_10_reg),
                                                                                               .wr_req_desc_5_wuser_11_reg(wr_req_desc_5_wuser_11_reg),
                                                                                               .wr_req_desc_5_wuser_12_reg(wr_req_desc_5_wuser_12_reg),
                                                                                               .wr_req_desc_5_wuser_13_reg(wr_req_desc_5_wuser_13_reg),
                                                                                               .wr_req_desc_5_wuser_14_reg(wr_req_desc_5_wuser_14_reg),
                                                                                               .wr_req_desc_5_wuser_15_reg(wr_req_desc_5_wuser_15_reg),
                                                                                               .wr_resp_desc_5_resp_reg(wr_resp_desc_5_resp_reg),
                                                                                               .wr_resp_desc_5_xid_0_reg(wr_resp_desc_5_xid_0_reg),
                                                                                               .wr_resp_desc_5_xid_1_reg(wr_resp_desc_5_xid_1_reg),
                                                                                               .wr_resp_desc_5_xid_2_reg(wr_resp_desc_5_xid_2_reg),
                                                                                               .wr_resp_desc_5_xid_3_reg(wr_resp_desc_5_xid_3_reg),
                                                                                               .wr_resp_desc_5_xuser_0_reg(wr_resp_desc_5_xuser_0_reg),
                                                                                               .wr_resp_desc_5_xuser_1_reg(wr_resp_desc_5_xuser_1_reg),
                                                                                               .wr_resp_desc_5_xuser_2_reg(wr_resp_desc_5_xuser_2_reg),
                                                                                               .wr_resp_desc_5_xuser_3_reg(wr_resp_desc_5_xuser_3_reg),
                                                                                               .wr_resp_desc_5_xuser_4_reg(wr_resp_desc_5_xuser_4_reg),
                                                                                               .wr_resp_desc_5_xuser_5_reg(wr_resp_desc_5_xuser_5_reg),
                                                                                               .wr_resp_desc_5_xuser_6_reg(wr_resp_desc_5_xuser_6_reg),
                                                                                               .wr_resp_desc_5_xuser_7_reg(wr_resp_desc_5_xuser_7_reg),
                                                                                               .wr_resp_desc_5_xuser_8_reg(wr_resp_desc_5_xuser_8_reg),
                                                                                               .wr_resp_desc_5_xuser_9_reg(wr_resp_desc_5_xuser_9_reg),
                                                                                               .wr_resp_desc_5_xuser_10_reg(wr_resp_desc_5_xuser_10_reg),
                                                                                               .wr_resp_desc_5_xuser_11_reg(wr_resp_desc_5_xuser_11_reg),
                                                                                               .wr_resp_desc_5_xuser_12_reg(wr_resp_desc_5_xuser_12_reg),
                                                                                               .wr_resp_desc_5_xuser_13_reg(wr_resp_desc_5_xuser_13_reg),
                                                                                               .wr_resp_desc_5_xuser_14_reg(wr_resp_desc_5_xuser_14_reg),
                                                                                               .wr_resp_desc_5_xuser_15_reg(wr_resp_desc_5_xuser_15_reg),
                                                                                               .sn_req_desc_5_attr_reg(sn_req_desc_5_attr_reg),
                                                                                               .sn_req_desc_5_acaddr_0_reg(sn_req_desc_5_acaddr_0_reg),
                                                                                               .sn_req_desc_5_acaddr_1_reg(sn_req_desc_5_acaddr_1_reg),
                                                                                               .sn_req_desc_5_acaddr_2_reg(sn_req_desc_5_acaddr_2_reg),
                                                                                               .sn_req_desc_5_acaddr_3_reg(sn_req_desc_5_acaddr_3_reg),
                                                                                               .sn_resp_desc_5_resp_reg(sn_resp_desc_5_resp_reg),
                                                                                               .rd_req_desc_6_txn_type_reg(rd_req_desc_6_txn_type_reg),
                                                                                               .rd_req_desc_6_size_reg(rd_req_desc_6_size_reg),
                                                                                               .rd_req_desc_6_axsize_reg(rd_req_desc_6_axsize_reg),
                                                                                               .rd_req_desc_6_attr_reg(rd_req_desc_6_attr_reg),
                                                                                               .rd_req_desc_6_axaddr_0_reg(rd_req_desc_6_axaddr_0_reg),
                                                                                               .rd_req_desc_6_axaddr_1_reg(rd_req_desc_6_axaddr_1_reg),
                                                                                               .rd_req_desc_6_axaddr_2_reg(rd_req_desc_6_axaddr_2_reg),
                                                                                               .rd_req_desc_6_axaddr_3_reg(rd_req_desc_6_axaddr_3_reg),
                                                                                               .rd_req_desc_6_axid_0_reg(rd_req_desc_6_axid_0_reg),
                                                                                               .rd_req_desc_6_axid_1_reg(rd_req_desc_6_axid_1_reg),
                                                                                               .rd_req_desc_6_axid_2_reg(rd_req_desc_6_axid_2_reg),
                                                                                               .rd_req_desc_6_axid_3_reg(rd_req_desc_6_axid_3_reg),
                                                                                               .rd_req_desc_6_axuser_0_reg(rd_req_desc_6_axuser_0_reg),
                                                                                               .rd_req_desc_6_axuser_1_reg(rd_req_desc_6_axuser_1_reg),
                                                                                               .rd_req_desc_6_axuser_2_reg(rd_req_desc_6_axuser_2_reg),
                                                                                               .rd_req_desc_6_axuser_3_reg(rd_req_desc_6_axuser_3_reg),
                                                                                               .rd_req_desc_6_axuser_4_reg(rd_req_desc_6_axuser_4_reg),
                                                                                               .rd_req_desc_6_axuser_5_reg(rd_req_desc_6_axuser_5_reg),
                                                                                               .rd_req_desc_6_axuser_6_reg(rd_req_desc_6_axuser_6_reg),
                                                                                               .rd_req_desc_6_axuser_7_reg(rd_req_desc_6_axuser_7_reg),
                                                                                               .rd_req_desc_6_axuser_8_reg(rd_req_desc_6_axuser_8_reg),
                                                                                               .rd_req_desc_6_axuser_9_reg(rd_req_desc_6_axuser_9_reg),
                                                                                               .rd_req_desc_6_axuser_10_reg(rd_req_desc_6_axuser_10_reg),
                                                                                               .rd_req_desc_6_axuser_11_reg(rd_req_desc_6_axuser_11_reg),
                                                                                               .rd_req_desc_6_axuser_12_reg(rd_req_desc_6_axuser_12_reg),
                                                                                               .rd_req_desc_6_axuser_13_reg(rd_req_desc_6_axuser_13_reg),
                                                                                               .rd_req_desc_6_axuser_14_reg(rd_req_desc_6_axuser_14_reg),
                                                                                               .rd_req_desc_6_axuser_15_reg(rd_req_desc_6_axuser_15_reg),
                                                                                               .rd_resp_desc_6_data_offset_reg(rd_resp_desc_6_data_offset_reg),
                                                                                               .rd_resp_desc_6_data_size_reg(rd_resp_desc_6_data_size_reg),
                                                                                               .rd_resp_desc_6_data_host_addr_0_reg(rd_resp_desc_6_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_6_data_host_addr_1_reg(rd_resp_desc_6_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_6_data_host_addr_2_reg(rd_resp_desc_6_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_6_data_host_addr_3_reg(rd_resp_desc_6_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_6_resp_reg(rd_resp_desc_6_resp_reg),
                                                                                               .rd_resp_desc_6_xid_0_reg(rd_resp_desc_6_xid_0_reg),
                                                                                               .rd_resp_desc_6_xid_1_reg(rd_resp_desc_6_xid_1_reg),
                                                                                               .rd_resp_desc_6_xid_2_reg(rd_resp_desc_6_xid_2_reg),
                                                                                               .rd_resp_desc_6_xid_3_reg(rd_resp_desc_6_xid_3_reg),
                                                                                               .rd_resp_desc_6_xuser_0_reg(rd_resp_desc_6_xuser_0_reg),
                                                                                               .rd_resp_desc_6_xuser_1_reg(rd_resp_desc_6_xuser_1_reg),
                                                                                               .rd_resp_desc_6_xuser_2_reg(rd_resp_desc_6_xuser_2_reg),
                                                                                               .rd_resp_desc_6_xuser_3_reg(rd_resp_desc_6_xuser_3_reg),
                                                                                               .rd_resp_desc_6_xuser_4_reg(rd_resp_desc_6_xuser_4_reg),
                                                                                               .rd_resp_desc_6_xuser_5_reg(rd_resp_desc_6_xuser_5_reg),
                                                                                               .rd_resp_desc_6_xuser_6_reg(rd_resp_desc_6_xuser_6_reg),
                                                                                               .rd_resp_desc_6_xuser_7_reg(rd_resp_desc_6_xuser_7_reg),
                                                                                               .rd_resp_desc_6_xuser_8_reg(rd_resp_desc_6_xuser_8_reg),
                                                                                               .rd_resp_desc_6_xuser_9_reg(rd_resp_desc_6_xuser_9_reg),
                                                                                               .rd_resp_desc_6_xuser_10_reg(rd_resp_desc_6_xuser_10_reg),
                                                                                               .rd_resp_desc_6_xuser_11_reg(rd_resp_desc_6_xuser_11_reg),
                                                                                               .rd_resp_desc_6_xuser_12_reg(rd_resp_desc_6_xuser_12_reg),
                                                                                               .rd_resp_desc_6_xuser_13_reg(rd_resp_desc_6_xuser_13_reg),
                                                                                               .rd_resp_desc_6_xuser_14_reg(rd_resp_desc_6_xuser_14_reg),
                                                                                               .rd_resp_desc_6_xuser_15_reg(rd_resp_desc_6_xuser_15_reg),
                                                                                               .wr_req_desc_6_txn_type_reg(wr_req_desc_6_txn_type_reg),
                                                                                               .wr_req_desc_6_size_reg(wr_req_desc_6_size_reg),
                                                                                               .wr_req_desc_6_data_offset_reg(wr_req_desc_6_data_offset_reg),
                                                                                               .wr_req_desc_6_data_host_addr_0_reg(wr_req_desc_6_data_host_addr_0_reg),
                                                                                               .wr_req_desc_6_data_host_addr_1_reg(wr_req_desc_6_data_host_addr_1_reg),
                                                                                               .wr_req_desc_6_data_host_addr_2_reg(wr_req_desc_6_data_host_addr_2_reg),
                                                                                               .wr_req_desc_6_data_host_addr_3_reg(wr_req_desc_6_data_host_addr_3_reg),
                                                                                               .wr_req_desc_6_wstrb_host_addr_0_reg(wr_req_desc_6_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_6_wstrb_host_addr_1_reg(wr_req_desc_6_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_6_wstrb_host_addr_2_reg(wr_req_desc_6_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_6_wstrb_host_addr_3_reg(wr_req_desc_6_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_6_axsize_reg(wr_req_desc_6_axsize_reg),
                                                                                               .wr_req_desc_6_attr_reg(wr_req_desc_6_attr_reg),
                                                                                               .wr_req_desc_6_axaddr_0_reg(wr_req_desc_6_axaddr_0_reg),
                                                                                               .wr_req_desc_6_axaddr_1_reg(wr_req_desc_6_axaddr_1_reg),
                                                                                               .wr_req_desc_6_axaddr_2_reg(wr_req_desc_6_axaddr_2_reg),
                                                                                               .wr_req_desc_6_axaddr_3_reg(wr_req_desc_6_axaddr_3_reg),
                                                                                               .wr_req_desc_6_axid_0_reg(wr_req_desc_6_axid_0_reg),
                                                                                               .wr_req_desc_6_axid_1_reg(wr_req_desc_6_axid_1_reg),
                                                                                               .wr_req_desc_6_axid_2_reg(wr_req_desc_6_axid_2_reg),
                                                                                               .wr_req_desc_6_axid_3_reg(wr_req_desc_6_axid_3_reg),
                                                                                               .wr_req_desc_6_axuser_0_reg(wr_req_desc_6_axuser_0_reg),
                                                                                               .wr_req_desc_6_axuser_1_reg(wr_req_desc_6_axuser_1_reg),
                                                                                               .wr_req_desc_6_axuser_2_reg(wr_req_desc_6_axuser_2_reg),
                                                                                               .wr_req_desc_6_axuser_3_reg(wr_req_desc_6_axuser_3_reg),
                                                                                               .wr_req_desc_6_axuser_4_reg(wr_req_desc_6_axuser_4_reg),
                                                                                               .wr_req_desc_6_axuser_5_reg(wr_req_desc_6_axuser_5_reg),
                                                                                               .wr_req_desc_6_axuser_6_reg(wr_req_desc_6_axuser_6_reg),
                                                                                               .wr_req_desc_6_axuser_7_reg(wr_req_desc_6_axuser_7_reg),
                                                                                               .wr_req_desc_6_axuser_8_reg(wr_req_desc_6_axuser_8_reg),
                                                                                               .wr_req_desc_6_axuser_9_reg(wr_req_desc_6_axuser_9_reg),
                                                                                               .wr_req_desc_6_axuser_10_reg(wr_req_desc_6_axuser_10_reg),
                                                                                               .wr_req_desc_6_axuser_11_reg(wr_req_desc_6_axuser_11_reg),
                                                                                               .wr_req_desc_6_axuser_12_reg(wr_req_desc_6_axuser_12_reg),
                                                                                               .wr_req_desc_6_axuser_13_reg(wr_req_desc_6_axuser_13_reg),
                                                                                               .wr_req_desc_6_axuser_14_reg(wr_req_desc_6_axuser_14_reg),
                                                                                               .wr_req_desc_6_axuser_15_reg(wr_req_desc_6_axuser_15_reg),
                                                                                               .wr_req_desc_6_wuser_0_reg(wr_req_desc_6_wuser_0_reg),
                                                                                               .wr_req_desc_6_wuser_1_reg(wr_req_desc_6_wuser_1_reg),
                                                                                               .wr_req_desc_6_wuser_2_reg(wr_req_desc_6_wuser_2_reg),
                                                                                               .wr_req_desc_6_wuser_3_reg(wr_req_desc_6_wuser_3_reg),
                                                                                               .wr_req_desc_6_wuser_4_reg(wr_req_desc_6_wuser_4_reg),
                                                                                               .wr_req_desc_6_wuser_5_reg(wr_req_desc_6_wuser_5_reg),
                                                                                               .wr_req_desc_6_wuser_6_reg(wr_req_desc_6_wuser_6_reg),
                                                                                               .wr_req_desc_6_wuser_7_reg(wr_req_desc_6_wuser_7_reg),
                                                                                               .wr_req_desc_6_wuser_8_reg(wr_req_desc_6_wuser_8_reg),
                                                                                               .wr_req_desc_6_wuser_9_reg(wr_req_desc_6_wuser_9_reg),
                                                                                               .wr_req_desc_6_wuser_10_reg(wr_req_desc_6_wuser_10_reg),
                                                                                               .wr_req_desc_6_wuser_11_reg(wr_req_desc_6_wuser_11_reg),
                                                                                               .wr_req_desc_6_wuser_12_reg(wr_req_desc_6_wuser_12_reg),
                                                                                               .wr_req_desc_6_wuser_13_reg(wr_req_desc_6_wuser_13_reg),
                                                                                               .wr_req_desc_6_wuser_14_reg(wr_req_desc_6_wuser_14_reg),
                                                                                               .wr_req_desc_6_wuser_15_reg(wr_req_desc_6_wuser_15_reg),
                                                                                               .wr_resp_desc_6_resp_reg(wr_resp_desc_6_resp_reg),
                                                                                               .wr_resp_desc_6_xid_0_reg(wr_resp_desc_6_xid_0_reg),
                                                                                               .wr_resp_desc_6_xid_1_reg(wr_resp_desc_6_xid_1_reg),
                                                                                               .wr_resp_desc_6_xid_2_reg(wr_resp_desc_6_xid_2_reg),
                                                                                               .wr_resp_desc_6_xid_3_reg(wr_resp_desc_6_xid_3_reg),
                                                                                               .wr_resp_desc_6_xuser_0_reg(wr_resp_desc_6_xuser_0_reg),
                                                                                               .wr_resp_desc_6_xuser_1_reg(wr_resp_desc_6_xuser_1_reg),
                                                                                               .wr_resp_desc_6_xuser_2_reg(wr_resp_desc_6_xuser_2_reg),
                                                                                               .wr_resp_desc_6_xuser_3_reg(wr_resp_desc_6_xuser_3_reg),
                                                                                               .wr_resp_desc_6_xuser_4_reg(wr_resp_desc_6_xuser_4_reg),
                                                                                               .wr_resp_desc_6_xuser_5_reg(wr_resp_desc_6_xuser_5_reg),
                                                                                               .wr_resp_desc_6_xuser_6_reg(wr_resp_desc_6_xuser_6_reg),
                                                                                               .wr_resp_desc_6_xuser_7_reg(wr_resp_desc_6_xuser_7_reg),
                                                                                               .wr_resp_desc_6_xuser_8_reg(wr_resp_desc_6_xuser_8_reg),
                                                                                               .wr_resp_desc_6_xuser_9_reg(wr_resp_desc_6_xuser_9_reg),
                                                                                               .wr_resp_desc_6_xuser_10_reg(wr_resp_desc_6_xuser_10_reg),
                                                                                               .wr_resp_desc_6_xuser_11_reg(wr_resp_desc_6_xuser_11_reg),
                                                                                               .wr_resp_desc_6_xuser_12_reg(wr_resp_desc_6_xuser_12_reg),
                                                                                               .wr_resp_desc_6_xuser_13_reg(wr_resp_desc_6_xuser_13_reg),
                                                                                               .wr_resp_desc_6_xuser_14_reg(wr_resp_desc_6_xuser_14_reg),
                                                                                               .wr_resp_desc_6_xuser_15_reg(wr_resp_desc_6_xuser_15_reg),
                                                                                               .sn_req_desc_6_attr_reg(sn_req_desc_6_attr_reg),
                                                                                               .sn_req_desc_6_acaddr_0_reg(sn_req_desc_6_acaddr_0_reg),
                                                                                               .sn_req_desc_6_acaddr_1_reg(sn_req_desc_6_acaddr_1_reg),
                                                                                               .sn_req_desc_6_acaddr_2_reg(sn_req_desc_6_acaddr_2_reg),
                                                                                               .sn_req_desc_6_acaddr_3_reg(sn_req_desc_6_acaddr_3_reg),
                                                                                               .sn_resp_desc_6_resp_reg(sn_resp_desc_6_resp_reg),
                                                                                               .rd_req_desc_7_txn_type_reg(rd_req_desc_7_txn_type_reg),
                                                                                               .rd_req_desc_7_size_reg(rd_req_desc_7_size_reg),
                                                                                               .rd_req_desc_7_axsize_reg(rd_req_desc_7_axsize_reg),
                                                                                               .rd_req_desc_7_attr_reg(rd_req_desc_7_attr_reg),
                                                                                               .rd_req_desc_7_axaddr_0_reg(rd_req_desc_7_axaddr_0_reg),
                                                                                               .rd_req_desc_7_axaddr_1_reg(rd_req_desc_7_axaddr_1_reg),
                                                                                               .rd_req_desc_7_axaddr_2_reg(rd_req_desc_7_axaddr_2_reg),
                                                                                               .rd_req_desc_7_axaddr_3_reg(rd_req_desc_7_axaddr_3_reg),
                                                                                               .rd_req_desc_7_axid_0_reg(rd_req_desc_7_axid_0_reg),
                                                                                               .rd_req_desc_7_axid_1_reg(rd_req_desc_7_axid_1_reg),
                                                                                               .rd_req_desc_7_axid_2_reg(rd_req_desc_7_axid_2_reg),
                                                                                               .rd_req_desc_7_axid_3_reg(rd_req_desc_7_axid_3_reg),
                                                                                               .rd_req_desc_7_axuser_0_reg(rd_req_desc_7_axuser_0_reg),
                                                                                               .rd_req_desc_7_axuser_1_reg(rd_req_desc_7_axuser_1_reg),
                                                                                               .rd_req_desc_7_axuser_2_reg(rd_req_desc_7_axuser_2_reg),
                                                                                               .rd_req_desc_7_axuser_3_reg(rd_req_desc_7_axuser_3_reg),
                                                                                               .rd_req_desc_7_axuser_4_reg(rd_req_desc_7_axuser_4_reg),
                                                                                               .rd_req_desc_7_axuser_5_reg(rd_req_desc_7_axuser_5_reg),
                                                                                               .rd_req_desc_7_axuser_6_reg(rd_req_desc_7_axuser_6_reg),
                                                                                               .rd_req_desc_7_axuser_7_reg(rd_req_desc_7_axuser_7_reg),
                                                                                               .rd_req_desc_7_axuser_8_reg(rd_req_desc_7_axuser_8_reg),
                                                                                               .rd_req_desc_7_axuser_9_reg(rd_req_desc_7_axuser_9_reg),
                                                                                               .rd_req_desc_7_axuser_10_reg(rd_req_desc_7_axuser_10_reg),
                                                                                               .rd_req_desc_7_axuser_11_reg(rd_req_desc_7_axuser_11_reg),
                                                                                               .rd_req_desc_7_axuser_12_reg(rd_req_desc_7_axuser_12_reg),
                                                                                               .rd_req_desc_7_axuser_13_reg(rd_req_desc_7_axuser_13_reg),
                                                                                               .rd_req_desc_7_axuser_14_reg(rd_req_desc_7_axuser_14_reg),
                                                                                               .rd_req_desc_7_axuser_15_reg(rd_req_desc_7_axuser_15_reg),
                                                                                               .rd_resp_desc_7_data_offset_reg(rd_resp_desc_7_data_offset_reg),
                                                                                               .rd_resp_desc_7_data_size_reg(rd_resp_desc_7_data_size_reg),
                                                                                               .rd_resp_desc_7_data_host_addr_0_reg(rd_resp_desc_7_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_7_data_host_addr_1_reg(rd_resp_desc_7_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_7_data_host_addr_2_reg(rd_resp_desc_7_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_7_data_host_addr_3_reg(rd_resp_desc_7_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_7_resp_reg(rd_resp_desc_7_resp_reg),
                                                                                               .rd_resp_desc_7_xid_0_reg(rd_resp_desc_7_xid_0_reg),
                                                                                               .rd_resp_desc_7_xid_1_reg(rd_resp_desc_7_xid_1_reg),
                                                                                               .rd_resp_desc_7_xid_2_reg(rd_resp_desc_7_xid_2_reg),
                                                                                               .rd_resp_desc_7_xid_3_reg(rd_resp_desc_7_xid_3_reg),
                                                                                               .rd_resp_desc_7_xuser_0_reg(rd_resp_desc_7_xuser_0_reg),
                                                                                               .rd_resp_desc_7_xuser_1_reg(rd_resp_desc_7_xuser_1_reg),
                                                                                               .rd_resp_desc_7_xuser_2_reg(rd_resp_desc_7_xuser_2_reg),
                                                                                               .rd_resp_desc_7_xuser_3_reg(rd_resp_desc_7_xuser_3_reg),
                                                                                               .rd_resp_desc_7_xuser_4_reg(rd_resp_desc_7_xuser_4_reg),
                                                                                               .rd_resp_desc_7_xuser_5_reg(rd_resp_desc_7_xuser_5_reg),
                                                                                               .rd_resp_desc_7_xuser_6_reg(rd_resp_desc_7_xuser_6_reg),
                                                                                               .rd_resp_desc_7_xuser_7_reg(rd_resp_desc_7_xuser_7_reg),
                                                                                               .rd_resp_desc_7_xuser_8_reg(rd_resp_desc_7_xuser_8_reg),
                                                                                               .rd_resp_desc_7_xuser_9_reg(rd_resp_desc_7_xuser_9_reg),
                                                                                               .rd_resp_desc_7_xuser_10_reg(rd_resp_desc_7_xuser_10_reg),
                                                                                               .rd_resp_desc_7_xuser_11_reg(rd_resp_desc_7_xuser_11_reg),
                                                                                               .rd_resp_desc_7_xuser_12_reg(rd_resp_desc_7_xuser_12_reg),
                                                                                               .rd_resp_desc_7_xuser_13_reg(rd_resp_desc_7_xuser_13_reg),
                                                                                               .rd_resp_desc_7_xuser_14_reg(rd_resp_desc_7_xuser_14_reg),
                                                                                               .rd_resp_desc_7_xuser_15_reg(rd_resp_desc_7_xuser_15_reg),
                                                                                               .wr_req_desc_7_txn_type_reg(wr_req_desc_7_txn_type_reg),
                                                                                               .wr_req_desc_7_size_reg(wr_req_desc_7_size_reg),
                                                                                               .wr_req_desc_7_data_offset_reg(wr_req_desc_7_data_offset_reg),
                                                                                               .wr_req_desc_7_data_host_addr_0_reg(wr_req_desc_7_data_host_addr_0_reg),
                                                                                               .wr_req_desc_7_data_host_addr_1_reg(wr_req_desc_7_data_host_addr_1_reg),
                                                                                               .wr_req_desc_7_data_host_addr_2_reg(wr_req_desc_7_data_host_addr_2_reg),
                                                                                               .wr_req_desc_7_data_host_addr_3_reg(wr_req_desc_7_data_host_addr_3_reg),
                                                                                               .wr_req_desc_7_wstrb_host_addr_0_reg(wr_req_desc_7_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_7_wstrb_host_addr_1_reg(wr_req_desc_7_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_7_wstrb_host_addr_2_reg(wr_req_desc_7_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_7_wstrb_host_addr_3_reg(wr_req_desc_7_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_7_axsize_reg(wr_req_desc_7_axsize_reg),
                                                                                               .wr_req_desc_7_attr_reg(wr_req_desc_7_attr_reg),
                                                                                               .wr_req_desc_7_axaddr_0_reg(wr_req_desc_7_axaddr_0_reg),
                                                                                               .wr_req_desc_7_axaddr_1_reg(wr_req_desc_7_axaddr_1_reg),
                                                                                               .wr_req_desc_7_axaddr_2_reg(wr_req_desc_7_axaddr_2_reg),
                                                                                               .wr_req_desc_7_axaddr_3_reg(wr_req_desc_7_axaddr_3_reg),
                                                                                               .wr_req_desc_7_axid_0_reg(wr_req_desc_7_axid_0_reg),
                                                                                               .wr_req_desc_7_axid_1_reg(wr_req_desc_7_axid_1_reg),
                                                                                               .wr_req_desc_7_axid_2_reg(wr_req_desc_7_axid_2_reg),
                                                                                               .wr_req_desc_7_axid_3_reg(wr_req_desc_7_axid_3_reg),
                                                                                               .wr_req_desc_7_axuser_0_reg(wr_req_desc_7_axuser_0_reg),
                                                                                               .wr_req_desc_7_axuser_1_reg(wr_req_desc_7_axuser_1_reg),
                                                                                               .wr_req_desc_7_axuser_2_reg(wr_req_desc_7_axuser_2_reg),
                                                                                               .wr_req_desc_7_axuser_3_reg(wr_req_desc_7_axuser_3_reg),
                                                                                               .wr_req_desc_7_axuser_4_reg(wr_req_desc_7_axuser_4_reg),
                                                                                               .wr_req_desc_7_axuser_5_reg(wr_req_desc_7_axuser_5_reg),
                                                                                               .wr_req_desc_7_axuser_6_reg(wr_req_desc_7_axuser_6_reg),
                                                                                               .wr_req_desc_7_axuser_7_reg(wr_req_desc_7_axuser_7_reg),
                                                                                               .wr_req_desc_7_axuser_8_reg(wr_req_desc_7_axuser_8_reg),
                                                                                               .wr_req_desc_7_axuser_9_reg(wr_req_desc_7_axuser_9_reg),
                                                                                               .wr_req_desc_7_axuser_10_reg(wr_req_desc_7_axuser_10_reg),
                                                                                               .wr_req_desc_7_axuser_11_reg(wr_req_desc_7_axuser_11_reg),
                                                                                               .wr_req_desc_7_axuser_12_reg(wr_req_desc_7_axuser_12_reg),
                                                                                               .wr_req_desc_7_axuser_13_reg(wr_req_desc_7_axuser_13_reg),
                                                                                               .wr_req_desc_7_axuser_14_reg(wr_req_desc_7_axuser_14_reg),
                                                                                               .wr_req_desc_7_axuser_15_reg(wr_req_desc_7_axuser_15_reg),
                                                                                               .wr_req_desc_7_wuser_0_reg(wr_req_desc_7_wuser_0_reg),
                                                                                               .wr_req_desc_7_wuser_1_reg(wr_req_desc_7_wuser_1_reg),
                                                                                               .wr_req_desc_7_wuser_2_reg(wr_req_desc_7_wuser_2_reg),
                                                                                               .wr_req_desc_7_wuser_3_reg(wr_req_desc_7_wuser_3_reg),
                                                                                               .wr_req_desc_7_wuser_4_reg(wr_req_desc_7_wuser_4_reg),
                                                                                               .wr_req_desc_7_wuser_5_reg(wr_req_desc_7_wuser_5_reg),
                                                                                               .wr_req_desc_7_wuser_6_reg(wr_req_desc_7_wuser_6_reg),
                                                                                               .wr_req_desc_7_wuser_7_reg(wr_req_desc_7_wuser_7_reg),
                                                                                               .wr_req_desc_7_wuser_8_reg(wr_req_desc_7_wuser_8_reg),
                                                                                               .wr_req_desc_7_wuser_9_reg(wr_req_desc_7_wuser_9_reg),
                                                                                               .wr_req_desc_7_wuser_10_reg(wr_req_desc_7_wuser_10_reg),
                                                                                               .wr_req_desc_7_wuser_11_reg(wr_req_desc_7_wuser_11_reg),
                                                                                               .wr_req_desc_7_wuser_12_reg(wr_req_desc_7_wuser_12_reg),
                                                                                               .wr_req_desc_7_wuser_13_reg(wr_req_desc_7_wuser_13_reg),
                                                                                               .wr_req_desc_7_wuser_14_reg(wr_req_desc_7_wuser_14_reg),
                                                                                               .wr_req_desc_7_wuser_15_reg(wr_req_desc_7_wuser_15_reg),
                                                                                               .wr_resp_desc_7_resp_reg(wr_resp_desc_7_resp_reg),
                                                                                               .wr_resp_desc_7_xid_0_reg(wr_resp_desc_7_xid_0_reg),
                                                                                               .wr_resp_desc_7_xid_1_reg(wr_resp_desc_7_xid_1_reg),
                                                                                               .wr_resp_desc_7_xid_2_reg(wr_resp_desc_7_xid_2_reg),
                                                                                               .wr_resp_desc_7_xid_3_reg(wr_resp_desc_7_xid_3_reg),
                                                                                               .wr_resp_desc_7_xuser_0_reg(wr_resp_desc_7_xuser_0_reg),
                                                                                               .wr_resp_desc_7_xuser_1_reg(wr_resp_desc_7_xuser_1_reg),
                                                                                               .wr_resp_desc_7_xuser_2_reg(wr_resp_desc_7_xuser_2_reg),
                                                                                               .wr_resp_desc_7_xuser_3_reg(wr_resp_desc_7_xuser_3_reg),
                                                                                               .wr_resp_desc_7_xuser_4_reg(wr_resp_desc_7_xuser_4_reg),
                                                                                               .wr_resp_desc_7_xuser_5_reg(wr_resp_desc_7_xuser_5_reg),
                                                                                               .wr_resp_desc_7_xuser_6_reg(wr_resp_desc_7_xuser_6_reg),
                                                                                               .wr_resp_desc_7_xuser_7_reg(wr_resp_desc_7_xuser_7_reg),
                                                                                               .wr_resp_desc_7_xuser_8_reg(wr_resp_desc_7_xuser_8_reg),
                                                                                               .wr_resp_desc_7_xuser_9_reg(wr_resp_desc_7_xuser_9_reg),
                                                                                               .wr_resp_desc_7_xuser_10_reg(wr_resp_desc_7_xuser_10_reg),
                                                                                               .wr_resp_desc_7_xuser_11_reg(wr_resp_desc_7_xuser_11_reg),
                                                                                               .wr_resp_desc_7_xuser_12_reg(wr_resp_desc_7_xuser_12_reg),
                                                                                               .wr_resp_desc_7_xuser_13_reg(wr_resp_desc_7_xuser_13_reg),
                                                                                               .wr_resp_desc_7_xuser_14_reg(wr_resp_desc_7_xuser_14_reg),
                                                                                               .wr_resp_desc_7_xuser_15_reg(wr_resp_desc_7_xuser_15_reg),
                                                                                               .sn_req_desc_7_attr_reg(sn_req_desc_7_attr_reg),
                                                                                               .sn_req_desc_7_acaddr_0_reg(sn_req_desc_7_acaddr_0_reg),
                                                                                               .sn_req_desc_7_acaddr_1_reg(sn_req_desc_7_acaddr_1_reg),
                                                                                               .sn_req_desc_7_acaddr_2_reg(sn_req_desc_7_acaddr_2_reg),
                                                                                               .sn_req_desc_7_acaddr_3_reg(sn_req_desc_7_acaddr_3_reg),
                                                                                               .sn_resp_desc_7_resp_reg(sn_resp_desc_7_resp_reg),
                                                                                               .rd_req_desc_8_txn_type_reg(rd_req_desc_8_txn_type_reg),
                                                                                               .rd_req_desc_8_size_reg(rd_req_desc_8_size_reg),
                                                                                               .rd_req_desc_8_axsize_reg(rd_req_desc_8_axsize_reg),
                                                                                               .rd_req_desc_8_attr_reg(rd_req_desc_8_attr_reg),
                                                                                               .rd_req_desc_8_axaddr_0_reg(rd_req_desc_8_axaddr_0_reg),
                                                                                               .rd_req_desc_8_axaddr_1_reg(rd_req_desc_8_axaddr_1_reg),
                                                                                               .rd_req_desc_8_axaddr_2_reg(rd_req_desc_8_axaddr_2_reg),
                                                                                               .rd_req_desc_8_axaddr_3_reg(rd_req_desc_8_axaddr_3_reg),
                                                                                               .rd_req_desc_8_axid_0_reg(rd_req_desc_8_axid_0_reg),
                                                                                               .rd_req_desc_8_axid_1_reg(rd_req_desc_8_axid_1_reg),
                                                                                               .rd_req_desc_8_axid_2_reg(rd_req_desc_8_axid_2_reg),
                                                                                               .rd_req_desc_8_axid_3_reg(rd_req_desc_8_axid_3_reg),
                                                                                               .rd_req_desc_8_axuser_0_reg(rd_req_desc_8_axuser_0_reg),
                                                                                               .rd_req_desc_8_axuser_1_reg(rd_req_desc_8_axuser_1_reg),
                                                                                               .rd_req_desc_8_axuser_2_reg(rd_req_desc_8_axuser_2_reg),
                                                                                               .rd_req_desc_8_axuser_3_reg(rd_req_desc_8_axuser_3_reg),
                                                                                               .rd_req_desc_8_axuser_4_reg(rd_req_desc_8_axuser_4_reg),
                                                                                               .rd_req_desc_8_axuser_5_reg(rd_req_desc_8_axuser_5_reg),
                                                                                               .rd_req_desc_8_axuser_6_reg(rd_req_desc_8_axuser_6_reg),
                                                                                               .rd_req_desc_8_axuser_7_reg(rd_req_desc_8_axuser_7_reg),
                                                                                               .rd_req_desc_8_axuser_8_reg(rd_req_desc_8_axuser_8_reg),
                                                                                               .rd_req_desc_8_axuser_9_reg(rd_req_desc_8_axuser_9_reg),
                                                                                               .rd_req_desc_8_axuser_10_reg(rd_req_desc_8_axuser_10_reg),
                                                                                               .rd_req_desc_8_axuser_11_reg(rd_req_desc_8_axuser_11_reg),
                                                                                               .rd_req_desc_8_axuser_12_reg(rd_req_desc_8_axuser_12_reg),
                                                                                               .rd_req_desc_8_axuser_13_reg(rd_req_desc_8_axuser_13_reg),
                                                                                               .rd_req_desc_8_axuser_14_reg(rd_req_desc_8_axuser_14_reg),
                                                                                               .rd_req_desc_8_axuser_15_reg(rd_req_desc_8_axuser_15_reg),
                                                                                               .rd_resp_desc_8_data_offset_reg(rd_resp_desc_8_data_offset_reg),
                                                                                               .rd_resp_desc_8_data_size_reg(rd_resp_desc_8_data_size_reg),
                                                                                               .rd_resp_desc_8_data_host_addr_0_reg(rd_resp_desc_8_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_8_data_host_addr_1_reg(rd_resp_desc_8_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_8_data_host_addr_2_reg(rd_resp_desc_8_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_8_data_host_addr_3_reg(rd_resp_desc_8_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_8_resp_reg(rd_resp_desc_8_resp_reg),
                                                                                               .rd_resp_desc_8_xid_0_reg(rd_resp_desc_8_xid_0_reg),
                                                                                               .rd_resp_desc_8_xid_1_reg(rd_resp_desc_8_xid_1_reg),
                                                                                               .rd_resp_desc_8_xid_2_reg(rd_resp_desc_8_xid_2_reg),
                                                                                               .rd_resp_desc_8_xid_3_reg(rd_resp_desc_8_xid_3_reg),
                                                                                               .rd_resp_desc_8_xuser_0_reg(rd_resp_desc_8_xuser_0_reg),
                                                                                               .rd_resp_desc_8_xuser_1_reg(rd_resp_desc_8_xuser_1_reg),
                                                                                               .rd_resp_desc_8_xuser_2_reg(rd_resp_desc_8_xuser_2_reg),
                                                                                               .rd_resp_desc_8_xuser_3_reg(rd_resp_desc_8_xuser_3_reg),
                                                                                               .rd_resp_desc_8_xuser_4_reg(rd_resp_desc_8_xuser_4_reg),
                                                                                               .rd_resp_desc_8_xuser_5_reg(rd_resp_desc_8_xuser_5_reg),
                                                                                               .rd_resp_desc_8_xuser_6_reg(rd_resp_desc_8_xuser_6_reg),
                                                                                               .rd_resp_desc_8_xuser_7_reg(rd_resp_desc_8_xuser_7_reg),
                                                                                               .rd_resp_desc_8_xuser_8_reg(rd_resp_desc_8_xuser_8_reg),
                                                                                               .rd_resp_desc_8_xuser_9_reg(rd_resp_desc_8_xuser_9_reg),
                                                                                               .rd_resp_desc_8_xuser_10_reg(rd_resp_desc_8_xuser_10_reg),
                                                                                               .rd_resp_desc_8_xuser_11_reg(rd_resp_desc_8_xuser_11_reg),
                                                                                               .rd_resp_desc_8_xuser_12_reg(rd_resp_desc_8_xuser_12_reg),
                                                                                               .rd_resp_desc_8_xuser_13_reg(rd_resp_desc_8_xuser_13_reg),
                                                                                               .rd_resp_desc_8_xuser_14_reg(rd_resp_desc_8_xuser_14_reg),
                                                                                               .rd_resp_desc_8_xuser_15_reg(rd_resp_desc_8_xuser_15_reg),
                                                                                               .wr_req_desc_8_txn_type_reg(wr_req_desc_8_txn_type_reg),
                                                                                               .wr_req_desc_8_size_reg(wr_req_desc_8_size_reg),
                                                                                               .wr_req_desc_8_data_offset_reg(wr_req_desc_8_data_offset_reg),
                                                                                               .wr_req_desc_8_data_host_addr_0_reg(wr_req_desc_8_data_host_addr_0_reg),
                                                                                               .wr_req_desc_8_data_host_addr_1_reg(wr_req_desc_8_data_host_addr_1_reg),
                                                                                               .wr_req_desc_8_data_host_addr_2_reg(wr_req_desc_8_data_host_addr_2_reg),
                                                                                               .wr_req_desc_8_data_host_addr_3_reg(wr_req_desc_8_data_host_addr_3_reg),
                                                                                               .wr_req_desc_8_wstrb_host_addr_0_reg(wr_req_desc_8_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_8_wstrb_host_addr_1_reg(wr_req_desc_8_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_8_wstrb_host_addr_2_reg(wr_req_desc_8_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_8_wstrb_host_addr_3_reg(wr_req_desc_8_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_8_axsize_reg(wr_req_desc_8_axsize_reg),
                                                                                               .wr_req_desc_8_attr_reg(wr_req_desc_8_attr_reg),
                                                                                               .wr_req_desc_8_axaddr_0_reg(wr_req_desc_8_axaddr_0_reg),
                                                                                               .wr_req_desc_8_axaddr_1_reg(wr_req_desc_8_axaddr_1_reg),
                                                                                               .wr_req_desc_8_axaddr_2_reg(wr_req_desc_8_axaddr_2_reg),
                                                                                               .wr_req_desc_8_axaddr_3_reg(wr_req_desc_8_axaddr_3_reg),
                                                                                               .wr_req_desc_8_axid_0_reg(wr_req_desc_8_axid_0_reg),
                                                                                               .wr_req_desc_8_axid_1_reg(wr_req_desc_8_axid_1_reg),
                                                                                               .wr_req_desc_8_axid_2_reg(wr_req_desc_8_axid_2_reg),
                                                                                               .wr_req_desc_8_axid_3_reg(wr_req_desc_8_axid_3_reg),
                                                                                               .wr_req_desc_8_axuser_0_reg(wr_req_desc_8_axuser_0_reg),
                                                                                               .wr_req_desc_8_axuser_1_reg(wr_req_desc_8_axuser_1_reg),
                                                                                               .wr_req_desc_8_axuser_2_reg(wr_req_desc_8_axuser_2_reg),
                                                                                               .wr_req_desc_8_axuser_3_reg(wr_req_desc_8_axuser_3_reg),
                                                                                               .wr_req_desc_8_axuser_4_reg(wr_req_desc_8_axuser_4_reg),
                                                                                               .wr_req_desc_8_axuser_5_reg(wr_req_desc_8_axuser_5_reg),
                                                                                               .wr_req_desc_8_axuser_6_reg(wr_req_desc_8_axuser_6_reg),
                                                                                               .wr_req_desc_8_axuser_7_reg(wr_req_desc_8_axuser_7_reg),
                                                                                               .wr_req_desc_8_axuser_8_reg(wr_req_desc_8_axuser_8_reg),
                                                                                               .wr_req_desc_8_axuser_9_reg(wr_req_desc_8_axuser_9_reg),
                                                                                               .wr_req_desc_8_axuser_10_reg(wr_req_desc_8_axuser_10_reg),
                                                                                               .wr_req_desc_8_axuser_11_reg(wr_req_desc_8_axuser_11_reg),
                                                                                               .wr_req_desc_8_axuser_12_reg(wr_req_desc_8_axuser_12_reg),
                                                                                               .wr_req_desc_8_axuser_13_reg(wr_req_desc_8_axuser_13_reg),
                                                                                               .wr_req_desc_8_axuser_14_reg(wr_req_desc_8_axuser_14_reg),
                                                                                               .wr_req_desc_8_axuser_15_reg(wr_req_desc_8_axuser_15_reg),
                                                                                               .wr_req_desc_8_wuser_0_reg(wr_req_desc_8_wuser_0_reg),
                                                                                               .wr_req_desc_8_wuser_1_reg(wr_req_desc_8_wuser_1_reg),
                                                                                               .wr_req_desc_8_wuser_2_reg(wr_req_desc_8_wuser_2_reg),
                                                                                               .wr_req_desc_8_wuser_3_reg(wr_req_desc_8_wuser_3_reg),
                                                                                               .wr_req_desc_8_wuser_4_reg(wr_req_desc_8_wuser_4_reg),
                                                                                               .wr_req_desc_8_wuser_5_reg(wr_req_desc_8_wuser_5_reg),
                                                                                               .wr_req_desc_8_wuser_6_reg(wr_req_desc_8_wuser_6_reg),
                                                                                               .wr_req_desc_8_wuser_7_reg(wr_req_desc_8_wuser_7_reg),
                                                                                               .wr_req_desc_8_wuser_8_reg(wr_req_desc_8_wuser_8_reg),
                                                                                               .wr_req_desc_8_wuser_9_reg(wr_req_desc_8_wuser_9_reg),
                                                                                               .wr_req_desc_8_wuser_10_reg(wr_req_desc_8_wuser_10_reg),
                                                                                               .wr_req_desc_8_wuser_11_reg(wr_req_desc_8_wuser_11_reg),
                                                                                               .wr_req_desc_8_wuser_12_reg(wr_req_desc_8_wuser_12_reg),
                                                                                               .wr_req_desc_8_wuser_13_reg(wr_req_desc_8_wuser_13_reg),
                                                                                               .wr_req_desc_8_wuser_14_reg(wr_req_desc_8_wuser_14_reg),
                                                                                               .wr_req_desc_8_wuser_15_reg(wr_req_desc_8_wuser_15_reg),
                                                                                               .wr_resp_desc_8_resp_reg(wr_resp_desc_8_resp_reg),
                                                                                               .wr_resp_desc_8_xid_0_reg(wr_resp_desc_8_xid_0_reg),
                                                                                               .wr_resp_desc_8_xid_1_reg(wr_resp_desc_8_xid_1_reg),
                                                                                               .wr_resp_desc_8_xid_2_reg(wr_resp_desc_8_xid_2_reg),
                                                                                               .wr_resp_desc_8_xid_3_reg(wr_resp_desc_8_xid_3_reg),
                                                                                               .wr_resp_desc_8_xuser_0_reg(wr_resp_desc_8_xuser_0_reg),
                                                                                               .wr_resp_desc_8_xuser_1_reg(wr_resp_desc_8_xuser_1_reg),
                                                                                               .wr_resp_desc_8_xuser_2_reg(wr_resp_desc_8_xuser_2_reg),
                                                                                               .wr_resp_desc_8_xuser_3_reg(wr_resp_desc_8_xuser_3_reg),
                                                                                               .wr_resp_desc_8_xuser_4_reg(wr_resp_desc_8_xuser_4_reg),
                                                                                               .wr_resp_desc_8_xuser_5_reg(wr_resp_desc_8_xuser_5_reg),
                                                                                               .wr_resp_desc_8_xuser_6_reg(wr_resp_desc_8_xuser_6_reg),
                                                                                               .wr_resp_desc_8_xuser_7_reg(wr_resp_desc_8_xuser_7_reg),
                                                                                               .wr_resp_desc_8_xuser_8_reg(wr_resp_desc_8_xuser_8_reg),
                                                                                               .wr_resp_desc_8_xuser_9_reg(wr_resp_desc_8_xuser_9_reg),
                                                                                               .wr_resp_desc_8_xuser_10_reg(wr_resp_desc_8_xuser_10_reg),
                                                                                               .wr_resp_desc_8_xuser_11_reg(wr_resp_desc_8_xuser_11_reg),
                                                                                               .wr_resp_desc_8_xuser_12_reg(wr_resp_desc_8_xuser_12_reg),
                                                                                               .wr_resp_desc_8_xuser_13_reg(wr_resp_desc_8_xuser_13_reg),
                                                                                               .wr_resp_desc_8_xuser_14_reg(wr_resp_desc_8_xuser_14_reg),
                                                                                               .wr_resp_desc_8_xuser_15_reg(wr_resp_desc_8_xuser_15_reg),
                                                                                               .sn_req_desc_8_attr_reg(sn_req_desc_8_attr_reg),
                                                                                               .sn_req_desc_8_acaddr_0_reg(sn_req_desc_8_acaddr_0_reg),
                                                                                               .sn_req_desc_8_acaddr_1_reg(sn_req_desc_8_acaddr_1_reg),
                                                                                               .sn_req_desc_8_acaddr_2_reg(sn_req_desc_8_acaddr_2_reg),
                                                                                               .sn_req_desc_8_acaddr_3_reg(sn_req_desc_8_acaddr_3_reg),
                                                                                               .sn_resp_desc_8_resp_reg(sn_resp_desc_8_resp_reg),
                                                                                               .rd_req_desc_9_txn_type_reg(rd_req_desc_9_txn_type_reg),
                                                                                               .rd_req_desc_9_size_reg(rd_req_desc_9_size_reg),
                                                                                               .rd_req_desc_9_axsize_reg(rd_req_desc_9_axsize_reg),
                                                                                               .rd_req_desc_9_attr_reg(rd_req_desc_9_attr_reg),
                                                                                               .rd_req_desc_9_axaddr_0_reg(rd_req_desc_9_axaddr_0_reg),
                                                                                               .rd_req_desc_9_axaddr_1_reg(rd_req_desc_9_axaddr_1_reg),
                                                                                               .rd_req_desc_9_axaddr_2_reg(rd_req_desc_9_axaddr_2_reg),
                                                                                               .rd_req_desc_9_axaddr_3_reg(rd_req_desc_9_axaddr_3_reg),
                                                                                               .rd_req_desc_9_axid_0_reg(rd_req_desc_9_axid_0_reg),
                                                                                               .rd_req_desc_9_axid_1_reg(rd_req_desc_9_axid_1_reg),
                                                                                               .rd_req_desc_9_axid_2_reg(rd_req_desc_9_axid_2_reg),
                                                                                               .rd_req_desc_9_axid_3_reg(rd_req_desc_9_axid_3_reg),
                                                                                               .rd_req_desc_9_axuser_0_reg(rd_req_desc_9_axuser_0_reg),
                                                                                               .rd_req_desc_9_axuser_1_reg(rd_req_desc_9_axuser_1_reg),
                                                                                               .rd_req_desc_9_axuser_2_reg(rd_req_desc_9_axuser_2_reg),
                                                                                               .rd_req_desc_9_axuser_3_reg(rd_req_desc_9_axuser_3_reg),
                                                                                               .rd_req_desc_9_axuser_4_reg(rd_req_desc_9_axuser_4_reg),
                                                                                               .rd_req_desc_9_axuser_5_reg(rd_req_desc_9_axuser_5_reg),
                                                                                               .rd_req_desc_9_axuser_6_reg(rd_req_desc_9_axuser_6_reg),
                                                                                               .rd_req_desc_9_axuser_7_reg(rd_req_desc_9_axuser_7_reg),
                                                                                               .rd_req_desc_9_axuser_8_reg(rd_req_desc_9_axuser_8_reg),
                                                                                               .rd_req_desc_9_axuser_9_reg(rd_req_desc_9_axuser_9_reg),
                                                                                               .rd_req_desc_9_axuser_10_reg(rd_req_desc_9_axuser_10_reg),
                                                                                               .rd_req_desc_9_axuser_11_reg(rd_req_desc_9_axuser_11_reg),
                                                                                               .rd_req_desc_9_axuser_12_reg(rd_req_desc_9_axuser_12_reg),
                                                                                               .rd_req_desc_9_axuser_13_reg(rd_req_desc_9_axuser_13_reg),
                                                                                               .rd_req_desc_9_axuser_14_reg(rd_req_desc_9_axuser_14_reg),
                                                                                               .rd_req_desc_9_axuser_15_reg(rd_req_desc_9_axuser_15_reg),
                                                                                               .rd_resp_desc_9_data_offset_reg(rd_resp_desc_9_data_offset_reg),
                                                                                               .rd_resp_desc_9_data_size_reg(rd_resp_desc_9_data_size_reg),
                                                                                               .rd_resp_desc_9_data_host_addr_0_reg(rd_resp_desc_9_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_9_data_host_addr_1_reg(rd_resp_desc_9_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_9_data_host_addr_2_reg(rd_resp_desc_9_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_9_data_host_addr_3_reg(rd_resp_desc_9_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_9_resp_reg(rd_resp_desc_9_resp_reg),
                                                                                               .rd_resp_desc_9_xid_0_reg(rd_resp_desc_9_xid_0_reg),
                                                                                               .rd_resp_desc_9_xid_1_reg(rd_resp_desc_9_xid_1_reg),
                                                                                               .rd_resp_desc_9_xid_2_reg(rd_resp_desc_9_xid_2_reg),
                                                                                               .rd_resp_desc_9_xid_3_reg(rd_resp_desc_9_xid_3_reg),
                                                                                               .rd_resp_desc_9_xuser_0_reg(rd_resp_desc_9_xuser_0_reg),
                                                                                               .rd_resp_desc_9_xuser_1_reg(rd_resp_desc_9_xuser_1_reg),
                                                                                               .rd_resp_desc_9_xuser_2_reg(rd_resp_desc_9_xuser_2_reg),
                                                                                               .rd_resp_desc_9_xuser_3_reg(rd_resp_desc_9_xuser_3_reg),
                                                                                               .rd_resp_desc_9_xuser_4_reg(rd_resp_desc_9_xuser_4_reg),
                                                                                               .rd_resp_desc_9_xuser_5_reg(rd_resp_desc_9_xuser_5_reg),
                                                                                               .rd_resp_desc_9_xuser_6_reg(rd_resp_desc_9_xuser_6_reg),
                                                                                               .rd_resp_desc_9_xuser_7_reg(rd_resp_desc_9_xuser_7_reg),
                                                                                               .rd_resp_desc_9_xuser_8_reg(rd_resp_desc_9_xuser_8_reg),
                                                                                               .rd_resp_desc_9_xuser_9_reg(rd_resp_desc_9_xuser_9_reg),
                                                                                               .rd_resp_desc_9_xuser_10_reg(rd_resp_desc_9_xuser_10_reg),
                                                                                               .rd_resp_desc_9_xuser_11_reg(rd_resp_desc_9_xuser_11_reg),
                                                                                               .rd_resp_desc_9_xuser_12_reg(rd_resp_desc_9_xuser_12_reg),
                                                                                               .rd_resp_desc_9_xuser_13_reg(rd_resp_desc_9_xuser_13_reg),
                                                                                               .rd_resp_desc_9_xuser_14_reg(rd_resp_desc_9_xuser_14_reg),
                                                                                               .rd_resp_desc_9_xuser_15_reg(rd_resp_desc_9_xuser_15_reg),
                                                                                               .wr_req_desc_9_txn_type_reg(wr_req_desc_9_txn_type_reg),
                                                                                               .wr_req_desc_9_size_reg(wr_req_desc_9_size_reg),
                                                                                               .wr_req_desc_9_data_offset_reg(wr_req_desc_9_data_offset_reg),
                                                                                               .wr_req_desc_9_data_host_addr_0_reg(wr_req_desc_9_data_host_addr_0_reg),
                                                                                               .wr_req_desc_9_data_host_addr_1_reg(wr_req_desc_9_data_host_addr_1_reg),
                                                                                               .wr_req_desc_9_data_host_addr_2_reg(wr_req_desc_9_data_host_addr_2_reg),
                                                                                               .wr_req_desc_9_data_host_addr_3_reg(wr_req_desc_9_data_host_addr_3_reg),
                                                                                               .wr_req_desc_9_wstrb_host_addr_0_reg(wr_req_desc_9_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_9_wstrb_host_addr_1_reg(wr_req_desc_9_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_9_wstrb_host_addr_2_reg(wr_req_desc_9_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_9_wstrb_host_addr_3_reg(wr_req_desc_9_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_9_axsize_reg(wr_req_desc_9_axsize_reg),
                                                                                               .wr_req_desc_9_attr_reg(wr_req_desc_9_attr_reg),
                                                                                               .wr_req_desc_9_axaddr_0_reg(wr_req_desc_9_axaddr_0_reg),
                                                                                               .wr_req_desc_9_axaddr_1_reg(wr_req_desc_9_axaddr_1_reg),
                                                                                               .wr_req_desc_9_axaddr_2_reg(wr_req_desc_9_axaddr_2_reg),
                                                                                               .wr_req_desc_9_axaddr_3_reg(wr_req_desc_9_axaddr_3_reg),
                                                                                               .wr_req_desc_9_axid_0_reg(wr_req_desc_9_axid_0_reg),
                                                                                               .wr_req_desc_9_axid_1_reg(wr_req_desc_9_axid_1_reg),
                                                                                               .wr_req_desc_9_axid_2_reg(wr_req_desc_9_axid_2_reg),
                                                                                               .wr_req_desc_9_axid_3_reg(wr_req_desc_9_axid_3_reg),
                                                                                               .wr_req_desc_9_axuser_0_reg(wr_req_desc_9_axuser_0_reg),
                                                                                               .wr_req_desc_9_axuser_1_reg(wr_req_desc_9_axuser_1_reg),
                                                                                               .wr_req_desc_9_axuser_2_reg(wr_req_desc_9_axuser_2_reg),
                                                                                               .wr_req_desc_9_axuser_3_reg(wr_req_desc_9_axuser_3_reg),
                                                                                               .wr_req_desc_9_axuser_4_reg(wr_req_desc_9_axuser_4_reg),
                                                                                               .wr_req_desc_9_axuser_5_reg(wr_req_desc_9_axuser_5_reg),
                                                                                               .wr_req_desc_9_axuser_6_reg(wr_req_desc_9_axuser_6_reg),
                                                                                               .wr_req_desc_9_axuser_7_reg(wr_req_desc_9_axuser_7_reg),
                                                                                               .wr_req_desc_9_axuser_8_reg(wr_req_desc_9_axuser_8_reg),
                                                                                               .wr_req_desc_9_axuser_9_reg(wr_req_desc_9_axuser_9_reg),
                                                                                               .wr_req_desc_9_axuser_10_reg(wr_req_desc_9_axuser_10_reg),
                                                                                               .wr_req_desc_9_axuser_11_reg(wr_req_desc_9_axuser_11_reg),
                                                                                               .wr_req_desc_9_axuser_12_reg(wr_req_desc_9_axuser_12_reg),
                                                                                               .wr_req_desc_9_axuser_13_reg(wr_req_desc_9_axuser_13_reg),
                                                                                               .wr_req_desc_9_axuser_14_reg(wr_req_desc_9_axuser_14_reg),
                                                                                               .wr_req_desc_9_axuser_15_reg(wr_req_desc_9_axuser_15_reg),
                                                                                               .wr_req_desc_9_wuser_0_reg(wr_req_desc_9_wuser_0_reg),
                                                                                               .wr_req_desc_9_wuser_1_reg(wr_req_desc_9_wuser_1_reg),
                                                                                               .wr_req_desc_9_wuser_2_reg(wr_req_desc_9_wuser_2_reg),
                                                                                               .wr_req_desc_9_wuser_3_reg(wr_req_desc_9_wuser_3_reg),
                                                                                               .wr_req_desc_9_wuser_4_reg(wr_req_desc_9_wuser_4_reg),
                                                                                               .wr_req_desc_9_wuser_5_reg(wr_req_desc_9_wuser_5_reg),
                                                                                               .wr_req_desc_9_wuser_6_reg(wr_req_desc_9_wuser_6_reg),
                                                                                               .wr_req_desc_9_wuser_7_reg(wr_req_desc_9_wuser_7_reg),
                                                                                               .wr_req_desc_9_wuser_8_reg(wr_req_desc_9_wuser_8_reg),
                                                                                               .wr_req_desc_9_wuser_9_reg(wr_req_desc_9_wuser_9_reg),
                                                                                               .wr_req_desc_9_wuser_10_reg(wr_req_desc_9_wuser_10_reg),
                                                                                               .wr_req_desc_9_wuser_11_reg(wr_req_desc_9_wuser_11_reg),
                                                                                               .wr_req_desc_9_wuser_12_reg(wr_req_desc_9_wuser_12_reg),
                                                                                               .wr_req_desc_9_wuser_13_reg(wr_req_desc_9_wuser_13_reg),
                                                                                               .wr_req_desc_9_wuser_14_reg(wr_req_desc_9_wuser_14_reg),
                                                                                               .wr_req_desc_9_wuser_15_reg(wr_req_desc_9_wuser_15_reg),
                                                                                               .wr_resp_desc_9_resp_reg(wr_resp_desc_9_resp_reg),
                                                                                               .wr_resp_desc_9_xid_0_reg(wr_resp_desc_9_xid_0_reg),
                                                                                               .wr_resp_desc_9_xid_1_reg(wr_resp_desc_9_xid_1_reg),
                                                                                               .wr_resp_desc_9_xid_2_reg(wr_resp_desc_9_xid_2_reg),
                                                                                               .wr_resp_desc_9_xid_3_reg(wr_resp_desc_9_xid_3_reg),
                                                                                               .wr_resp_desc_9_xuser_0_reg(wr_resp_desc_9_xuser_0_reg),
                                                                                               .wr_resp_desc_9_xuser_1_reg(wr_resp_desc_9_xuser_1_reg),
                                                                                               .wr_resp_desc_9_xuser_2_reg(wr_resp_desc_9_xuser_2_reg),
                                                                                               .wr_resp_desc_9_xuser_3_reg(wr_resp_desc_9_xuser_3_reg),
                                                                                               .wr_resp_desc_9_xuser_4_reg(wr_resp_desc_9_xuser_4_reg),
                                                                                               .wr_resp_desc_9_xuser_5_reg(wr_resp_desc_9_xuser_5_reg),
                                                                                               .wr_resp_desc_9_xuser_6_reg(wr_resp_desc_9_xuser_6_reg),
                                                                                               .wr_resp_desc_9_xuser_7_reg(wr_resp_desc_9_xuser_7_reg),
                                                                                               .wr_resp_desc_9_xuser_8_reg(wr_resp_desc_9_xuser_8_reg),
                                                                                               .wr_resp_desc_9_xuser_9_reg(wr_resp_desc_9_xuser_9_reg),
                                                                                               .wr_resp_desc_9_xuser_10_reg(wr_resp_desc_9_xuser_10_reg),
                                                                                               .wr_resp_desc_9_xuser_11_reg(wr_resp_desc_9_xuser_11_reg),
                                                                                               .wr_resp_desc_9_xuser_12_reg(wr_resp_desc_9_xuser_12_reg),
                                                                                               .wr_resp_desc_9_xuser_13_reg(wr_resp_desc_9_xuser_13_reg),
                                                                                               .wr_resp_desc_9_xuser_14_reg(wr_resp_desc_9_xuser_14_reg),
                                                                                               .wr_resp_desc_9_xuser_15_reg(wr_resp_desc_9_xuser_15_reg),
                                                                                               .sn_req_desc_9_attr_reg(sn_req_desc_9_attr_reg),
                                                                                               .sn_req_desc_9_acaddr_0_reg(sn_req_desc_9_acaddr_0_reg),
                                                                                               .sn_req_desc_9_acaddr_1_reg(sn_req_desc_9_acaddr_1_reg),
                                                                                               .sn_req_desc_9_acaddr_2_reg(sn_req_desc_9_acaddr_2_reg),
                                                                                               .sn_req_desc_9_acaddr_3_reg(sn_req_desc_9_acaddr_3_reg),
                                                                                               .sn_resp_desc_9_resp_reg(sn_resp_desc_9_resp_reg),
                                                                                               .rd_req_desc_a_txn_type_reg(rd_req_desc_a_txn_type_reg),
                                                                                               .rd_req_desc_a_size_reg(rd_req_desc_a_size_reg),
                                                                                               .rd_req_desc_a_axsize_reg(rd_req_desc_a_axsize_reg),
                                                                                               .rd_req_desc_a_attr_reg(rd_req_desc_a_attr_reg),
                                                                                               .rd_req_desc_a_axaddr_0_reg(rd_req_desc_a_axaddr_0_reg),
                                                                                               .rd_req_desc_a_axaddr_1_reg(rd_req_desc_a_axaddr_1_reg),
                                                                                               .rd_req_desc_a_axaddr_2_reg(rd_req_desc_a_axaddr_2_reg),
                                                                                               .rd_req_desc_a_axaddr_3_reg(rd_req_desc_a_axaddr_3_reg),
                                                                                               .rd_req_desc_a_axid_0_reg(rd_req_desc_a_axid_0_reg),
                                                                                               .rd_req_desc_a_axid_1_reg(rd_req_desc_a_axid_1_reg),
                                                                                               .rd_req_desc_a_axid_2_reg(rd_req_desc_a_axid_2_reg),
                                                                                               .rd_req_desc_a_axid_3_reg(rd_req_desc_a_axid_3_reg),
                                                                                               .rd_req_desc_a_axuser_0_reg(rd_req_desc_a_axuser_0_reg),
                                                                                               .rd_req_desc_a_axuser_1_reg(rd_req_desc_a_axuser_1_reg),
                                                                                               .rd_req_desc_a_axuser_2_reg(rd_req_desc_a_axuser_2_reg),
                                                                                               .rd_req_desc_a_axuser_3_reg(rd_req_desc_a_axuser_3_reg),
                                                                                               .rd_req_desc_a_axuser_4_reg(rd_req_desc_a_axuser_4_reg),
                                                                                               .rd_req_desc_a_axuser_5_reg(rd_req_desc_a_axuser_5_reg),
                                                                                               .rd_req_desc_a_axuser_6_reg(rd_req_desc_a_axuser_6_reg),
                                                                                               .rd_req_desc_a_axuser_7_reg(rd_req_desc_a_axuser_7_reg),
                                                                                               .rd_req_desc_a_axuser_8_reg(rd_req_desc_a_axuser_8_reg),
                                                                                               .rd_req_desc_a_axuser_9_reg(rd_req_desc_a_axuser_9_reg),
                                                                                               .rd_req_desc_a_axuser_10_reg(rd_req_desc_a_axuser_10_reg),
                                                                                               .rd_req_desc_a_axuser_11_reg(rd_req_desc_a_axuser_11_reg),
                                                                                               .rd_req_desc_a_axuser_12_reg(rd_req_desc_a_axuser_12_reg),
                                                                                               .rd_req_desc_a_axuser_13_reg(rd_req_desc_a_axuser_13_reg),
                                                                                               .rd_req_desc_a_axuser_14_reg(rd_req_desc_a_axuser_14_reg),
                                                                                               .rd_req_desc_a_axuser_15_reg(rd_req_desc_a_axuser_15_reg),
                                                                                               .rd_resp_desc_a_data_offset_reg(rd_resp_desc_a_data_offset_reg),
                                                                                               .rd_resp_desc_a_data_size_reg(rd_resp_desc_a_data_size_reg),
                                                                                               .rd_resp_desc_a_data_host_addr_0_reg(rd_resp_desc_a_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_a_data_host_addr_1_reg(rd_resp_desc_a_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_a_data_host_addr_2_reg(rd_resp_desc_a_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_a_data_host_addr_3_reg(rd_resp_desc_a_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_a_resp_reg(rd_resp_desc_a_resp_reg),
                                                                                               .rd_resp_desc_a_xid_0_reg(rd_resp_desc_a_xid_0_reg),
                                                                                               .rd_resp_desc_a_xid_1_reg(rd_resp_desc_a_xid_1_reg),
                                                                                               .rd_resp_desc_a_xid_2_reg(rd_resp_desc_a_xid_2_reg),
                                                                                               .rd_resp_desc_a_xid_3_reg(rd_resp_desc_a_xid_3_reg),
                                                                                               .rd_resp_desc_a_xuser_0_reg(rd_resp_desc_a_xuser_0_reg),
                                                                                               .rd_resp_desc_a_xuser_1_reg(rd_resp_desc_a_xuser_1_reg),
                                                                                               .rd_resp_desc_a_xuser_2_reg(rd_resp_desc_a_xuser_2_reg),
                                                                                               .rd_resp_desc_a_xuser_3_reg(rd_resp_desc_a_xuser_3_reg),
                                                                                               .rd_resp_desc_a_xuser_4_reg(rd_resp_desc_a_xuser_4_reg),
                                                                                               .rd_resp_desc_a_xuser_5_reg(rd_resp_desc_a_xuser_5_reg),
                                                                                               .rd_resp_desc_a_xuser_6_reg(rd_resp_desc_a_xuser_6_reg),
                                                                                               .rd_resp_desc_a_xuser_7_reg(rd_resp_desc_a_xuser_7_reg),
                                                                                               .rd_resp_desc_a_xuser_8_reg(rd_resp_desc_a_xuser_8_reg),
                                                                                               .rd_resp_desc_a_xuser_9_reg(rd_resp_desc_a_xuser_9_reg),
                                                                                               .rd_resp_desc_a_xuser_10_reg(rd_resp_desc_a_xuser_10_reg),
                                                                                               .rd_resp_desc_a_xuser_11_reg(rd_resp_desc_a_xuser_11_reg),
                                                                                               .rd_resp_desc_a_xuser_12_reg(rd_resp_desc_a_xuser_12_reg),
                                                                                               .rd_resp_desc_a_xuser_13_reg(rd_resp_desc_a_xuser_13_reg),
                                                                                               .rd_resp_desc_a_xuser_14_reg(rd_resp_desc_a_xuser_14_reg),
                                                                                               .rd_resp_desc_a_xuser_15_reg(rd_resp_desc_a_xuser_15_reg),
                                                                                               .wr_req_desc_a_txn_type_reg(wr_req_desc_a_txn_type_reg),
                                                                                               .wr_req_desc_a_size_reg(wr_req_desc_a_size_reg),
                                                                                               .wr_req_desc_a_data_offset_reg(wr_req_desc_a_data_offset_reg),
                                                                                               .wr_req_desc_a_data_host_addr_0_reg(wr_req_desc_a_data_host_addr_0_reg),
                                                                                               .wr_req_desc_a_data_host_addr_1_reg(wr_req_desc_a_data_host_addr_1_reg),
                                                                                               .wr_req_desc_a_data_host_addr_2_reg(wr_req_desc_a_data_host_addr_2_reg),
                                                                                               .wr_req_desc_a_data_host_addr_3_reg(wr_req_desc_a_data_host_addr_3_reg),
                                                                                               .wr_req_desc_a_wstrb_host_addr_0_reg(wr_req_desc_a_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_a_wstrb_host_addr_1_reg(wr_req_desc_a_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_a_wstrb_host_addr_2_reg(wr_req_desc_a_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_a_wstrb_host_addr_3_reg(wr_req_desc_a_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_a_axsize_reg(wr_req_desc_a_axsize_reg),
                                                                                               .wr_req_desc_a_attr_reg(wr_req_desc_a_attr_reg),
                                                                                               .wr_req_desc_a_axaddr_0_reg(wr_req_desc_a_axaddr_0_reg),
                                                                                               .wr_req_desc_a_axaddr_1_reg(wr_req_desc_a_axaddr_1_reg),
                                                                                               .wr_req_desc_a_axaddr_2_reg(wr_req_desc_a_axaddr_2_reg),
                                                                                               .wr_req_desc_a_axaddr_3_reg(wr_req_desc_a_axaddr_3_reg),
                                                                                               .wr_req_desc_a_axid_0_reg(wr_req_desc_a_axid_0_reg),
                                                                                               .wr_req_desc_a_axid_1_reg(wr_req_desc_a_axid_1_reg),
                                                                                               .wr_req_desc_a_axid_2_reg(wr_req_desc_a_axid_2_reg),
                                                                                               .wr_req_desc_a_axid_3_reg(wr_req_desc_a_axid_3_reg),
                                                                                               .wr_req_desc_a_axuser_0_reg(wr_req_desc_a_axuser_0_reg),
                                                                                               .wr_req_desc_a_axuser_1_reg(wr_req_desc_a_axuser_1_reg),
                                                                                               .wr_req_desc_a_axuser_2_reg(wr_req_desc_a_axuser_2_reg),
                                                                                               .wr_req_desc_a_axuser_3_reg(wr_req_desc_a_axuser_3_reg),
                                                                                               .wr_req_desc_a_axuser_4_reg(wr_req_desc_a_axuser_4_reg),
                                                                                               .wr_req_desc_a_axuser_5_reg(wr_req_desc_a_axuser_5_reg),
                                                                                               .wr_req_desc_a_axuser_6_reg(wr_req_desc_a_axuser_6_reg),
                                                                                               .wr_req_desc_a_axuser_7_reg(wr_req_desc_a_axuser_7_reg),
                                                                                               .wr_req_desc_a_axuser_8_reg(wr_req_desc_a_axuser_8_reg),
                                                                                               .wr_req_desc_a_axuser_9_reg(wr_req_desc_a_axuser_9_reg),
                                                                                               .wr_req_desc_a_axuser_10_reg(wr_req_desc_a_axuser_10_reg),
                                                                                               .wr_req_desc_a_axuser_11_reg(wr_req_desc_a_axuser_11_reg),
                                                                                               .wr_req_desc_a_axuser_12_reg(wr_req_desc_a_axuser_12_reg),
                                                                                               .wr_req_desc_a_axuser_13_reg(wr_req_desc_a_axuser_13_reg),
                                                                                               .wr_req_desc_a_axuser_14_reg(wr_req_desc_a_axuser_14_reg),
                                                                                               .wr_req_desc_a_axuser_15_reg(wr_req_desc_a_axuser_15_reg),
                                                                                               .wr_req_desc_a_wuser_0_reg(wr_req_desc_a_wuser_0_reg),
                                                                                               .wr_req_desc_a_wuser_1_reg(wr_req_desc_a_wuser_1_reg),
                                                                                               .wr_req_desc_a_wuser_2_reg(wr_req_desc_a_wuser_2_reg),
                                                                                               .wr_req_desc_a_wuser_3_reg(wr_req_desc_a_wuser_3_reg),
                                                                                               .wr_req_desc_a_wuser_4_reg(wr_req_desc_a_wuser_4_reg),
                                                                                               .wr_req_desc_a_wuser_5_reg(wr_req_desc_a_wuser_5_reg),
                                                                                               .wr_req_desc_a_wuser_6_reg(wr_req_desc_a_wuser_6_reg),
                                                                                               .wr_req_desc_a_wuser_7_reg(wr_req_desc_a_wuser_7_reg),
                                                                                               .wr_req_desc_a_wuser_8_reg(wr_req_desc_a_wuser_8_reg),
                                                                                               .wr_req_desc_a_wuser_9_reg(wr_req_desc_a_wuser_9_reg),
                                                                                               .wr_req_desc_a_wuser_10_reg(wr_req_desc_a_wuser_10_reg),
                                                                                               .wr_req_desc_a_wuser_11_reg(wr_req_desc_a_wuser_11_reg),
                                                                                               .wr_req_desc_a_wuser_12_reg(wr_req_desc_a_wuser_12_reg),
                                                                                               .wr_req_desc_a_wuser_13_reg(wr_req_desc_a_wuser_13_reg),
                                                                                               .wr_req_desc_a_wuser_14_reg(wr_req_desc_a_wuser_14_reg),
                                                                                               .wr_req_desc_a_wuser_15_reg(wr_req_desc_a_wuser_15_reg),
                                                                                               .wr_resp_desc_a_resp_reg(wr_resp_desc_a_resp_reg),
                                                                                               .wr_resp_desc_a_xid_0_reg(wr_resp_desc_a_xid_0_reg),
                                                                                               .wr_resp_desc_a_xid_1_reg(wr_resp_desc_a_xid_1_reg),
                                                                                               .wr_resp_desc_a_xid_2_reg(wr_resp_desc_a_xid_2_reg),
                                                                                               .wr_resp_desc_a_xid_3_reg(wr_resp_desc_a_xid_3_reg),
                                                                                               .wr_resp_desc_a_xuser_0_reg(wr_resp_desc_a_xuser_0_reg),
                                                                                               .wr_resp_desc_a_xuser_1_reg(wr_resp_desc_a_xuser_1_reg),
                                                                                               .wr_resp_desc_a_xuser_2_reg(wr_resp_desc_a_xuser_2_reg),
                                                                                               .wr_resp_desc_a_xuser_3_reg(wr_resp_desc_a_xuser_3_reg),
                                                                                               .wr_resp_desc_a_xuser_4_reg(wr_resp_desc_a_xuser_4_reg),
                                                                                               .wr_resp_desc_a_xuser_5_reg(wr_resp_desc_a_xuser_5_reg),
                                                                                               .wr_resp_desc_a_xuser_6_reg(wr_resp_desc_a_xuser_6_reg),
                                                                                               .wr_resp_desc_a_xuser_7_reg(wr_resp_desc_a_xuser_7_reg),
                                                                                               .wr_resp_desc_a_xuser_8_reg(wr_resp_desc_a_xuser_8_reg),
                                                                                               .wr_resp_desc_a_xuser_9_reg(wr_resp_desc_a_xuser_9_reg),
                                                                                               .wr_resp_desc_a_xuser_10_reg(wr_resp_desc_a_xuser_10_reg),
                                                                                               .wr_resp_desc_a_xuser_11_reg(wr_resp_desc_a_xuser_11_reg),
                                                                                               .wr_resp_desc_a_xuser_12_reg(wr_resp_desc_a_xuser_12_reg),
                                                                                               .wr_resp_desc_a_xuser_13_reg(wr_resp_desc_a_xuser_13_reg),
                                                                                               .wr_resp_desc_a_xuser_14_reg(wr_resp_desc_a_xuser_14_reg),
                                                                                               .wr_resp_desc_a_xuser_15_reg(wr_resp_desc_a_xuser_15_reg),
                                                                                               .sn_req_desc_a_attr_reg(sn_req_desc_a_attr_reg),
                                                                                               .sn_req_desc_a_acaddr_0_reg(sn_req_desc_a_acaddr_0_reg),
                                                                                               .sn_req_desc_a_acaddr_1_reg(sn_req_desc_a_acaddr_1_reg),
                                                                                               .sn_req_desc_a_acaddr_2_reg(sn_req_desc_a_acaddr_2_reg),
                                                                                               .sn_req_desc_a_acaddr_3_reg(sn_req_desc_a_acaddr_3_reg),
                                                                                               .sn_resp_desc_a_resp_reg(sn_resp_desc_a_resp_reg),
                                                                                               .rd_req_desc_b_txn_type_reg(rd_req_desc_b_txn_type_reg),
                                                                                               .rd_req_desc_b_size_reg(rd_req_desc_b_size_reg),
                                                                                               .rd_req_desc_b_axsize_reg(rd_req_desc_b_axsize_reg),
                                                                                               .rd_req_desc_b_attr_reg(rd_req_desc_b_attr_reg),
                                                                                               .rd_req_desc_b_axaddr_0_reg(rd_req_desc_b_axaddr_0_reg),
                                                                                               .rd_req_desc_b_axaddr_1_reg(rd_req_desc_b_axaddr_1_reg),
                                                                                               .rd_req_desc_b_axaddr_2_reg(rd_req_desc_b_axaddr_2_reg),
                                                                                               .rd_req_desc_b_axaddr_3_reg(rd_req_desc_b_axaddr_3_reg),
                                                                                               .rd_req_desc_b_axid_0_reg(rd_req_desc_b_axid_0_reg),
                                                                                               .rd_req_desc_b_axid_1_reg(rd_req_desc_b_axid_1_reg),
                                                                                               .rd_req_desc_b_axid_2_reg(rd_req_desc_b_axid_2_reg),
                                                                                               .rd_req_desc_b_axid_3_reg(rd_req_desc_b_axid_3_reg),
                                                                                               .rd_req_desc_b_axuser_0_reg(rd_req_desc_b_axuser_0_reg),
                                                                                               .rd_req_desc_b_axuser_1_reg(rd_req_desc_b_axuser_1_reg),
                                                                                               .rd_req_desc_b_axuser_2_reg(rd_req_desc_b_axuser_2_reg),
                                                                                               .rd_req_desc_b_axuser_3_reg(rd_req_desc_b_axuser_3_reg),
                                                                                               .rd_req_desc_b_axuser_4_reg(rd_req_desc_b_axuser_4_reg),
                                                                                               .rd_req_desc_b_axuser_5_reg(rd_req_desc_b_axuser_5_reg),
                                                                                               .rd_req_desc_b_axuser_6_reg(rd_req_desc_b_axuser_6_reg),
                                                                                               .rd_req_desc_b_axuser_7_reg(rd_req_desc_b_axuser_7_reg),
                                                                                               .rd_req_desc_b_axuser_8_reg(rd_req_desc_b_axuser_8_reg),
                                                                                               .rd_req_desc_b_axuser_9_reg(rd_req_desc_b_axuser_9_reg),
                                                                                               .rd_req_desc_b_axuser_10_reg(rd_req_desc_b_axuser_10_reg),
                                                                                               .rd_req_desc_b_axuser_11_reg(rd_req_desc_b_axuser_11_reg),
                                                                                               .rd_req_desc_b_axuser_12_reg(rd_req_desc_b_axuser_12_reg),
                                                                                               .rd_req_desc_b_axuser_13_reg(rd_req_desc_b_axuser_13_reg),
                                                                                               .rd_req_desc_b_axuser_14_reg(rd_req_desc_b_axuser_14_reg),
                                                                                               .rd_req_desc_b_axuser_15_reg(rd_req_desc_b_axuser_15_reg),
                                                                                               .rd_resp_desc_b_data_offset_reg(rd_resp_desc_b_data_offset_reg),
                                                                                               .rd_resp_desc_b_data_size_reg(rd_resp_desc_b_data_size_reg),
                                                                                               .rd_resp_desc_b_data_host_addr_0_reg(rd_resp_desc_b_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_b_data_host_addr_1_reg(rd_resp_desc_b_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_b_data_host_addr_2_reg(rd_resp_desc_b_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_b_data_host_addr_3_reg(rd_resp_desc_b_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_b_resp_reg(rd_resp_desc_b_resp_reg),
                                                                                               .rd_resp_desc_b_xid_0_reg(rd_resp_desc_b_xid_0_reg),
                                                                                               .rd_resp_desc_b_xid_1_reg(rd_resp_desc_b_xid_1_reg),
                                                                                               .rd_resp_desc_b_xid_2_reg(rd_resp_desc_b_xid_2_reg),
                                                                                               .rd_resp_desc_b_xid_3_reg(rd_resp_desc_b_xid_3_reg),
                                                                                               .rd_resp_desc_b_xuser_0_reg(rd_resp_desc_b_xuser_0_reg),
                                                                                               .rd_resp_desc_b_xuser_1_reg(rd_resp_desc_b_xuser_1_reg),
                                                                                               .rd_resp_desc_b_xuser_2_reg(rd_resp_desc_b_xuser_2_reg),
                                                                                               .rd_resp_desc_b_xuser_3_reg(rd_resp_desc_b_xuser_3_reg),
                                                                                               .rd_resp_desc_b_xuser_4_reg(rd_resp_desc_b_xuser_4_reg),
                                                                                               .rd_resp_desc_b_xuser_5_reg(rd_resp_desc_b_xuser_5_reg),
                                                                                               .rd_resp_desc_b_xuser_6_reg(rd_resp_desc_b_xuser_6_reg),
                                                                                               .rd_resp_desc_b_xuser_7_reg(rd_resp_desc_b_xuser_7_reg),
                                                                                               .rd_resp_desc_b_xuser_8_reg(rd_resp_desc_b_xuser_8_reg),
                                                                                               .rd_resp_desc_b_xuser_9_reg(rd_resp_desc_b_xuser_9_reg),
                                                                                               .rd_resp_desc_b_xuser_10_reg(rd_resp_desc_b_xuser_10_reg),
                                                                                               .rd_resp_desc_b_xuser_11_reg(rd_resp_desc_b_xuser_11_reg),
                                                                                               .rd_resp_desc_b_xuser_12_reg(rd_resp_desc_b_xuser_12_reg),
                                                                                               .rd_resp_desc_b_xuser_13_reg(rd_resp_desc_b_xuser_13_reg),
                                                                                               .rd_resp_desc_b_xuser_14_reg(rd_resp_desc_b_xuser_14_reg),
                                                                                               .rd_resp_desc_b_xuser_15_reg(rd_resp_desc_b_xuser_15_reg),
                                                                                               .wr_req_desc_b_txn_type_reg(wr_req_desc_b_txn_type_reg),
                                                                                               .wr_req_desc_b_size_reg(wr_req_desc_b_size_reg),
                                                                                               .wr_req_desc_b_data_offset_reg(wr_req_desc_b_data_offset_reg),
                                                                                               .wr_req_desc_b_data_host_addr_0_reg(wr_req_desc_b_data_host_addr_0_reg),
                                                                                               .wr_req_desc_b_data_host_addr_1_reg(wr_req_desc_b_data_host_addr_1_reg),
                                                                                               .wr_req_desc_b_data_host_addr_2_reg(wr_req_desc_b_data_host_addr_2_reg),
                                                                                               .wr_req_desc_b_data_host_addr_3_reg(wr_req_desc_b_data_host_addr_3_reg),
                                                                                               .wr_req_desc_b_wstrb_host_addr_0_reg(wr_req_desc_b_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_b_wstrb_host_addr_1_reg(wr_req_desc_b_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_b_wstrb_host_addr_2_reg(wr_req_desc_b_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_b_wstrb_host_addr_3_reg(wr_req_desc_b_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_b_axsize_reg(wr_req_desc_b_axsize_reg),
                                                                                               .wr_req_desc_b_attr_reg(wr_req_desc_b_attr_reg),
                                                                                               .wr_req_desc_b_axaddr_0_reg(wr_req_desc_b_axaddr_0_reg),
                                                                                               .wr_req_desc_b_axaddr_1_reg(wr_req_desc_b_axaddr_1_reg),
                                                                                               .wr_req_desc_b_axaddr_2_reg(wr_req_desc_b_axaddr_2_reg),
                                                                                               .wr_req_desc_b_axaddr_3_reg(wr_req_desc_b_axaddr_3_reg),
                                                                                               .wr_req_desc_b_axid_0_reg(wr_req_desc_b_axid_0_reg),
                                                                                               .wr_req_desc_b_axid_1_reg(wr_req_desc_b_axid_1_reg),
                                                                                               .wr_req_desc_b_axid_2_reg(wr_req_desc_b_axid_2_reg),
                                                                                               .wr_req_desc_b_axid_3_reg(wr_req_desc_b_axid_3_reg),
                                                                                               .wr_req_desc_b_axuser_0_reg(wr_req_desc_b_axuser_0_reg),
                                                                                               .wr_req_desc_b_axuser_1_reg(wr_req_desc_b_axuser_1_reg),
                                                                                               .wr_req_desc_b_axuser_2_reg(wr_req_desc_b_axuser_2_reg),
                                                                                               .wr_req_desc_b_axuser_3_reg(wr_req_desc_b_axuser_3_reg),
                                                                                               .wr_req_desc_b_axuser_4_reg(wr_req_desc_b_axuser_4_reg),
                                                                                               .wr_req_desc_b_axuser_5_reg(wr_req_desc_b_axuser_5_reg),
                                                                                               .wr_req_desc_b_axuser_6_reg(wr_req_desc_b_axuser_6_reg),
                                                                                               .wr_req_desc_b_axuser_7_reg(wr_req_desc_b_axuser_7_reg),
                                                                                               .wr_req_desc_b_axuser_8_reg(wr_req_desc_b_axuser_8_reg),
                                                                                               .wr_req_desc_b_axuser_9_reg(wr_req_desc_b_axuser_9_reg),
                                                                                               .wr_req_desc_b_axuser_10_reg(wr_req_desc_b_axuser_10_reg),
                                                                                               .wr_req_desc_b_axuser_11_reg(wr_req_desc_b_axuser_11_reg),
                                                                                               .wr_req_desc_b_axuser_12_reg(wr_req_desc_b_axuser_12_reg),
                                                                                               .wr_req_desc_b_axuser_13_reg(wr_req_desc_b_axuser_13_reg),
                                                                                               .wr_req_desc_b_axuser_14_reg(wr_req_desc_b_axuser_14_reg),
                                                                                               .wr_req_desc_b_axuser_15_reg(wr_req_desc_b_axuser_15_reg),
                                                                                               .wr_req_desc_b_wuser_0_reg(wr_req_desc_b_wuser_0_reg),
                                                                                               .wr_req_desc_b_wuser_1_reg(wr_req_desc_b_wuser_1_reg),
                                                                                               .wr_req_desc_b_wuser_2_reg(wr_req_desc_b_wuser_2_reg),
                                                                                               .wr_req_desc_b_wuser_3_reg(wr_req_desc_b_wuser_3_reg),
                                                                                               .wr_req_desc_b_wuser_4_reg(wr_req_desc_b_wuser_4_reg),
                                                                                               .wr_req_desc_b_wuser_5_reg(wr_req_desc_b_wuser_5_reg),
                                                                                               .wr_req_desc_b_wuser_6_reg(wr_req_desc_b_wuser_6_reg),
                                                                                               .wr_req_desc_b_wuser_7_reg(wr_req_desc_b_wuser_7_reg),
                                                                                               .wr_req_desc_b_wuser_8_reg(wr_req_desc_b_wuser_8_reg),
                                                                                               .wr_req_desc_b_wuser_9_reg(wr_req_desc_b_wuser_9_reg),
                                                                                               .wr_req_desc_b_wuser_10_reg(wr_req_desc_b_wuser_10_reg),
                                                                                               .wr_req_desc_b_wuser_11_reg(wr_req_desc_b_wuser_11_reg),
                                                                                               .wr_req_desc_b_wuser_12_reg(wr_req_desc_b_wuser_12_reg),
                                                                                               .wr_req_desc_b_wuser_13_reg(wr_req_desc_b_wuser_13_reg),
                                                                                               .wr_req_desc_b_wuser_14_reg(wr_req_desc_b_wuser_14_reg),
                                                                                               .wr_req_desc_b_wuser_15_reg(wr_req_desc_b_wuser_15_reg),
                                                                                               .wr_resp_desc_b_resp_reg(wr_resp_desc_b_resp_reg),
                                                                                               .wr_resp_desc_b_xid_0_reg(wr_resp_desc_b_xid_0_reg),
                                                                                               .wr_resp_desc_b_xid_1_reg(wr_resp_desc_b_xid_1_reg),
                                                                                               .wr_resp_desc_b_xid_2_reg(wr_resp_desc_b_xid_2_reg),
                                                                                               .wr_resp_desc_b_xid_3_reg(wr_resp_desc_b_xid_3_reg),
                                                                                               .wr_resp_desc_b_xuser_0_reg(wr_resp_desc_b_xuser_0_reg),
                                                                                               .wr_resp_desc_b_xuser_1_reg(wr_resp_desc_b_xuser_1_reg),
                                                                                               .wr_resp_desc_b_xuser_2_reg(wr_resp_desc_b_xuser_2_reg),
                                                                                               .wr_resp_desc_b_xuser_3_reg(wr_resp_desc_b_xuser_3_reg),
                                                                                               .wr_resp_desc_b_xuser_4_reg(wr_resp_desc_b_xuser_4_reg),
                                                                                               .wr_resp_desc_b_xuser_5_reg(wr_resp_desc_b_xuser_5_reg),
                                                                                               .wr_resp_desc_b_xuser_6_reg(wr_resp_desc_b_xuser_6_reg),
                                                                                               .wr_resp_desc_b_xuser_7_reg(wr_resp_desc_b_xuser_7_reg),
                                                                                               .wr_resp_desc_b_xuser_8_reg(wr_resp_desc_b_xuser_8_reg),
                                                                                               .wr_resp_desc_b_xuser_9_reg(wr_resp_desc_b_xuser_9_reg),
                                                                                               .wr_resp_desc_b_xuser_10_reg(wr_resp_desc_b_xuser_10_reg),
                                                                                               .wr_resp_desc_b_xuser_11_reg(wr_resp_desc_b_xuser_11_reg),
                                                                                               .wr_resp_desc_b_xuser_12_reg(wr_resp_desc_b_xuser_12_reg),
                                                                                               .wr_resp_desc_b_xuser_13_reg(wr_resp_desc_b_xuser_13_reg),
                                                                                               .wr_resp_desc_b_xuser_14_reg(wr_resp_desc_b_xuser_14_reg),
                                                                                               .wr_resp_desc_b_xuser_15_reg(wr_resp_desc_b_xuser_15_reg),
                                                                                               .sn_req_desc_b_attr_reg(sn_req_desc_b_attr_reg),
                                                                                               .sn_req_desc_b_acaddr_0_reg(sn_req_desc_b_acaddr_0_reg),
                                                                                               .sn_req_desc_b_acaddr_1_reg(sn_req_desc_b_acaddr_1_reg),
                                                                                               .sn_req_desc_b_acaddr_2_reg(sn_req_desc_b_acaddr_2_reg),
                                                                                               .sn_req_desc_b_acaddr_3_reg(sn_req_desc_b_acaddr_3_reg),
                                                                                               .sn_resp_desc_b_resp_reg(sn_resp_desc_b_resp_reg),
                                                                                               .rd_req_desc_c_txn_type_reg(rd_req_desc_c_txn_type_reg),
                                                                                               .rd_req_desc_c_size_reg(rd_req_desc_c_size_reg),
                                                                                               .rd_req_desc_c_axsize_reg(rd_req_desc_c_axsize_reg),
                                                                                               .rd_req_desc_c_attr_reg(rd_req_desc_c_attr_reg),
                                                                                               .rd_req_desc_c_axaddr_0_reg(rd_req_desc_c_axaddr_0_reg),
                                                                                               .rd_req_desc_c_axaddr_1_reg(rd_req_desc_c_axaddr_1_reg),
                                                                                               .rd_req_desc_c_axaddr_2_reg(rd_req_desc_c_axaddr_2_reg),
                                                                                               .rd_req_desc_c_axaddr_3_reg(rd_req_desc_c_axaddr_3_reg),
                                                                                               .rd_req_desc_c_axid_0_reg(rd_req_desc_c_axid_0_reg),
                                                                                               .rd_req_desc_c_axid_1_reg(rd_req_desc_c_axid_1_reg),
                                                                                               .rd_req_desc_c_axid_2_reg(rd_req_desc_c_axid_2_reg),
                                                                                               .rd_req_desc_c_axid_3_reg(rd_req_desc_c_axid_3_reg),
                                                                                               .rd_req_desc_c_axuser_0_reg(rd_req_desc_c_axuser_0_reg),
                                                                                               .rd_req_desc_c_axuser_1_reg(rd_req_desc_c_axuser_1_reg),
                                                                                               .rd_req_desc_c_axuser_2_reg(rd_req_desc_c_axuser_2_reg),
                                                                                               .rd_req_desc_c_axuser_3_reg(rd_req_desc_c_axuser_3_reg),
                                                                                               .rd_req_desc_c_axuser_4_reg(rd_req_desc_c_axuser_4_reg),
                                                                                               .rd_req_desc_c_axuser_5_reg(rd_req_desc_c_axuser_5_reg),
                                                                                               .rd_req_desc_c_axuser_6_reg(rd_req_desc_c_axuser_6_reg),
                                                                                               .rd_req_desc_c_axuser_7_reg(rd_req_desc_c_axuser_7_reg),
                                                                                               .rd_req_desc_c_axuser_8_reg(rd_req_desc_c_axuser_8_reg),
                                                                                               .rd_req_desc_c_axuser_9_reg(rd_req_desc_c_axuser_9_reg),
                                                                                               .rd_req_desc_c_axuser_10_reg(rd_req_desc_c_axuser_10_reg),
                                                                                               .rd_req_desc_c_axuser_11_reg(rd_req_desc_c_axuser_11_reg),
                                                                                               .rd_req_desc_c_axuser_12_reg(rd_req_desc_c_axuser_12_reg),
                                                                                               .rd_req_desc_c_axuser_13_reg(rd_req_desc_c_axuser_13_reg),
                                                                                               .rd_req_desc_c_axuser_14_reg(rd_req_desc_c_axuser_14_reg),
                                                                                               .rd_req_desc_c_axuser_15_reg(rd_req_desc_c_axuser_15_reg),
                                                                                               .rd_resp_desc_c_data_offset_reg(rd_resp_desc_c_data_offset_reg),
                                                                                               .rd_resp_desc_c_data_size_reg(rd_resp_desc_c_data_size_reg),
                                                                                               .rd_resp_desc_c_data_host_addr_0_reg(rd_resp_desc_c_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_c_data_host_addr_1_reg(rd_resp_desc_c_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_c_data_host_addr_2_reg(rd_resp_desc_c_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_c_data_host_addr_3_reg(rd_resp_desc_c_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_c_resp_reg(rd_resp_desc_c_resp_reg),
                                                                                               .rd_resp_desc_c_xid_0_reg(rd_resp_desc_c_xid_0_reg),
                                                                                               .rd_resp_desc_c_xid_1_reg(rd_resp_desc_c_xid_1_reg),
                                                                                               .rd_resp_desc_c_xid_2_reg(rd_resp_desc_c_xid_2_reg),
                                                                                               .rd_resp_desc_c_xid_3_reg(rd_resp_desc_c_xid_3_reg),
                                                                                               .rd_resp_desc_c_xuser_0_reg(rd_resp_desc_c_xuser_0_reg),
                                                                                               .rd_resp_desc_c_xuser_1_reg(rd_resp_desc_c_xuser_1_reg),
                                                                                               .rd_resp_desc_c_xuser_2_reg(rd_resp_desc_c_xuser_2_reg),
                                                                                               .rd_resp_desc_c_xuser_3_reg(rd_resp_desc_c_xuser_3_reg),
                                                                                               .rd_resp_desc_c_xuser_4_reg(rd_resp_desc_c_xuser_4_reg),
                                                                                               .rd_resp_desc_c_xuser_5_reg(rd_resp_desc_c_xuser_5_reg),
                                                                                               .rd_resp_desc_c_xuser_6_reg(rd_resp_desc_c_xuser_6_reg),
                                                                                               .rd_resp_desc_c_xuser_7_reg(rd_resp_desc_c_xuser_7_reg),
                                                                                               .rd_resp_desc_c_xuser_8_reg(rd_resp_desc_c_xuser_8_reg),
                                                                                               .rd_resp_desc_c_xuser_9_reg(rd_resp_desc_c_xuser_9_reg),
                                                                                               .rd_resp_desc_c_xuser_10_reg(rd_resp_desc_c_xuser_10_reg),
                                                                                               .rd_resp_desc_c_xuser_11_reg(rd_resp_desc_c_xuser_11_reg),
                                                                                               .rd_resp_desc_c_xuser_12_reg(rd_resp_desc_c_xuser_12_reg),
                                                                                               .rd_resp_desc_c_xuser_13_reg(rd_resp_desc_c_xuser_13_reg),
                                                                                               .rd_resp_desc_c_xuser_14_reg(rd_resp_desc_c_xuser_14_reg),
                                                                                               .rd_resp_desc_c_xuser_15_reg(rd_resp_desc_c_xuser_15_reg),
                                                                                               .wr_req_desc_c_txn_type_reg(wr_req_desc_c_txn_type_reg),
                                                                                               .wr_req_desc_c_size_reg(wr_req_desc_c_size_reg),
                                                                                               .wr_req_desc_c_data_offset_reg(wr_req_desc_c_data_offset_reg),
                                                                                               .wr_req_desc_c_data_host_addr_0_reg(wr_req_desc_c_data_host_addr_0_reg),
                                                                                               .wr_req_desc_c_data_host_addr_1_reg(wr_req_desc_c_data_host_addr_1_reg),
                                                                                               .wr_req_desc_c_data_host_addr_2_reg(wr_req_desc_c_data_host_addr_2_reg),
                                                                                               .wr_req_desc_c_data_host_addr_3_reg(wr_req_desc_c_data_host_addr_3_reg),
                                                                                               .wr_req_desc_c_wstrb_host_addr_0_reg(wr_req_desc_c_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_c_wstrb_host_addr_1_reg(wr_req_desc_c_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_c_wstrb_host_addr_2_reg(wr_req_desc_c_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_c_wstrb_host_addr_3_reg(wr_req_desc_c_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_c_axsize_reg(wr_req_desc_c_axsize_reg),
                                                                                               .wr_req_desc_c_attr_reg(wr_req_desc_c_attr_reg),
                                                                                               .wr_req_desc_c_axaddr_0_reg(wr_req_desc_c_axaddr_0_reg),
                                                                                               .wr_req_desc_c_axaddr_1_reg(wr_req_desc_c_axaddr_1_reg),
                                                                                               .wr_req_desc_c_axaddr_2_reg(wr_req_desc_c_axaddr_2_reg),
                                                                                               .wr_req_desc_c_axaddr_3_reg(wr_req_desc_c_axaddr_3_reg),
                                                                                               .wr_req_desc_c_axid_0_reg(wr_req_desc_c_axid_0_reg),
                                                                                               .wr_req_desc_c_axid_1_reg(wr_req_desc_c_axid_1_reg),
                                                                                               .wr_req_desc_c_axid_2_reg(wr_req_desc_c_axid_2_reg),
                                                                                               .wr_req_desc_c_axid_3_reg(wr_req_desc_c_axid_3_reg),
                                                                                               .wr_req_desc_c_axuser_0_reg(wr_req_desc_c_axuser_0_reg),
                                                                                               .wr_req_desc_c_axuser_1_reg(wr_req_desc_c_axuser_1_reg),
                                                                                               .wr_req_desc_c_axuser_2_reg(wr_req_desc_c_axuser_2_reg),
                                                                                               .wr_req_desc_c_axuser_3_reg(wr_req_desc_c_axuser_3_reg),
                                                                                               .wr_req_desc_c_axuser_4_reg(wr_req_desc_c_axuser_4_reg),
                                                                                               .wr_req_desc_c_axuser_5_reg(wr_req_desc_c_axuser_5_reg),
                                                                                               .wr_req_desc_c_axuser_6_reg(wr_req_desc_c_axuser_6_reg),
                                                                                               .wr_req_desc_c_axuser_7_reg(wr_req_desc_c_axuser_7_reg),
                                                                                               .wr_req_desc_c_axuser_8_reg(wr_req_desc_c_axuser_8_reg),
                                                                                               .wr_req_desc_c_axuser_9_reg(wr_req_desc_c_axuser_9_reg),
                                                                                               .wr_req_desc_c_axuser_10_reg(wr_req_desc_c_axuser_10_reg),
                                                                                               .wr_req_desc_c_axuser_11_reg(wr_req_desc_c_axuser_11_reg),
                                                                                               .wr_req_desc_c_axuser_12_reg(wr_req_desc_c_axuser_12_reg),
                                                                                               .wr_req_desc_c_axuser_13_reg(wr_req_desc_c_axuser_13_reg),
                                                                                               .wr_req_desc_c_axuser_14_reg(wr_req_desc_c_axuser_14_reg),
                                                                                               .wr_req_desc_c_axuser_15_reg(wr_req_desc_c_axuser_15_reg),
                                                                                               .wr_req_desc_c_wuser_0_reg(wr_req_desc_c_wuser_0_reg),
                                                                                               .wr_req_desc_c_wuser_1_reg(wr_req_desc_c_wuser_1_reg),
                                                                                               .wr_req_desc_c_wuser_2_reg(wr_req_desc_c_wuser_2_reg),
                                                                                               .wr_req_desc_c_wuser_3_reg(wr_req_desc_c_wuser_3_reg),
                                                                                               .wr_req_desc_c_wuser_4_reg(wr_req_desc_c_wuser_4_reg),
                                                                                               .wr_req_desc_c_wuser_5_reg(wr_req_desc_c_wuser_5_reg),
                                                                                               .wr_req_desc_c_wuser_6_reg(wr_req_desc_c_wuser_6_reg),
                                                                                               .wr_req_desc_c_wuser_7_reg(wr_req_desc_c_wuser_7_reg),
                                                                                               .wr_req_desc_c_wuser_8_reg(wr_req_desc_c_wuser_8_reg),
                                                                                               .wr_req_desc_c_wuser_9_reg(wr_req_desc_c_wuser_9_reg),
                                                                                               .wr_req_desc_c_wuser_10_reg(wr_req_desc_c_wuser_10_reg),
                                                                                               .wr_req_desc_c_wuser_11_reg(wr_req_desc_c_wuser_11_reg),
                                                                                               .wr_req_desc_c_wuser_12_reg(wr_req_desc_c_wuser_12_reg),
                                                                                               .wr_req_desc_c_wuser_13_reg(wr_req_desc_c_wuser_13_reg),
                                                                                               .wr_req_desc_c_wuser_14_reg(wr_req_desc_c_wuser_14_reg),
                                                                                               .wr_req_desc_c_wuser_15_reg(wr_req_desc_c_wuser_15_reg),
                                                                                               .wr_resp_desc_c_resp_reg(wr_resp_desc_c_resp_reg),
                                                                                               .wr_resp_desc_c_xid_0_reg(wr_resp_desc_c_xid_0_reg),
                                                                                               .wr_resp_desc_c_xid_1_reg(wr_resp_desc_c_xid_1_reg),
                                                                                               .wr_resp_desc_c_xid_2_reg(wr_resp_desc_c_xid_2_reg),
                                                                                               .wr_resp_desc_c_xid_3_reg(wr_resp_desc_c_xid_3_reg),
                                                                                               .wr_resp_desc_c_xuser_0_reg(wr_resp_desc_c_xuser_0_reg),
                                                                                               .wr_resp_desc_c_xuser_1_reg(wr_resp_desc_c_xuser_1_reg),
                                                                                               .wr_resp_desc_c_xuser_2_reg(wr_resp_desc_c_xuser_2_reg),
                                                                                               .wr_resp_desc_c_xuser_3_reg(wr_resp_desc_c_xuser_3_reg),
                                                                                               .wr_resp_desc_c_xuser_4_reg(wr_resp_desc_c_xuser_4_reg),
                                                                                               .wr_resp_desc_c_xuser_5_reg(wr_resp_desc_c_xuser_5_reg),
                                                                                               .wr_resp_desc_c_xuser_6_reg(wr_resp_desc_c_xuser_6_reg),
                                                                                               .wr_resp_desc_c_xuser_7_reg(wr_resp_desc_c_xuser_7_reg),
                                                                                               .wr_resp_desc_c_xuser_8_reg(wr_resp_desc_c_xuser_8_reg),
                                                                                               .wr_resp_desc_c_xuser_9_reg(wr_resp_desc_c_xuser_9_reg),
                                                                                               .wr_resp_desc_c_xuser_10_reg(wr_resp_desc_c_xuser_10_reg),
                                                                                               .wr_resp_desc_c_xuser_11_reg(wr_resp_desc_c_xuser_11_reg),
                                                                                               .wr_resp_desc_c_xuser_12_reg(wr_resp_desc_c_xuser_12_reg),
                                                                                               .wr_resp_desc_c_xuser_13_reg(wr_resp_desc_c_xuser_13_reg),
                                                                                               .wr_resp_desc_c_xuser_14_reg(wr_resp_desc_c_xuser_14_reg),
                                                                                               .wr_resp_desc_c_xuser_15_reg(wr_resp_desc_c_xuser_15_reg),
                                                                                               .sn_req_desc_c_attr_reg(sn_req_desc_c_attr_reg),
                                                                                               .sn_req_desc_c_acaddr_0_reg(sn_req_desc_c_acaddr_0_reg),
                                                                                               .sn_req_desc_c_acaddr_1_reg(sn_req_desc_c_acaddr_1_reg),
                                                                                               .sn_req_desc_c_acaddr_2_reg(sn_req_desc_c_acaddr_2_reg),
                                                                                               .sn_req_desc_c_acaddr_3_reg(sn_req_desc_c_acaddr_3_reg),
                                                                                               .sn_resp_desc_c_resp_reg(sn_resp_desc_c_resp_reg),
                                                                                               .rd_req_desc_d_txn_type_reg(rd_req_desc_d_txn_type_reg),
                                                                                               .rd_req_desc_d_size_reg(rd_req_desc_d_size_reg),
                                                                                               .rd_req_desc_d_axsize_reg(rd_req_desc_d_axsize_reg),
                                                                                               .rd_req_desc_d_attr_reg(rd_req_desc_d_attr_reg),
                                                                                               .rd_req_desc_d_axaddr_0_reg(rd_req_desc_d_axaddr_0_reg),
                                                                                               .rd_req_desc_d_axaddr_1_reg(rd_req_desc_d_axaddr_1_reg),
                                                                                               .rd_req_desc_d_axaddr_2_reg(rd_req_desc_d_axaddr_2_reg),
                                                                                               .rd_req_desc_d_axaddr_3_reg(rd_req_desc_d_axaddr_3_reg),
                                                                                               .rd_req_desc_d_axid_0_reg(rd_req_desc_d_axid_0_reg),
                                                                                               .rd_req_desc_d_axid_1_reg(rd_req_desc_d_axid_1_reg),
                                                                                               .rd_req_desc_d_axid_2_reg(rd_req_desc_d_axid_2_reg),
                                                                                               .rd_req_desc_d_axid_3_reg(rd_req_desc_d_axid_3_reg),
                                                                                               .rd_req_desc_d_axuser_0_reg(rd_req_desc_d_axuser_0_reg),
                                                                                               .rd_req_desc_d_axuser_1_reg(rd_req_desc_d_axuser_1_reg),
                                                                                               .rd_req_desc_d_axuser_2_reg(rd_req_desc_d_axuser_2_reg),
                                                                                               .rd_req_desc_d_axuser_3_reg(rd_req_desc_d_axuser_3_reg),
                                                                                               .rd_req_desc_d_axuser_4_reg(rd_req_desc_d_axuser_4_reg),
                                                                                               .rd_req_desc_d_axuser_5_reg(rd_req_desc_d_axuser_5_reg),
                                                                                               .rd_req_desc_d_axuser_6_reg(rd_req_desc_d_axuser_6_reg),
                                                                                               .rd_req_desc_d_axuser_7_reg(rd_req_desc_d_axuser_7_reg),
                                                                                               .rd_req_desc_d_axuser_8_reg(rd_req_desc_d_axuser_8_reg),
                                                                                               .rd_req_desc_d_axuser_9_reg(rd_req_desc_d_axuser_9_reg),
                                                                                               .rd_req_desc_d_axuser_10_reg(rd_req_desc_d_axuser_10_reg),
                                                                                               .rd_req_desc_d_axuser_11_reg(rd_req_desc_d_axuser_11_reg),
                                                                                               .rd_req_desc_d_axuser_12_reg(rd_req_desc_d_axuser_12_reg),
                                                                                               .rd_req_desc_d_axuser_13_reg(rd_req_desc_d_axuser_13_reg),
                                                                                               .rd_req_desc_d_axuser_14_reg(rd_req_desc_d_axuser_14_reg),
                                                                                               .rd_req_desc_d_axuser_15_reg(rd_req_desc_d_axuser_15_reg),
                                                                                               .rd_resp_desc_d_data_offset_reg(rd_resp_desc_d_data_offset_reg),
                                                                                               .rd_resp_desc_d_data_size_reg(rd_resp_desc_d_data_size_reg),
                                                                                               .rd_resp_desc_d_data_host_addr_0_reg(rd_resp_desc_d_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_d_data_host_addr_1_reg(rd_resp_desc_d_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_d_data_host_addr_2_reg(rd_resp_desc_d_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_d_data_host_addr_3_reg(rd_resp_desc_d_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_d_resp_reg(rd_resp_desc_d_resp_reg),
                                                                                               .rd_resp_desc_d_xid_0_reg(rd_resp_desc_d_xid_0_reg),
                                                                                               .rd_resp_desc_d_xid_1_reg(rd_resp_desc_d_xid_1_reg),
                                                                                               .rd_resp_desc_d_xid_2_reg(rd_resp_desc_d_xid_2_reg),
                                                                                               .rd_resp_desc_d_xid_3_reg(rd_resp_desc_d_xid_3_reg),
                                                                                               .rd_resp_desc_d_xuser_0_reg(rd_resp_desc_d_xuser_0_reg),
                                                                                               .rd_resp_desc_d_xuser_1_reg(rd_resp_desc_d_xuser_1_reg),
                                                                                               .rd_resp_desc_d_xuser_2_reg(rd_resp_desc_d_xuser_2_reg),
                                                                                               .rd_resp_desc_d_xuser_3_reg(rd_resp_desc_d_xuser_3_reg),
                                                                                               .rd_resp_desc_d_xuser_4_reg(rd_resp_desc_d_xuser_4_reg),
                                                                                               .rd_resp_desc_d_xuser_5_reg(rd_resp_desc_d_xuser_5_reg),
                                                                                               .rd_resp_desc_d_xuser_6_reg(rd_resp_desc_d_xuser_6_reg),
                                                                                               .rd_resp_desc_d_xuser_7_reg(rd_resp_desc_d_xuser_7_reg),
                                                                                               .rd_resp_desc_d_xuser_8_reg(rd_resp_desc_d_xuser_8_reg),
                                                                                               .rd_resp_desc_d_xuser_9_reg(rd_resp_desc_d_xuser_9_reg),
                                                                                               .rd_resp_desc_d_xuser_10_reg(rd_resp_desc_d_xuser_10_reg),
                                                                                               .rd_resp_desc_d_xuser_11_reg(rd_resp_desc_d_xuser_11_reg),
                                                                                               .rd_resp_desc_d_xuser_12_reg(rd_resp_desc_d_xuser_12_reg),
                                                                                               .rd_resp_desc_d_xuser_13_reg(rd_resp_desc_d_xuser_13_reg),
                                                                                               .rd_resp_desc_d_xuser_14_reg(rd_resp_desc_d_xuser_14_reg),
                                                                                               .rd_resp_desc_d_xuser_15_reg(rd_resp_desc_d_xuser_15_reg),
                                                                                               .wr_req_desc_d_txn_type_reg(wr_req_desc_d_txn_type_reg),
                                                                                               .wr_req_desc_d_size_reg(wr_req_desc_d_size_reg),
                                                                                               .wr_req_desc_d_data_offset_reg(wr_req_desc_d_data_offset_reg),
                                                                                               .wr_req_desc_d_data_host_addr_0_reg(wr_req_desc_d_data_host_addr_0_reg),
                                                                                               .wr_req_desc_d_data_host_addr_1_reg(wr_req_desc_d_data_host_addr_1_reg),
                                                                                               .wr_req_desc_d_data_host_addr_2_reg(wr_req_desc_d_data_host_addr_2_reg),
                                                                                               .wr_req_desc_d_data_host_addr_3_reg(wr_req_desc_d_data_host_addr_3_reg),
                                                                                               .wr_req_desc_d_wstrb_host_addr_0_reg(wr_req_desc_d_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_d_wstrb_host_addr_1_reg(wr_req_desc_d_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_d_wstrb_host_addr_2_reg(wr_req_desc_d_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_d_wstrb_host_addr_3_reg(wr_req_desc_d_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_d_axsize_reg(wr_req_desc_d_axsize_reg),
                                                                                               .wr_req_desc_d_attr_reg(wr_req_desc_d_attr_reg),
                                                                                               .wr_req_desc_d_axaddr_0_reg(wr_req_desc_d_axaddr_0_reg),
                                                                                               .wr_req_desc_d_axaddr_1_reg(wr_req_desc_d_axaddr_1_reg),
                                                                                               .wr_req_desc_d_axaddr_2_reg(wr_req_desc_d_axaddr_2_reg),
                                                                                               .wr_req_desc_d_axaddr_3_reg(wr_req_desc_d_axaddr_3_reg),
                                                                                               .wr_req_desc_d_axid_0_reg(wr_req_desc_d_axid_0_reg),
                                                                                               .wr_req_desc_d_axid_1_reg(wr_req_desc_d_axid_1_reg),
                                                                                               .wr_req_desc_d_axid_2_reg(wr_req_desc_d_axid_2_reg),
                                                                                               .wr_req_desc_d_axid_3_reg(wr_req_desc_d_axid_3_reg),
                                                                                               .wr_req_desc_d_axuser_0_reg(wr_req_desc_d_axuser_0_reg),
                                                                                               .wr_req_desc_d_axuser_1_reg(wr_req_desc_d_axuser_1_reg),
                                                                                               .wr_req_desc_d_axuser_2_reg(wr_req_desc_d_axuser_2_reg),
                                                                                               .wr_req_desc_d_axuser_3_reg(wr_req_desc_d_axuser_3_reg),
                                                                                               .wr_req_desc_d_axuser_4_reg(wr_req_desc_d_axuser_4_reg),
                                                                                               .wr_req_desc_d_axuser_5_reg(wr_req_desc_d_axuser_5_reg),
                                                                                               .wr_req_desc_d_axuser_6_reg(wr_req_desc_d_axuser_6_reg),
                                                                                               .wr_req_desc_d_axuser_7_reg(wr_req_desc_d_axuser_7_reg),
                                                                                               .wr_req_desc_d_axuser_8_reg(wr_req_desc_d_axuser_8_reg),
                                                                                               .wr_req_desc_d_axuser_9_reg(wr_req_desc_d_axuser_9_reg),
                                                                                               .wr_req_desc_d_axuser_10_reg(wr_req_desc_d_axuser_10_reg),
                                                                                               .wr_req_desc_d_axuser_11_reg(wr_req_desc_d_axuser_11_reg),
                                                                                               .wr_req_desc_d_axuser_12_reg(wr_req_desc_d_axuser_12_reg),
                                                                                               .wr_req_desc_d_axuser_13_reg(wr_req_desc_d_axuser_13_reg),
                                                                                               .wr_req_desc_d_axuser_14_reg(wr_req_desc_d_axuser_14_reg),
                                                                                               .wr_req_desc_d_axuser_15_reg(wr_req_desc_d_axuser_15_reg),
                                                                                               .wr_req_desc_d_wuser_0_reg(wr_req_desc_d_wuser_0_reg),
                                                                                               .wr_req_desc_d_wuser_1_reg(wr_req_desc_d_wuser_1_reg),
                                                                                               .wr_req_desc_d_wuser_2_reg(wr_req_desc_d_wuser_2_reg),
                                                                                               .wr_req_desc_d_wuser_3_reg(wr_req_desc_d_wuser_3_reg),
                                                                                               .wr_req_desc_d_wuser_4_reg(wr_req_desc_d_wuser_4_reg),
                                                                                               .wr_req_desc_d_wuser_5_reg(wr_req_desc_d_wuser_5_reg),
                                                                                               .wr_req_desc_d_wuser_6_reg(wr_req_desc_d_wuser_6_reg),
                                                                                               .wr_req_desc_d_wuser_7_reg(wr_req_desc_d_wuser_7_reg),
                                                                                               .wr_req_desc_d_wuser_8_reg(wr_req_desc_d_wuser_8_reg),
                                                                                               .wr_req_desc_d_wuser_9_reg(wr_req_desc_d_wuser_9_reg),
                                                                                               .wr_req_desc_d_wuser_10_reg(wr_req_desc_d_wuser_10_reg),
                                                                                               .wr_req_desc_d_wuser_11_reg(wr_req_desc_d_wuser_11_reg),
                                                                                               .wr_req_desc_d_wuser_12_reg(wr_req_desc_d_wuser_12_reg),
                                                                                               .wr_req_desc_d_wuser_13_reg(wr_req_desc_d_wuser_13_reg),
                                                                                               .wr_req_desc_d_wuser_14_reg(wr_req_desc_d_wuser_14_reg),
                                                                                               .wr_req_desc_d_wuser_15_reg(wr_req_desc_d_wuser_15_reg),
                                                                                               .wr_resp_desc_d_resp_reg(wr_resp_desc_d_resp_reg),
                                                                                               .wr_resp_desc_d_xid_0_reg(wr_resp_desc_d_xid_0_reg),
                                                                                               .wr_resp_desc_d_xid_1_reg(wr_resp_desc_d_xid_1_reg),
                                                                                               .wr_resp_desc_d_xid_2_reg(wr_resp_desc_d_xid_2_reg),
                                                                                               .wr_resp_desc_d_xid_3_reg(wr_resp_desc_d_xid_3_reg),
                                                                                               .wr_resp_desc_d_xuser_0_reg(wr_resp_desc_d_xuser_0_reg),
                                                                                               .wr_resp_desc_d_xuser_1_reg(wr_resp_desc_d_xuser_1_reg),
                                                                                               .wr_resp_desc_d_xuser_2_reg(wr_resp_desc_d_xuser_2_reg),
                                                                                               .wr_resp_desc_d_xuser_3_reg(wr_resp_desc_d_xuser_3_reg),
                                                                                               .wr_resp_desc_d_xuser_4_reg(wr_resp_desc_d_xuser_4_reg),
                                                                                               .wr_resp_desc_d_xuser_5_reg(wr_resp_desc_d_xuser_5_reg),
                                                                                               .wr_resp_desc_d_xuser_6_reg(wr_resp_desc_d_xuser_6_reg),
                                                                                               .wr_resp_desc_d_xuser_7_reg(wr_resp_desc_d_xuser_7_reg),
                                                                                               .wr_resp_desc_d_xuser_8_reg(wr_resp_desc_d_xuser_8_reg),
                                                                                               .wr_resp_desc_d_xuser_9_reg(wr_resp_desc_d_xuser_9_reg),
                                                                                               .wr_resp_desc_d_xuser_10_reg(wr_resp_desc_d_xuser_10_reg),
                                                                                               .wr_resp_desc_d_xuser_11_reg(wr_resp_desc_d_xuser_11_reg),
                                                                                               .wr_resp_desc_d_xuser_12_reg(wr_resp_desc_d_xuser_12_reg),
                                                                                               .wr_resp_desc_d_xuser_13_reg(wr_resp_desc_d_xuser_13_reg),
                                                                                               .wr_resp_desc_d_xuser_14_reg(wr_resp_desc_d_xuser_14_reg),
                                                                                               .wr_resp_desc_d_xuser_15_reg(wr_resp_desc_d_xuser_15_reg),
                                                                                               .sn_req_desc_d_attr_reg(sn_req_desc_d_attr_reg),
                                                                                               .sn_req_desc_d_acaddr_0_reg(sn_req_desc_d_acaddr_0_reg),
                                                                                               .sn_req_desc_d_acaddr_1_reg(sn_req_desc_d_acaddr_1_reg),
                                                                                               .sn_req_desc_d_acaddr_2_reg(sn_req_desc_d_acaddr_2_reg),
                                                                                               .sn_req_desc_d_acaddr_3_reg(sn_req_desc_d_acaddr_3_reg),
                                                                                               .sn_resp_desc_d_resp_reg(sn_resp_desc_d_resp_reg),
                                                                                               .rd_req_desc_e_txn_type_reg(rd_req_desc_e_txn_type_reg),
                                                                                               .rd_req_desc_e_size_reg(rd_req_desc_e_size_reg),
                                                                                               .rd_req_desc_e_axsize_reg(rd_req_desc_e_axsize_reg),
                                                                                               .rd_req_desc_e_attr_reg(rd_req_desc_e_attr_reg),
                                                                                               .rd_req_desc_e_axaddr_0_reg(rd_req_desc_e_axaddr_0_reg),
                                                                                               .rd_req_desc_e_axaddr_1_reg(rd_req_desc_e_axaddr_1_reg),
                                                                                               .rd_req_desc_e_axaddr_2_reg(rd_req_desc_e_axaddr_2_reg),
                                                                                               .rd_req_desc_e_axaddr_3_reg(rd_req_desc_e_axaddr_3_reg),
                                                                                               .rd_req_desc_e_axid_0_reg(rd_req_desc_e_axid_0_reg),
                                                                                               .rd_req_desc_e_axid_1_reg(rd_req_desc_e_axid_1_reg),
                                                                                               .rd_req_desc_e_axid_2_reg(rd_req_desc_e_axid_2_reg),
                                                                                               .rd_req_desc_e_axid_3_reg(rd_req_desc_e_axid_3_reg),
                                                                                               .rd_req_desc_e_axuser_0_reg(rd_req_desc_e_axuser_0_reg),
                                                                                               .rd_req_desc_e_axuser_1_reg(rd_req_desc_e_axuser_1_reg),
                                                                                               .rd_req_desc_e_axuser_2_reg(rd_req_desc_e_axuser_2_reg),
                                                                                               .rd_req_desc_e_axuser_3_reg(rd_req_desc_e_axuser_3_reg),
                                                                                               .rd_req_desc_e_axuser_4_reg(rd_req_desc_e_axuser_4_reg),
                                                                                               .rd_req_desc_e_axuser_5_reg(rd_req_desc_e_axuser_5_reg),
                                                                                               .rd_req_desc_e_axuser_6_reg(rd_req_desc_e_axuser_6_reg),
                                                                                               .rd_req_desc_e_axuser_7_reg(rd_req_desc_e_axuser_7_reg),
                                                                                               .rd_req_desc_e_axuser_8_reg(rd_req_desc_e_axuser_8_reg),
                                                                                               .rd_req_desc_e_axuser_9_reg(rd_req_desc_e_axuser_9_reg),
                                                                                               .rd_req_desc_e_axuser_10_reg(rd_req_desc_e_axuser_10_reg),
                                                                                               .rd_req_desc_e_axuser_11_reg(rd_req_desc_e_axuser_11_reg),
                                                                                               .rd_req_desc_e_axuser_12_reg(rd_req_desc_e_axuser_12_reg),
                                                                                               .rd_req_desc_e_axuser_13_reg(rd_req_desc_e_axuser_13_reg),
                                                                                               .rd_req_desc_e_axuser_14_reg(rd_req_desc_e_axuser_14_reg),
                                                                                               .rd_req_desc_e_axuser_15_reg(rd_req_desc_e_axuser_15_reg),
                                                                                               .rd_resp_desc_e_data_offset_reg(rd_resp_desc_e_data_offset_reg),
                                                                                               .rd_resp_desc_e_data_size_reg(rd_resp_desc_e_data_size_reg),
                                                                                               .rd_resp_desc_e_data_host_addr_0_reg(rd_resp_desc_e_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_e_data_host_addr_1_reg(rd_resp_desc_e_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_e_data_host_addr_2_reg(rd_resp_desc_e_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_e_data_host_addr_3_reg(rd_resp_desc_e_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_e_resp_reg(rd_resp_desc_e_resp_reg),
                                                                                               .rd_resp_desc_e_xid_0_reg(rd_resp_desc_e_xid_0_reg),
                                                                                               .rd_resp_desc_e_xid_1_reg(rd_resp_desc_e_xid_1_reg),
                                                                                               .rd_resp_desc_e_xid_2_reg(rd_resp_desc_e_xid_2_reg),
                                                                                               .rd_resp_desc_e_xid_3_reg(rd_resp_desc_e_xid_3_reg),
                                                                                               .rd_resp_desc_e_xuser_0_reg(rd_resp_desc_e_xuser_0_reg),
                                                                                               .rd_resp_desc_e_xuser_1_reg(rd_resp_desc_e_xuser_1_reg),
                                                                                               .rd_resp_desc_e_xuser_2_reg(rd_resp_desc_e_xuser_2_reg),
                                                                                               .rd_resp_desc_e_xuser_3_reg(rd_resp_desc_e_xuser_3_reg),
                                                                                               .rd_resp_desc_e_xuser_4_reg(rd_resp_desc_e_xuser_4_reg),
                                                                                               .rd_resp_desc_e_xuser_5_reg(rd_resp_desc_e_xuser_5_reg),
                                                                                               .rd_resp_desc_e_xuser_6_reg(rd_resp_desc_e_xuser_6_reg),
                                                                                               .rd_resp_desc_e_xuser_7_reg(rd_resp_desc_e_xuser_7_reg),
                                                                                               .rd_resp_desc_e_xuser_8_reg(rd_resp_desc_e_xuser_8_reg),
                                                                                               .rd_resp_desc_e_xuser_9_reg(rd_resp_desc_e_xuser_9_reg),
                                                                                               .rd_resp_desc_e_xuser_10_reg(rd_resp_desc_e_xuser_10_reg),
                                                                                               .rd_resp_desc_e_xuser_11_reg(rd_resp_desc_e_xuser_11_reg),
                                                                                               .rd_resp_desc_e_xuser_12_reg(rd_resp_desc_e_xuser_12_reg),
                                                                                               .rd_resp_desc_e_xuser_13_reg(rd_resp_desc_e_xuser_13_reg),
                                                                                               .rd_resp_desc_e_xuser_14_reg(rd_resp_desc_e_xuser_14_reg),
                                                                                               .rd_resp_desc_e_xuser_15_reg(rd_resp_desc_e_xuser_15_reg),
                                                                                               .wr_req_desc_e_txn_type_reg(wr_req_desc_e_txn_type_reg),
                                                                                               .wr_req_desc_e_size_reg(wr_req_desc_e_size_reg),
                                                                                               .wr_req_desc_e_data_offset_reg(wr_req_desc_e_data_offset_reg),
                                                                                               .wr_req_desc_e_data_host_addr_0_reg(wr_req_desc_e_data_host_addr_0_reg),
                                                                                               .wr_req_desc_e_data_host_addr_1_reg(wr_req_desc_e_data_host_addr_1_reg),
                                                                                               .wr_req_desc_e_data_host_addr_2_reg(wr_req_desc_e_data_host_addr_2_reg),
                                                                                               .wr_req_desc_e_data_host_addr_3_reg(wr_req_desc_e_data_host_addr_3_reg),
                                                                                               .wr_req_desc_e_wstrb_host_addr_0_reg(wr_req_desc_e_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_e_wstrb_host_addr_1_reg(wr_req_desc_e_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_e_wstrb_host_addr_2_reg(wr_req_desc_e_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_e_wstrb_host_addr_3_reg(wr_req_desc_e_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_e_axsize_reg(wr_req_desc_e_axsize_reg),
                                                                                               .wr_req_desc_e_attr_reg(wr_req_desc_e_attr_reg),
                                                                                               .wr_req_desc_e_axaddr_0_reg(wr_req_desc_e_axaddr_0_reg),
                                                                                               .wr_req_desc_e_axaddr_1_reg(wr_req_desc_e_axaddr_1_reg),
                                                                                               .wr_req_desc_e_axaddr_2_reg(wr_req_desc_e_axaddr_2_reg),
                                                                                               .wr_req_desc_e_axaddr_3_reg(wr_req_desc_e_axaddr_3_reg),
                                                                                               .wr_req_desc_e_axid_0_reg(wr_req_desc_e_axid_0_reg),
                                                                                               .wr_req_desc_e_axid_1_reg(wr_req_desc_e_axid_1_reg),
                                                                                               .wr_req_desc_e_axid_2_reg(wr_req_desc_e_axid_2_reg),
                                                                                               .wr_req_desc_e_axid_3_reg(wr_req_desc_e_axid_3_reg),
                                                                                               .wr_req_desc_e_axuser_0_reg(wr_req_desc_e_axuser_0_reg),
                                                                                               .wr_req_desc_e_axuser_1_reg(wr_req_desc_e_axuser_1_reg),
                                                                                               .wr_req_desc_e_axuser_2_reg(wr_req_desc_e_axuser_2_reg),
                                                                                               .wr_req_desc_e_axuser_3_reg(wr_req_desc_e_axuser_3_reg),
                                                                                               .wr_req_desc_e_axuser_4_reg(wr_req_desc_e_axuser_4_reg),
                                                                                               .wr_req_desc_e_axuser_5_reg(wr_req_desc_e_axuser_5_reg),
                                                                                               .wr_req_desc_e_axuser_6_reg(wr_req_desc_e_axuser_6_reg),
                                                                                               .wr_req_desc_e_axuser_7_reg(wr_req_desc_e_axuser_7_reg),
                                                                                               .wr_req_desc_e_axuser_8_reg(wr_req_desc_e_axuser_8_reg),
                                                                                               .wr_req_desc_e_axuser_9_reg(wr_req_desc_e_axuser_9_reg),
                                                                                               .wr_req_desc_e_axuser_10_reg(wr_req_desc_e_axuser_10_reg),
                                                                                               .wr_req_desc_e_axuser_11_reg(wr_req_desc_e_axuser_11_reg),
                                                                                               .wr_req_desc_e_axuser_12_reg(wr_req_desc_e_axuser_12_reg),
                                                                                               .wr_req_desc_e_axuser_13_reg(wr_req_desc_e_axuser_13_reg),
                                                                                               .wr_req_desc_e_axuser_14_reg(wr_req_desc_e_axuser_14_reg),
                                                                                               .wr_req_desc_e_axuser_15_reg(wr_req_desc_e_axuser_15_reg),
                                                                                               .wr_req_desc_e_wuser_0_reg(wr_req_desc_e_wuser_0_reg),
                                                                                               .wr_req_desc_e_wuser_1_reg(wr_req_desc_e_wuser_1_reg),
                                                                                               .wr_req_desc_e_wuser_2_reg(wr_req_desc_e_wuser_2_reg),
                                                                                               .wr_req_desc_e_wuser_3_reg(wr_req_desc_e_wuser_3_reg),
                                                                                               .wr_req_desc_e_wuser_4_reg(wr_req_desc_e_wuser_4_reg),
                                                                                               .wr_req_desc_e_wuser_5_reg(wr_req_desc_e_wuser_5_reg),
                                                                                               .wr_req_desc_e_wuser_6_reg(wr_req_desc_e_wuser_6_reg),
                                                                                               .wr_req_desc_e_wuser_7_reg(wr_req_desc_e_wuser_7_reg),
                                                                                               .wr_req_desc_e_wuser_8_reg(wr_req_desc_e_wuser_8_reg),
                                                                                               .wr_req_desc_e_wuser_9_reg(wr_req_desc_e_wuser_9_reg),
                                                                                               .wr_req_desc_e_wuser_10_reg(wr_req_desc_e_wuser_10_reg),
                                                                                               .wr_req_desc_e_wuser_11_reg(wr_req_desc_e_wuser_11_reg),
                                                                                               .wr_req_desc_e_wuser_12_reg(wr_req_desc_e_wuser_12_reg),
                                                                                               .wr_req_desc_e_wuser_13_reg(wr_req_desc_e_wuser_13_reg),
                                                                                               .wr_req_desc_e_wuser_14_reg(wr_req_desc_e_wuser_14_reg),
                                                                                               .wr_req_desc_e_wuser_15_reg(wr_req_desc_e_wuser_15_reg),
                                                                                               .wr_resp_desc_e_resp_reg(wr_resp_desc_e_resp_reg),
                                                                                               .wr_resp_desc_e_xid_0_reg(wr_resp_desc_e_xid_0_reg),
                                                                                               .wr_resp_desc_e_xid_1_reg(wr_resp_desc_e_xid_1_reg),
                                                                                               .wr_resp_desc_e_xid_2_reg(wr_resp_desc_e_xid_2_reg),
                                                                                               .wr_resp_desc_e_xid_3_reg(wr_resp_desc_e_xid_3_reg),
                                                                                               .wr_resp_desc_e_xuser_0_reg(wr_resp_desc_e_xuser_0_reg),
                                                                                               .wr_resp_desc_e_xuser_1_reg(wr_resp_desc_e_xuser_1_reg),
                                                                                               .wr_resp_desc_e_xuser_2_reg(wr_resp_desc_e_xuser_2_reg),
                                                                                               .wr_resp_desc_e_xuser_3_reg(wr_resp_desc_e_xuser_3_reg),
                                                                                               .wr_resp_desc_e_xuser_4_reg(wr_resp_desc_e_xuser_4_reg),
                                                                                               .wr_resp_desc_e_xuser_5_reg(wr_resp_desc_e_xuser_5_reg),
                                                                                               .wr_resp_desc_e_xuser_6_reg(wr_resp_desc_e_xuser_6_reg),
                                                                                               .wr_resp_desc_e_xuser_7_reg(wr_resp_desc_e_xuser_7_reg),
                                                                                               .wr_resp_desc_e_xuser_8_reg(wr_resp_desc_e_xuser_8_reg),
                                                                                               .wr_resp_desc_e_xuser_9_reg(wr_resp_desc_e_xuser_9_reg),
                                                                                               .wr_resp_desc_e_xuser_10_reg(wr_resp_desc_e_xuser_10_reg),
                                                                                               .wr_resp_desc_e_xuser_11_reg(wr_resp_desc_e_xuser_11_reg),
                                                                                               .wr_resp_desc_e_xuser_12_reg(wr_resp_desc_e_xuser_12_reg),
                                                                                               .wr_resp_desc_e_xuser_13_reg(wr_resp_desc_e_xuser_13_reg),
                                                                                               .wr_resp_desc_e_xuser_14_reg(wr_resp_desc_e_xuser_14_reg),
                                                                                               .wr_resp_desc_e_xuser_15_reg(wr_resp_desc_e_xuser_15_reg),
                                                                                               .sn_req_desc_e_attr_reg(sn_req_desc_e_attr_reg),
                                                                                               .sn_req_desc_e_acaddr_0_reg(sn_req_desc_e_acaddr_0_reg),
                                                                                               .sn_req_desc_e_acaddr_1_reg(sn_req_desc_e_acaddr_1_reg),
                                                                                               .sn_req_desc_e_acaddr_2_reg(sn_req_desc_e_acaddr_2_reg),
                                                                                               .sn_req_desc_e_acaddr_3_reg(sn_req_desc_e_acaddr_3_reg),
                                                                                               .sn_resp_desc_e_resp_reg(sn_resp_desc_e_resp_reg),
                                                                                               .rd_req_desc_f_txn_type_reg(rd_req_desc_f_txn_type_reg),
                                                                                               .rd_req_desc_f_size_reg(rd_req_desc_f_size_reg),
                                                                                               .rd_req_desc_f_axsize_reg(rd_req_desc_f_axsize_reg),
                                                                                               .rd_req_desc_f_attr_reg(rd_req_desc_f_attr_reg),
                                                                                               .rd_req_desc_f_axaddr_0_reg(rd_req_desc_f_axaddr_0_reg),
                                                                                               .rd_req_desc_f_axaddr_1_reg(rd_req_desc_f_axaddr_1_reg),
                                                                                               .rd_req_desc_f_axaddr_2_reg(rd_req_desc_f_axaddr_2_reg),
                                                                                               .rd_req_desc_f_axaddr_3_reg(rd_req_desc_f_axaddr_3_reg),
                                                                                               .rd_req_desc_f_axid_0_reg(rd_req_desc_f_axid_0_reg),
                                                                                               .rd_req_desc_f_axid_1_reg(rd_req_desc_f_axid_1_reg),
                                                                                               .rd_req_desc_f_axid_2_reg(rd_req_desc_f_axid_2_reg),
                                                                                               .rd_req_desc_f_axid_3_reg(rd_req_desc_f_axid_3_reg),
                                                                                               .rd_req_desc_f_axuser_0_reg(rd_req_desc_f_axuser_0_reg),
                                                                                               .rd_req_desc_f_axuser_1_reg(rd_req_desc_f_axuser_1_reg),
                                                                                               .rd_req_desc_f_axuser_2_reg(rd_req_desc_f_axuser_2_reg),
                                                                                               .rd_req_desc_f_axuser_3_reg(rd_req_desc_f_axuser_3_reg),
                                                                                               .rd_req_desc_f_axuser_4_reg(rd_req_desc_f_axuser_4_reg),
                                                                                               .rd_req_desc_f_axuser_5_reg(rd_req_desc_f_axuser_5_reg),
                                                                                               .rd_req_desc_f_axuser_6_reg(rd_req_desc_f_axuser_6_reg),
                                                                                               .rd_req_desc_f_axuser_7_reg(rd_req_desc_f_axuser_7_reg),
                                                                                               .rd_req_desc_f_axuser_8_reg(rd_req_desc_f_axuser_8_reg),
                                                                                               .rd_req_desc_f_axuser_9_reg(rd_req_desc_f_axuser_9_reg),
                                                                                               .rd_req_desc_f_axuser_10_reg(rd_req_desc_f_axuser_10_reg),
                                                                                               .rd_req_desc_f_axuser_11_reg(rd_req_desc_f_axuser_11_reg),
                                                                                               .rd_req_desc_f_axuser_12_reg(rd_req_desc_f_axuser_12_reg),
                                                                                               .rd_req_desc_f_axuser_13_reg(rd_req_desc_f_axuser_13_reg),
                                                                                               .rd_req_desc_f_axuser_14_reg(rd_req_desc_f_axuser_14_reg),
                                                                                               .rd_req_desc_f_axuser_15_reg(rd_req_desc_f_axuser_15_reg),
                                                                                               .rd_resp_desc_f_data_offset_reg(rd_resp_desc_f_data_offset_reg),
                                                                                               .rd_resp_desc_f_data_size_reg(rd_resp_desc_f_data_size_reg),
                                                                                               .rd_resp_desc_f_data_host_addr_0_reg(rd_resp_desc_f_data_host_addr_0_reg),
                                                                                               .rd_resp_desc_f_data_host_addr_1_reg(rd_resp_desc_f_data_host_addr_1_reg),
                                                                                               .rd_resp_desc_f_data_host_addr_2_reg(rd_resp_desc_f_data_host_addr_2_reg),
                                                                                               .rd_resp_desc_f_data_host_addr_3_reg(rd_resp_desc_f_data_host_addr_3_reg),
                                                                                               .rd_resp_desc_f_resp_reg(rd_resp_desc_f_resp_reg),
                                                                                               .rd_resp_desc_f_xid_0_reg(rd_resp_desc_f_xid_0_reg),
                                                                                               .rd_resp_desc_f_xid_1_reg(rd_resp_desc_f_xid_1_reg),
                                                                                               .rd_resp_desc_f_xid_2_reg(rd_resp_desc_f_xid_2_reg),
                                                                                               .rd_resp_desc_f_xid_3_reg(rd_resp_desc_f_xid_3_reg),
                                                                                               .rd_resp_desc_f_xuser_0_reg(rd_resp_desc_f_xuser_0_reg),
                                                                                               .rd_resp_desc_f_xuser_1_reg(rd_resp_desc_f_xuser_1_reg),
                                                                                               .rd_resp_desc_f_xuser_2_reg(rd_resp_desc_f_xuser_2_reg),
                                                                                               .rd_resp_desc_f_xuser_3_reg(rd_resp_desc_f_xuser_3_reg),
                                                                                               .rd_resp_desc_f_xuser_4_reg(rd_resp_desc_f_xuser_4_reg),
                                                                                               .rd_resp_desc_f_xuser_5_reg(rd_resp_desc_f_xuser_5_reg),
                                                                                               .rd_resp_desc_f_xuser_6_reg(rd_resp_desc_f_xuser_6_reg),
                                                                                               .rd_resp_desc_f_xuser_7_reg(rd_resp_desc_f_xuser_7_reg),
                                                                                               .rd_resp_desc_f_xuser_8_reg(rd_resp_desc_f_xuser_8_reg),
                                                                                               .rd_resp_desc_f_xuser_9_reg(rd_resp_desc_f_xuser_9_reg),
                                                                                               .rd_resp_desc_f_xuser_10_reg(rd_resp_desc_f_xuser_10_reg),
                                                                                               .rd_resp_desc_f_xuser_11_reg(rd_resp_desc_f_xuser_11_reg),
                                                                                               .rd_resp_desc_f_xuser_12_reg(rd_resp_desc_f_xuser_12_reg),
                                                                                               .rd_resp_desc_f_xuser_13_reg(rd_resp_desc_f_xuser_13_reg),
                                                                                               .rd_resp_desc_f_xuser_14_reg(rd_resp_desc_f_xuser_14_reg),
                                                                                               .rd_resp_desc_f_xuser_15_reg(rd_resp_desc_f_xuser_15_reg),
                                                                                               .wr_req_desc_f_txn_type_reg(wr_req_desc_f_txn_type_reg),
                                                                                               .wr_req_desc_f_size_reg(wr_req_desc_f_size_reg),
                                                                                               .wr_req_desc_f_data_offset_reg(wr_req_desc_f_data_offset_reg),
                                                                                               .wr_req_desc_f_data_host_addr_0_reg(wr_req_desc_f_data_host_addr_0_reg),
                                                                                               .wr_req_desc_f_data_host_addr_1_reg(wr_req_desc_f_data_host_addr_1_reg),
                                                                                               .wr_req_desc_f_data_host_addr_2_reg(wr_req_desc_f_data_host_addr_2_reg),
                                                                                               .wr_req_desc_f_data_host_addr_3_reg(wr_req_desc_f_data_host_addr_3_reg),
                                                                                               .wr_req_desc_f_wstrb_host_addr_0_reg(wr_req_desc_f_wstrb_host_addr_0_reg),
                                                                                               .wr_req_desc_f_wstrb_host_addr_1_reg(wr_req_desc_f_wstrb_host_addr_1_reg),
                                                                                               .wr_req_desc_f_wstrb_host_addr_2_reg(wr_req_desc_f_wstrb_host_addr_2_reg),
                                                                                               .wr_req_desc_f_wstrb_host_addr_3_reg(wr_req_desc_f_wstrb_host_addr_3_reg),
                                                                                               .wr_req_desc_f_axsize_reg(wr_req_desc_f_axsize_reg),
                                                                                               .wr_req_desc_f_attr_reg(wr_req_desc_f_attr_reg),
                                                                                               .wr_req_desc_f_axaddr_0_reg(wr_req_desc_f_axaddr_0_reg),
                                                                                               .wr_req_desc_f_axaddr_1_reg(wr_req_desc_f_axaddr_1_reg),
                                                                                               .wr_req_desc_f_axaddr_2_reg(wr_req_desc_f_axaddr_2_reg),
                                                                                               .wr_req_desc_f_axaddr_3_reg(wr_req_desc_f_axaddr_3_reg),
                                                                                               .wr_req_desc_f_axid_0_reg(wr_req_desc_f_axid_0_reg),
                                                                                               .wr_req_desc_f_axid_1_reg(wr_req_desc_f_axid_1_reg),
                                                                                               .wr_req_desc_f_axid_2_reg(wr_req_desc_f_axid_2_reg),
                                                                                               .wr_req_desc_f_axid_3_reg(wr_req_desc_f_axid_3_reg),
                                                                                               .wr_req_desc_f_axuser_0_reg(wr_req_desc_f_axuser_0_reg),
                                                                                               .wr_req_desc_f_axuser_1_reg(wr_req_desc_f_axuser_1_reg),
                                                                                               .wr_req_desc_f_axuser_2_reg(wr_req_desc_f_axuser_2_reg),
                                                                                               .wr_req_desc_f_axuser_3_reg(wr_req_desc_f_axuser_3_reg),
                                                                                               .wr_req_desc_f_axuser_4_reg(wr_req_desc_f_axuser_4_reg),
                                                                                               .wr_req_desc_f_axuser_5_reg(wr_req_desc_f_axuser_5_reg),
                                                                                               .wr_req_desc_f_axuser_6_reg(wr_req_desc_f_axuser_6_reg),
                                                                                               .wr_req_desc_f_axuser_7_reg(wr_req_desc_f_axuser_7_reg),
                                                                                               .wr_req_desc_f_axuser_8_reg(wr_req_desc_f_axuser_8_reg),
                                                                                               .wr_req_desc_f_axuser_9_reg(wr_req_desc_f_axuser_9_reg),
                                                                                               .wr_req_desc_f_axuser_10_reg(wr_req_desc_f_axuser_10_reg),
                                                                                               .wr_req_desc_f_axuser_11_reg(wr_req_desc_f_axuser_11_reg),
                                                                                               .wr_req_desc_f_axuser_12_reg(wr_req_desc_f_axuser_12_reg),
                                                                                               .wr_req_desc_f_axuser_13_reg(wr_req_desc_f_axuser_13_reg),
                                                                                               .wr_req_desc_f_axuser_14_reg(wr_req_desc_f_axuser_14_reg),
                                                                                               .wr_req_desc_f_axuser_15_reg(wr_req_desc_f_axuser_15_reg),
                                                                                               .wr_req_desc_f_wuser_0_reg(wr_req_desc_f_wuser_0_reg),
                                                                                               .wr_req_desc_f_wuser_1_reg(wr_req_desc_f_wuser_1_reg),
                                                                                               .wr_req_desc_f_wuser_2_reg(wr_req_desc_f_wuser_2_reg),
                                                                                               .wr_req_desc_f_wuser_3_reg(wr_req_desc_f_wuser_3_reg),
                                                                                               .wr_req_desc_f_wuser_4_reg(wr_req_desc_f_wuser_4_reg),
                                                                                               .wr_req_desc_f_wuser_5_reg(wr_req_desc_f_wuser_5_reg),
                                                                                               .wr_req_desc_f_wuser_6_reg(wr_req_desc_f_wuser_6_reg),
                                                                                               .wr_req_desc_f_wuser_7_reg(wr_req_desc_f_wuser_7_reg),
                                                                                               .wr_req_desc_f_wuser_8_reg(wr_req_desc_f_wuser_8_reg),
                                                                                               .wr_req_desc_f_wuser_9_reg(wr_req_desc_f_wuser_9_reg),
                                                                                               .wr_req_desc_f_wuser_10_reg(wr_req_desc_f_wuser_10_reg),
                                                                                               .wr_req_desc_f_wuser_11_reg(wr_req_desc_f_wuser_11_reg),
                                                                                               .wr_req_desc_f_wuser_12_reg(wr_req_desc_f_wuser_12_reg),
                                                                                               .wr_req_desc_f_wuser_13_reg(wr_req_desc_f_wuser_13_reg),
                                                                                               .wr_req_desc_f_wuser_14_reg(wr_req_desc_f_wuser_14_reg),
                                                                                               .wr_req_desc_f_wuser_15_reg(wr_req_desc_f_wuser_15_reg),
                                                                                               .wr_resp_desc_f_resp_reg(wr_resp_desc_f_resp_reg),
                                                                                               .wr_resp_desc_f_xid_0_reg(wr_resp_desc_f_xid_0_reg),
                                                                                               .wr_resp_desc_f_xid_1_reg(wr_resp_desc_f_xid_1_reg),
                                                                                               .wr_resp_desc_f_xid_2_reg(wr_resp_desc_f_xid_2_reg),
                                                                                               .wr_resp_desc_f_xid_3_reg(wr_resp_desc_f_xid_3_reg),
                                                                                               .wr_resp_desc_f_xuser_0_reg(wr_resp_desc_f_xuser_0_reg),
                                                                                               .wr_resp_desc_f_xuser_1_reg(wr_resp_desc_f_xuser_1_reg),
                                                                                               .wr_resp_desc_f_xuser_2_reg(wr_resp_desc_f_xuser_2_reg),
                                                                                               .wr_resp_desc_f_xuser_3_reg(wr_resp_desc_f_xuser_3_reg),
                                                                                               .wr_resp_desc_f_xuser_4_reg(wr_resp_desc_f_xuser_4_reg),
                                                                                               .wr_resp_desc_f_xuser_5_reg(wr_resp_desc_f_xuser_5_reg),
                                                                                               .wr_resp_desc_f_xuser_6_reg(wr_resp_desc_f_xuser_6_reg),
                                                                                               .wr_resp_desc_f_xuser_7_reg(wr_resp_desc_f_xuser_7_reg),
                                                                                               .wr_resp_desc_f_xuser_8_reg(wr_resp_desc_f_xuser_8_reg),
                                                                                               .wr_resp_desc_f_xuser_9_reg(wr_resp_desc_f_xuser_9_reg),
                                                                                               .wr_resp_desc_f_xuser_10_reg(wr_resp_desc_f_xuser_10_reg),
                                                                                               .wr_resp_desc_f_xuser_11_reg(wr_resp_desc_f_xuser_11_reg),
                                                                                               .wr_resp_desc_f_xuser_12_reg(wr_resp_desc_f_xuser_12_reg),
                                                                                               .wr_resp_desc_f_xuser_13_reg(wr_resp_desc_f_xuser_13_reg),
                                                                                               .wr_resp_desc_f_xuser_14_reg(wr_resp_desc_f_xuser_14_reg),
                                                                                               .wr_resp_desc_f_xuser_15_reg(wr_resp_desc_f_xuser_15_reg),
                                                                                               .sn_req_desc_f_attr_reg(sn_req_desc_f_attr_reg),
                                                                                               .sn_req_desc_f_acaddr_0_reg(sn_req_desc_f_acaddr_0_reg),
                                                                                               .sn_req_desc_f_acaddr_1_reg(sn_req_desc_f_acaddr_1_reg),
                                                                                               .sn_req_desc_f_acaddr_2_reg(sn_req_desc_f_acaddr_2_reg),
                                                                                               .sn_req_desc_f_acaddr_3_reg(sn_req_desc_f_acaddr_3_reg),
                                                                                               .sn_resp_desc_f_resp_reg(sn_resp_desc_f_resp_reg),
                                                                                               .rb2uc_rd_data      (rb2uc_rd_data),
                                                                                               .rb2uc_rd_wstrb     (rb2uc_rd_wstrb),
                                                                                               .rb2uc_sn_data      (rb2uc_sn_data),
                                                                                               .rd_hm2uc_done      (rd_hm2uc_done),
                                                                                               .wr_hm2uc_done      (wr_hm2uc_done),
                                                                                               .rd_resp_fifo_pop_desc_conn(rd_resp_fifo_pop_desc_conn),
                                                                                               .wr_resp_fifo_pop_desc_conn(wr_resp_fifo_pop_desc_conn),
                                                                                               .sn_req_fifo_pop_desc_conn(sn_req_fifo_pop_desc_conn));

endmodule

// Local Variables:
// verilog-library-directories:("./")
// End:

