/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */
                       
assign int_desc_0_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[0];
assign int_desc_0_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[0];
assign int_desc_0_attr_axregion = int_desc_n_attr_axregion[0];
assign int_desc_0_attr_axqos = int_desc_n_attr_axqos[0];
assign int_desc_0_attr_axprot = int_desc_n_attr_axprot[0];
assign int_desc_0_attr_axcache = int_desc_n_attr_axcache[0];
assign int_desc_0_attr_axlock = int_desc_n_attr_axlock[0];
assign int_desc_0_attr_axburst = int_desc_n_attr_axburst[0];
assign int_desc_0_axid_0_axid = int_desc_n_axid_0_axid[0];
assign int_desc_0_axid_1_axid = int_desc_n_axid_1_axid[0];
assign int_desc_0_axid_2_axid = int_desc_n_axid_2_axid[0];
assign int_desc_0_axid_3_axid = int_desc_n_axid_3_axid[0];
assign int_desc_0_axuser_0_axuser = int_desc_n_axuser_0_axuser[0];
assign int_desc_0_axuser_1_axuser = int_desc_n_axuser_1_axuser[0];
assign int_desc_0_axuser_2_axuser = int_desc_n_axuser_2_axuser[0];
assign int_desc_0_axuser_3_axuser = int_desc_n_axuser_3_axuser[0];
assign int_desc_0_axuser_4_axuser = int_desc_n_axuser_4_axuser[0];
assign int_desc_0_axuser_5_axuser = int_desc_n_axuser_5_axuser[0];
assign int_desc_0_axuser_6_axuser = int_desc_n_axuser_6_axuser[0];
assign int_desc_0_axuser_7_axuser = int_desc_n_axuser_7_axuser[0];
assign int_desc_0_axuser_8_axuser = int_desc_n_axuser_8_axuser[0];
assign int_desc_0_axuser_9_axuser = int_desc_n_axuser_9_axuser[0];
assign int_desc_0_axuser_10_axuser = int_desc_n_axuser_10_axuser[0];
assign int_desc_0_axuser_11_axuser = int_desc_n_axuser_11_axuser[0];
assign int_desc_0_axuser_12_axuser = int_desc_n_axuser_12_axuser[0];
assign int_desc_0_axuser_13_axuser = int_desc_n_axuser_13_axuser[0];
assign int_desc_0_axuser_14_axuser = int_desc_n_axuser_14_axuser[0];
assign int_desc_0_axuser_15_axuser = int_desc_n_axuser_15_axuser[0];
assign int_desc_0_size_txn_size = int_desc_n_size_txn_size[0];
assign int_desc_0_axsize_axsize = int_desc_n_axsize_axsize[0];
assign int_desc_0_axaddr_0_addr = int_desc_n_axaddr_0_addr[0];
assign int_desc_0_axaddr_1_addr = int_desc_n_axaddr_1_addr[0];
assign int_desc_0_axaddr_2_addr = int_desc_n_axaddr_2_addr[0];
assign int_desc_0_axaddr_3_addr = int_desc_n_axaddr_3_addr[0];
assign int_desc_0_data_offset_addr = int_desc_n_data_offset_addr[0];
assign int_desc_0_wuser_0_wuser = int_desc_n_wuser_0_wuser[0];
assign int_desc_0_wuser_1_wuser = int_desc_n_wuser_1_wuser[0];
assign int_desc_0_wuser_2_wuser = int_desc_n_wuser_2_wuser[0];
assign int_desc_0_wuser_3_wuser = int_desc_n_wuser_3_wuser[0];
assign int_desc_0_wuser_4_wuser = int_desc_n_wuser_4_wuser[0];
assign int_desc_0_wuser_5_wuser = int_desc_n_wuser_5_wuser[0];
assign int_desc_0_wuser_6_wuser = int_desc_n_wuser_6_wuser[0];
assign int_desc_0_wuser_7_wuser = int_desc_n_wuser_7_wuser[0];
assign int_desc_0_wuser_8_wuser = int_desc_n_wuser_8_wuser[0];
assign int_desc_0_wuser_9_wuser = int_desc_n_wuser_9_wuser[0];
assign int_desc_0_wuser_10_wuser = int_desc_n_wuser_10_wuser[0];
assign int_desc_0_wuser_11_wuser = int_desc_n_wuser_11_wuser[0];
assign int_desc_0_wuser_12_wuser = int_desc_n_wuser_12_wuser[0];
assign int_desc_0_wuser_13_wuser = int_desc_n_wuser_13_wuser[0];
assign int_desc_0_wuser_14_wuser = int_desc_n_wuser_14_wuser[0];
assign int_desc_0_wuser_15_wuser = int_desc_n_wuser_15_wuser[0];
assign int_desc_1_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[1];
assign int_desc_1_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[1];
assign int_desc_1_attr_axregion = int_desc_n_attr_axregion[1];
assign int_desc_1_attr_axqos = int_desc_n_attr_axqos[1];
assign int_desc_1_attr_axprot = int_desc_n_attr_axprot[1];
assign int_desc_1_attr_axcache = int_desc_n_attr_axcache[1];
assign int_desc_1_attr_axlock = int_desc_n_attr_axlock[1];
assign int_desc_1_attr_axburst = int_desc_n_attr_axburst[1];
assign int_desc_1_axid_0_axid = int_desc_n_axid_0_axid[1];
assign int_desc_1_axid_1_axid = int_desc_n_axid_1_axid[1];
assign int_desc_1_axid_2_axid = int_desc_n_axid_2_axid[1];
assign int_desc_1_axid_3_axid = int_desc_n_axid_3_axid[1];
assign int_desc_1_axuser_0_axuser = int_desc_n_axuser_0_axuser[1];
assign int_desc_1_axuser_1_axuser = int_desc_n_axuser_1_axuser[1];
assign int_desc_1_axuser_2_axuser = int_desc_n_axuser_2_axuser[1];
assign int_desc_1_axuser_3_axuser = int_desc_n_axuser_3_axuser[1];
assign int_desc_1_axuser_4_axuser = int_desc_n_axuser_4_axuser[1];
assign int_desc_1_axuser_5_axuser = int_desc_n_axuser_5_axuser[1];
assign int_desc_1_axuser_6_axuser = int_desc_n_axuser_6_axuser[1];
assign int_desc_1_axuser_7_axuser = int_desc_n_axuser_7_axuser[1];
assign int_desc_1_axuser_8_axuser = int_desc_n_axuser_8_axuser[1];
assign int_desc_1_axuser_9_axuser = int_desc_n_axuser_9_axuser[1];
assign int_desc_1_axuser_10_axuser = int_desc_n_axuser_10_axuser[1];
assign int_desc_1_axuser_11_axuser = int_desc_n_axuser_11_axuser[1];
assign int_desc_1_axuser_12_axuser = int_desc_n_axuser_12_axuser[1];
assign int_desc_1_axuser_13_axuser = int_desc_n_axuser_13_axuser[1];
assign int_desc_1_axuser_14_axuser = int_desc_n_axuser_14_axuser[1];
assign int_desc_1_axuser_15_axuser = int_desc_n_axuser_15_axuser[1];
assign int_desc_1_size_txn_size = int_desc_n_size_txn_size[1];
assign int_desc_1_axsize_axsize = int_desc_n_axsize_axsize[1];
assign int_desc_1_axaddr_0_addr = int_desc_n_axaddr_0_addr[1];
assign int_desc_1_axaddr_1_addr = int_desc_n_axaddr_1_addr[1];
assign int_desc_1_axaddr_2_addr = int_desc_n_axaddr_2_addr[1];
assign int_desc_1_axaddr_3_addr = int_desc_n_axaddr_3_addr[1];
assign int_desc_1_data_offset_addr = int_desc_n_data_offset_addr[1];
assign int_desc_1_wuser_0_wuser = int_desc_n_wuser_0_wuser[1];
assign int_desc_1_wuser_1_wuser = int_desc_n_wuser_1_wuser[1];
assign int_desc_1_wuser_2_wuser = int_desc_n_wuser_2_wuser[1];
assign int_desc_1_wuser_3_wuser = int_desc_n_wuser_3_wuser[1];
assign int_desc_1_wuser_4_wuser = int_desc_n_wuser_4_wuser[1];
assign int_desc_1_wuser_5_wuser = int_desc_n_wuser_5_wuser[1];
assign int_desc_1_wuser_6_wuser = int_desc_n_wuser_6_wuser[1];
assign int_desc_1_wuser_7_wuser = int_desc_n_wuser_7_wuser[1];
assign int_desc_1_wuser_8_wuser = int_desc_n_wuser_8_wuser[1];
assign int_desc_1_wuser_9_wuser = int_desc_n_wuser_9_wuser[1];
assign int_desc_1_wuser_10_wuser = int_desc_n_wuser_10_wuser[1];
assign int_desc_1_wuser_11_wuser = int_desc_n_wuser_11_wuser[1];
assign int_desc_1_wuser_12_wuser = int_desc_n_wuser_12_wuser[1];
assign int_desc_1_wuser_13_wuser = int_desc_n_wuser_13_wuser[1];
assign int_desc_1_wuser_14_wuser = int_desc_n_wuser_14_wuser[1];
assign int_desc_1_wuser_15_wuser = int_desc_n_wuser_15_wuser[1];
assign int_desc_2_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[2];
assign int_desc_2_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[2];
assign int_desc_2_attr_axregion = int_desc_n_attr_axregion[2];
assign int_desc_2_attr_axqos = int_desc_n_attr_axqos[2];
assign int_desc_2_attr_axprot = int_desc_n_attr_axprot[2];
assign int_desc_2_attr_axcache = int_desc_n_attr_axcache[2];
assign int_desc_2_attr_axlock = int_desc_n_attr_axlock[2];
assign int_desc_2_attr_axburst = int_desc_n_attr_axburst[2];
assign int_desc_2_axid_0_axid = int_desc_n_axid_0_axid[2];
assign int_desc_2_axid_1_axid = int_desc_n_axid_1_axid[2];
assign int_desc_2_axid_2_axid = int_desc_n_axid_2_axid[2];
assign int_desc_2_axid_3_axid = int_desc_n_axid_3_axid[2];
assign int_desc_2_axuser_0_axuser = int_desc_n_axuser_0_axuser[2];
assign int_desc_2_axuser_1_axuser = int_desc_n_axuser_1_axuser[2];
assign int_desc_2_axuser_2_axuser = int_desc_n_axuser_2_axuser[2];
assign int_desc_2_axuser_3_axuser = int_desc_n_axuser_3_axuser[2];
assign int_desc_2_axuser_4_axuser = int_desc_n_axuser_4_axuser[2];
assign int_desc_2_axuser_5_axuser = int_desc_n_axuser_5_axuser[2];
assign int_desc_2_axuser_6_axuser = int_desc_n_axuser_6_axuser[2];
assign int_desc_2_axuser_7_axuser = int_desc_n_axuser_7_axuser[2];
assign int_desc_2_axuser_8_axuser = int_desc_n_axuser_8_axuser[2];
assign int_desc_2_axuser_9_axuser = int_desc_n_axuser_9_axuser[2];
assign int_desc_2_axuser_10_axuser = int_desc_n_axuser_10_axuser[2];
assign int_desc_2_axuser_11_axuser = int_desc_n_axuser_11_axuser[2];
assign int_desc_2_axuser_12_axuser = int_desc_n_axuser_12_axuser[2];
assign int_desc_2_axuser_13_axuser = int_desc_n_axuser_13_axuser[2];
assign int_desc_2_axuser_14_axuser = int_desc_n_axuser_14_axuser[2];
assign int_desc_2_axuser_15_axuser = int_desc_n_axuser_15_axuser[2];
assign int_desc_2_size_txn_size = int_desc_n_size_txn_size[2];
assign int_desc_2_axsize_axsize = int_desc_n_axsize_axsize[2];
assign int_desc_2_axaddr_0_addr = int_desc_n_axaddr_0_addr[2];
assign int_desc_2_axaddr_1_addr = int_desc_n_axaddr_1_addr[2];
assign int_desc_2_axaddr_2_addr = int_desc_n_axaddr_2_addr[2];
assign int_desc_2_axaddr_3_addr = int_desc_n_axaddr_3_addr[2];
assign int_desc_2_data_offset_addr = int_desc_n_data_offset_addr[2];
assign int_desc_2_wuser_0_wuser = int_desc_n_wuser_0_wuser[2];
assign int_desc_2_wuser_1_wuser = int_desc_n_wuser_1_wuser[2];
assign int_desc_2_wuser_2_wuser = int_desc_n_wuser_2_wuser[2];
assign int_desc_2_wuser_3_wuser = int_desc_n_wuser_3_wuser[2];
assign int_desc_2_wuser_4_wuser = int_desc_n_wuser_4_wuser[2];
assign int_desc_2_wuser_5_wuser = int_desc_n_wuser_5_wuser[2];
assign int_desc_2_wuser_6_wuser = int_desc_n_wuser_6_wuser[2];
assign int_desc_2_wuser_7_wuser = int_desc_n_wuser_7_wuser[2];
assign int_desc_2_wuser_8_wuser = int_desc_n_wuser_8_wuser[2];
assign int_desc_2_wuser_9_wuser = int_desc_n_wuser_9_wuser[2];
assign int_desc_2_wuser_10_wuser = int_desc_n_wuser_10_wuser[2];
assign int_desc_2_wuser_11_wuser = int_desc_n_wuser_11_wuser[2];
assign int_desc_2_wuser_12_wuser = int_desc_n_wuser_12_wuser[2];
assign int_desc_2_wuser_13_wuser = int_desc_n_wuser_13_wuser[2];
assign int_desc_2_wuser_14_wuser = int_desc_n_wuser_14_wuser[2];
assign int_desc_2_wuser_15_wuser = int_desc_n_wuser_15_wuser[2];
assign int_desc_3_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[3];
assign int_desc_3_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[3];
assign int_desc_3_attr_axregion = int_desc_n_attr_axregion[3];
assign int_desc_3_attr_axqos = int_desc_n_attr_axqos[3];
assign int_desc_3_attr_axprot = int_desc_n_attr_axprot[3];
assign int_desc_3_attr_axcache = int_desc_n_attr_axcache[3];
assign int_desc_3_attr_axlock = int_desc_n_attr_axlock[3];
assign int_desc_3_attr_axburst = int_desc_n_attr_axburst[3];
assign int_desc_3_axid_0_axid = int_desc_n_axid_0_axid[3];
assign int_desc_3_axid_1_axid = int_desc_n_axid_1_axid[3];
assign int_desc_3_axid_2_axid = int_desc_n_axid_2_axid[3];
assign int_desc_3_axid_3_axid = int_desc_n_axid_3_axid[3];
assign int_desc_3_axuser_0_axuser = int_desc_n_axuser_0_axuser[3];
assign int_desc_3_axuser_1_axuser = int_desc_n_axuser_1_axuser[3];
assign int_desc_3_axuser_2_axuser = int_desc_n_axuser_2_axuser[3];
assign int_desc_3_axuser_3_axuser = int_desc_n_axuser_3_axuser[3];
assign int_desc_3_axuser_4_axuser = int_desc_n_axuser_4_axuser[3];
assign int_desc_3_axuser_5_axuser = int_desc_n_axuser_5_axuser[3];
assign int_desc_3_axuser_6_axuser = int_desc_n_axuser_6_axuser[3];
assign int_desc_3_axuser_7_axuser = int_desc_n_axuser_7_axuser[3];
assign int_desc_3_axuser_8_axuser = int_desc_n_axuser_8_axuser[3];
assign int_desc_3_axuser_9_axuser = int_desc_n_axuser_9_axuser[3];
assign int_desc_3_axuser_10_axuser = int_desc_n_axuser_10_axuser[3];
assign int_desc_3_axuser_11_axuser = int_desc_n_axuser_11_axuser[3];
assign int_desc_3_axuser_12_axuser = int_desc_n_axuser_12_axuser[3];
assign int_desc_3_axuser_13_axuser = int_desc_n_axuser_13_axuser[3];
assign int_desc_3_axuser_14_axuser = int_desc_n_axuser_14_axuser[3];
assign int_desc_3_axuser_15_axuser = int_desc_n_axuser_15_axuser[3];
assign int_desc_3_size_txn_size = int_desc_n_size_txn_size[3];
assign int_desc_3_axsize_axsize = int_desc_n_axsize_axsize[3];
assign int_desc_3_axaddr_0_addr = int_desc_n_axaddr_0_addr[3];
assign int_desc_3_axaddr_1_addr = int_desc_n_axaddr_1_addr[3];
assign int_desc_3_axaddr_2_addr = int_desc_n_axaddr_2_addr[3];
assign int_desc_3_axaddr_3_addr = int_desc_n_axaddr_3_addr[3];
assign int_desc_3_data_offset_addr = int_desc_n_data_offset_addr[3];
assign int_desc_3_wuser_0_wuser = int_desc_n_wuser_0_wuser[3];
assign int_desc_3_wuser_1_wuser = int_desc_n_wuser_1_wuser[3];
assign int_desc_3_wuser_2_wuser = int_desc_n_wuser_2_wuser[3];
assign int_desc_3_wuser_3_wuser = int_desc_n_wuser_3_wuser[3];
assign int_desc_3_wuser_4_wuser = int_desc_n_wuser_4_wuser[3];
assign int_desc_3_wuser_5_wuser = int_desc_n_wuser_5_wuser[3];
assign int_desc_3_wuser_6_wuser = int_desc_n_wuser_6_wuser[3];
assign int_desc_3_wuser_7_wuser = int_desc_n_wuser_7_wuser[3];
assign int_desc_3_wuser_8_wuser = int_desc_n_wuser_8_wuser[3];
assign int_desc_3_wuser_9_wuser = int_desc_n_wuser_9_wuser[3];
assign int_desc_3_wuser_10_wuser = int_desc_n_wuser_10_wuser[3];
assign int_desc_3_wuser_11_wuser = int_desc_n_wuser_11_wuser[3];
assign int_desc_3_wuser_12_wuser = int_desc_n_wuser_12_wuser[3];
assign int_desc_3_wuser_13_wuser = int_desc_n_wuser_13_wuser[3];
assign int_desc_3_wuser_14_wuser = int_desc_n_wuser_14_wuser[3];
assign int_desc_3_wuser_15_wuser = int_desc_n_wuser_15_wuser[3];
assign int_desc_4_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[4];
assign int_desc_4_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[4];
assign int_desc_4_attr_axregion = int_desc_n_attr_axregion[4];
assign int_desc_4_attr_axqos = int_desc_n_attr_axqos[4];
assign int_desc_4_attr_axprot = int_desc_n_attr_axprot[4];
assign int_desc_4_attr_axcache = int_desc_n_attr_axcache[4];
assign int_desc_4_attr_axlock = int_desc_n_attr_axlock[4];
assign int_desc_4_attr_axburst = int_desc_n_attr_axburst[4];
assign int_desc_4_axid_0_axid = int_desc_n_axid_0_axid[4];
assign int_desc_4_axid_1_axid = int_desc_n_axid_1_axid[4];
assign int_desc_4_axid_2_axid = int_desc_n_axid_2_axid[4];
assign int_desc_4_axid_3_axid = int_desc_n_axid_3_axid[4];
assign int_desc_4_axuser_0_axuser = int_desc_n_axuser_0_axuser[4];
assign int_desc_4_axuser_1_axuser = int_desc_n_axuser_1_axuser[4];
assign int_desc_4_axuser_2_axuser = int_desc_n_axuser_2_axuser[4];
assign int_desc_4_axuser_3_axuser = int_desc_n_axuser_3_axuser[4];
assign int_desc_4_axuser_4_axuser = int_desc_n_axuser_4_axuser[4];
assign int_desc_4_axuser_5_axuser = int_desc_n_axuser_5_axuser[4];
assign int_desc_4_axuser_6_axuser = int_desc_n_axuser_6_axuser[4];
assign int_desc_4_axuser_7_axuser = int_desc_n_axuser_7_axuser[4];
assign int_desc_4_axuser_8_axuser = int_desc_n_axuser_8_axuser[4];
assign int_desc_4_axuser_9_axuser = int_desc_n_axuser_9_axuser[4];
assign int_desc_4_axuser_10_axuser = int_desc_n_axuser_10_axuser[4];
assign int_desc_4_axuser_11_axuser = int_desc_n_axuser_11_axuser[4];
assign int_desc_4_axuser_12_axuser = int_desc_n_axuser_12_axuser[4];
assign int_desc_4_axuser_13_axuser = int_desc_n_axuser_13_axuser[4];
assign int_desc_4_axuser_14_axuser = int_desc_n_axuser_14_axuser[4];
assign int_desc_4_axuser_15_axuser = int_desc_n_axuser_15_axuser[4];
assign int_desc_4_size_txn_size = int_desc_n_size_txn_size[4];
assign int_desc_4_axsize_axsize = int_desc_n_axsize_axsize[4];
assign int_desc_4_axaddr_0_addr = int_desc_n_axaddr_0_addr[4];
assign int_desc_4_axaddr_1_addr = int_desc_n_axaddr_1_addr[4];
assign int_desc_4_axaddr_2_addr = int_desc_n_axaddr_2_addr[4];
assign int_desc_4_axaddr_3_addr = int_desc_n_axaddr_3_addr[4];
assign int_desc_4_data_offset_addr = int_desc_n_data_offset_addr[4];
assign int_desc_4_wuser_0_wuser = int_desc_n_wuser_0_wuser[4];
assign int_desc_4_wuser_1_wuser = int_desc_n_wuser_1_wuser[4];
assign int_desc_4_wuser_2_wuser = int_desc_n_wuser_2_wuser[4];
assign int_desc_4_wuser_3_wuser = int_desc_n_wuser_3_wuser[4];
assign int_desc_4_wuser_4_wuser = int_desc_n_wuser_4_wuser[4];
assign int_desc_4_wuser_5_wuser = int_desc_n_wuser_5_wuser[4];
assign int_desc_4_wuser_6_wuser = int_desc_n_wuser_6_wuser[4];
assign int_desc_4_wuser_7_wuser = int_desc_n_wuser_7_wuser[4];
assign int_desc_4_wuser_8_wuser = int_desc_n_wuser_8_wuser[4];
assign int_desc_4_wuser_9_wuser = int_desc_n_wuser_9_wuser[4];
assign int_desc_4_wuser_10_wuser = int_desc_n_wuser_10_wuser[4];
assign int_desc_4_wuser_11_wuser = int_desc_n_wuser_11_wuser[4];
assign int_desc_4_wuser_12_wuser = int_desc_n_wuser_12_wuser[4];
assign int_desc_4_wuser_13_wuser = int_desc_n_wuser_13_wuser[4];
assign int_desc_4_wuser_14_wuser = int_desc_n_wuser_14_wuser[4];
assign int_desc_4_wuser_15_wuser = int_desc_n_wuser_15_wuser[4];
assign int_desc_5_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[5];
assign int_desc_5_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[5];
assign int_desc_5_attr_axregion = int_desc_n_attr_axregion[5];
assign int_desc_5_attr_axqos = int_desc_n_attr_axqos[5];
assign int_desc_5_attr_axprot = int_desc_n_attr_axprot[5];
assign int_desc_5_attr_axcache = int_desc_n_attr_axcache[5];
assign int_desc_5_attr_axlock = int_desc_n_attr_axlock[5];
assign int_desc_5_attr_axburst = int_desc_n_attr_axburst[5];
assign int_desc_5_axid_0_axid = int_desc_n_axid_0_axid[5];
assign int_desc_5_axid_1_axid = int_desc_n_axid_1_axid[5];
assign int_desc_5_axid_2_axid = int_desc_n_axid_2_axid[5];
assign int_desc_5_axid_3_axid = int_desc_n_axid_3_axid[5];
assign int_desc_5_axuser_0_axuser = int_desc_n_axuser_0_axuser[5];
assign int_desc_5_axuser_1_axuser = int_desc_n_axuser_1_axuser[5];
assign int_desc_5_axuser_2_axuser = int_desc_n_axuser_2_axuser[5];
assign int_desc_5_axuser_3_axuser = int_desc_n_axuser_3_axuser[5];
assign int_desc_5_axuser_4_axuser = int_desc_n_axuser_4_axuser[5];
assign int_desc_5_axuser_5_axuser = int_desc_n_axuser_5_axuser[5];
assign int_desc_5_axuser_6_axuser = int_desc_n_axuser_6_axuser[5];
assign int_desc_5_axuser_7_axuser = int_desc_n_axuser_7_axuser[5];
assign int_desc_5_axuser_8_axuser = int_desc_n_axuser_8_axuser[5];
assign int_desc_5_axuser_9_axuser = int_desc_n_axuser_9_axuser[5];
assign int_desc_5_axuser_10_axuser = int_desc_n_axuser_10_axuser[5];
assign int_desc_5_axuser_11_axuser = int_desc_n_axuser_11_axuser[5];
assign int_desc_5_axuser_12_axuser = int_desc_n_axuser_12_axuser[5];
assign int_desc_5_axuser_13_axuser = int_desc_n_axuser_13_axuser[5];
assign int_desc_5_axuser_14_axuser = int_desc_n_axuser_14_axuser[5];
assign int_desc_5_axuser_15_axuser = int_desc_n_axuser_15_axuser[5];
assign int_desc_5_size_txn_size = int_desc_n_size_txn_size[5];
assign int_desc_5_axsize_axsize = int_desc_n_axsize_axsize[5];
assign int_desc_5_axaddr_0_addr = int_desc_n_axaddr_0_addr[5];
assign int_desc_5_axaddr_1_addr = int_desc_n_axaddr_1_addr[5];
assign int_desc_5_axaddr_2_addr = int_desc_n_axaddr_2_addr[5];
assign int_desc_5_axaddr_3_addr = int_desc_n_axaddr_3_addr[5];
assign int_desc_5_data_offset_addr = int_desc_n_data_offset_addr[5];
assign int_desc_5_wuser_0_wuser = int_desc_n_wuser_0_wuser[5];
assign int_desc_5_wuser_1_wuser = int_desc_n_wuser_1_wuser[5];
assign int_desc_5_wuser_2_wuser = int_desc_n_wuser_2_wuser[5];
assign int_desc_5_wuser_3_wuser = int_desc_n_wuser_3_wuser[5];
assign int_desc_5_wuser_4_wuser = int_desc_n_wuser_4_wuser[5];
assign int_desc_5_wuser_5_wuser = int_desc_n_wuser_5_wuser[5];
assign int_desc_5_wuser_6_wuser = int_desc_n_wuser_6_wuser[5];
assign int_desc_5_wuser_7_wuser = int_desc_n_wuser_7_wuser[5];
assign int_desc_5_wuser_8_wuser = int_desc_n_wuser_8_wuser[5];
assign int_desc_5_wuser_9_wuser = int_desc_n_wuser_9_wuser[5];
assign int_desc_5_wuser_10_wuser = int_desc_n_wuser_10_wuser[5];
assign int_desc_5_wuser_11_wuser = int_desc_n_wuser_11_wuser[5];
assign int_desc_5_wuser_12_wuser = int_desc_n_wuser_12_wuser[5];
assign int_desc_5_wuser_13_wuser = int_desc_n_wuser_13_wuser[5];
assign int_desc_5_wuser_14_wuser = int_desc_n_wuser_14_wuser[5];
assign int_desc_5_wuser_15_wuser = int_desc_n_wuser_15_wuser[5];
assign int_desc_6_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[6];
assign int_desc_6_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[6];
assign int_desc_6_attr_axregion = int_desc_n_attr_axregion[6];
assign int_desc_6_attr_axqos = int_desc_n_attr_axqos[6];
assign int_desc_6_attr_axprot = int_desc_n_attr_axprot[6];
assign int_desc_6_attr_axcache = int_desc_n_attr_axcache[6];
assign int_desc_6_attr_axlock = int_desc_n_attr_axlock[6];
assign int_desc_6_attr_axburst = int_desc_n_attr_axburst[6];
assign int_desc_6_axid_0_axid = int_desc_n_axid_0_axid[6];
assign int_desc_6_axid_1_axid = int_desc_n_axid_1_axid[6];
assign int_desc_6_axid_2_axid = int_desc_n_axid_2_axid[6];
assign int_desc_6_axid_3_axid = int_desc_n_axid_3_axid[6];
assign int_desc_6_axuser_0_axuser = int_desc_n_axuser_0_axuser[6];
assign int_desc_6_axuser_1_axuser = int_desc_n_axuser_1_axuser[6];
assign int_desc_6_axuser_2_axuser = int_desc_n_axuser_2_axuser[6];
assign int_desc_6_axuser_3_axuser = int_desc_n_axuser_3_axuser[6];
assign int_desc_6_axuser_4_axuser = int_desc_n_axuser_4_axuser[6];
assign int_desc_6_axuser_5_axuser = int_desc_n_axuser_5_axuser[6];
assign int_desc_6_axuser_6_axuser = int_desc_n_axuser_6_axuser[6];
assign int_desc_6_axuser_7_axuser = int_desc_n_axuser_7_axuser[6];
assign int_desc_6_axuser_8_axuser = int_desc_n_axuser_8_axuser[6];
assign int_desc_6_axuser_9_axuser = int_desc_n_axuser_9_axuser[6];
assign int_desc_6_axuser_10_axuser = int_desc_n_axuser_10_axuser[6];
assign int_desc_6_axuser_11_axuser = int_desc_n_axuser_11_axuser[6];
assign int_desc_6_axuser_12_axuser = int_desc_n_axuser_12_axuser[6];
assign int_desc_6_axuser_13_axuser = int_desc_n_axuser_13_axuser[6];
assign int_desc_6_axuser_14_axuser = int_desc_n_axuser_14_axuser[6];
assign int_desc_6_axuser_15_axuser = int_desc_n_axuser_15_axuser[6];
assign int_desc_6_size_txn_size = int_desc_n_size_txn_size[6];
assign int_desc_6_axsize_axsize = int_desc_n_axsize_axsize[6];
assign int_desc_6_axaddr_0_addr = int_desc_n_axaddr_0_addr[6];
assign int_desc_6_axaddr_1_addr = int_desc_n_axaddr_1_addr[6];
assign int_desc_6_axaddr_2_addr = int_desc_n_axaddr_2_addr[6];
assign int_desc_6_axaddr_3_addr = int_desc_n_axaddr_3_addr[6];
assign int_desc_6_data_offset_addr = int_desc_n_data_offset_addr[6];
assign int_desc_6_wuser_0_wuser = int_desc_n_wuser_0_wuser[6];
assign int_desc_6_wuser_1_wuser = int_desc_n_wuser_1_wuser[6];
assign int_desc_6_wuser_2_wuser = int_desc_n_wuser_2_wuser[6];
assign int_desc_6_wuser_3_wuser = int_desc_n_wuser_3_wuser[6];
assign int_desc_6_wuser_4_wuser = int_desc_n_wuser_4_wuser[6];
assign int_desc_6_wuser_5_wuser = int_desc_n_wuser_5_wuser[6];
assign int_desc_6_wuser_6_wuser = int_desc_n_wuser_6_wuser[6];
assign int_desc_6_wuser_7_wuser = int_desc_n_wuser_7_wuser[6];
assign int_desc_6_wuser_8_wuser = int_desc_n_wuser_8_wuser[6];
assign int_desc_6_wuser_9_wuser = int_desc_n_wuser_9_wuser[6];
assign int_desc_6_wuser_10_wuser = int_desc_n_wuser_10_wuser[6];
assign int_desc_6_wuser_11_wuser = int_desc_n_wuser_11_wuser[6];
assign int_desc_6_wuser_12_wuser = int_desc_n_wuser_12_wuser[6];
assign int_desc_6_wuser_13_wuser = int_desc_n_wuser_13_wuser[6];
assign int_desc_6_wuser_14_wuser = int_desc_n_wuser_14_wuser[6];
assign int_desc_6_wuser_15_wuser = int_desc_n_wuser_15_wuser[6];
assign int_desc_7_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[7];
assign int_desc_7_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[7];
assign int_desc_7_attr_axregion = int_desc_n_attr_axregion[7];
assign int_desc_7_attr_axqos = int_desc_n_attr_axqos[7];
assign int_desc_7_attr_axprot = int_desc_n_attr_axprot[7];
assign int_desc_7_attr_axcache = int_desc_n_attr_axcache[7];
assign int_desc_7_attr_axlock = int_desc_n_attr_axlock[7];
assign int_desc_7_attr_axburst = int_desc_n_attr_axburst[7];
assign int_desc_7_axid_0_axid = int_desc_n_axid_0_axid[7];
assign int_desc_7_axid_1_axid = int_desc_n_axid_1_axid[7];
assign int_desc_7_axid_2_axid = int_desc_n_axid_2_axid[7];
assign int_desc_7_axid_3_axid = int_desc_n_axid_3_axid[7];
assign int_desc_7_axuser_0_axuser = int_desc_n_axuser_0_axuser[7];
assign int_desc_7_axuser_1_axuser = int_desc_n_axuser_1_axuser[7];
assign int_desc_7_axuser_2_axuser = int_desc_n_axuser_2_axuser[7];
assign int_desc_7_axuser_3_axuser = int_desc_n_axuser_3_axuser[7];
assign int_desc_7_axuser_4_axuser = int_desc_n_axuser_4_axuser[7];
assign int_desc_7_axuser_5_axuser = int_desc_n_axuser_5_axuser[7];
assign int_desc_7_axuser_6_axuser = int_desc_n_axuser_6_axuser[7];
assign int_desc_7_axuser_7_axuser = int_desc_n_axuser_7_axuser[7];
assign int_desc_7_axuser_8_axuser = int_desc_n_axuser_8_axuser[7];
assign int_desc_7_axuser_9_axuser = int_desc_n_axuser_9_axuser[7];
assign int_desc_7_axuser_10_axuser = int_desc_n_axuser_10_axuser[7];
assign int_desc_7_axuser_11_axuser = int_desc_n_axuser_11_axuser[7];
assign int_desc_7_axuser_12_axuser = int_desc_n_axuser_12_axuser[7];
assign int_desc_7_axuser_13_axuser = int_desc_n_axuser_13_axuser[7];
assign int_desc_7_axuser_14_axuser = int_desc_n_axuser_14_axuser[7];
assign int_desc_7_axuser_15_axuser = int_desc_n_axuser_15_axuser[7];
assign int_desc_7_size_txn_size = int_desc_n_size_txn_size[7];
assign int_desc_7_axsize_axsize = int_desc_n_axsize_axsize[7];
assign int_desc_7_axaddr_0_addr = int_desc_n_axaddr_0_addr[7];
assign int_desc_7_axaddr_1_addr = int_desc_n_axaddr_1_addr[7];
assign int_desc_7_axaddr_2_addr = int_desc_n_axaddr_2_addr[7];
assign int_desc_7_axaddr_3_addr = int_desc_n_axaddr_3_addr[7];
assign int_desc_7_data_offset_addr = int_desc_n_data_offset_addr[7];
assign int_desc_7_wuser_0_wuser = int_desc_n_wuser_0_wuser[7];
assign int_desc_7_wuser_1_wuser = int_desc_n_wuser_1_wuser[7];
assign int_desc_7_wuser_2_wuser = int_desc_n_wuser_2_wuser[7];
assign int_desc_7_wuser_3_wuser = int_desc_n_wuser_3_wuser[7];
assign int_desc_7_wuser_4_wuser = int_desc_n_wuser_4_wuser[7];
assign int_desc_7_wuser_5_wuser = int_desc_n_wuser_5_wuser[7];
assign int_desc_7_wuser_6_wuser = int_desc_n_wuser_6_wuser[7];
assign int_desc_7_wuser_7_wuser = int_desc_n_wuser_7_wuser[7];
assign int_desc_7_wuser_8_wuser = int_desc_n_wuser_8_wuser[7];
assign int_desc_7_wuser_9_wuser = int_desc_n_wuser_9_wuser[7];
assign int_desc_7_wuser_10_wuser = int_desc_n_wuser_10_wuser[7];
assign int_desc_7_wuser_11_wuser = int_desc_n_wuser_11_wuser[7];
assign int_desc_7_wuser_12_wuser = int_desc_n_wuser_12_wuser[7];
assign int_desc_7_wuser_13_wuser = int_desc_n_wuser_13_wuser[7];
assign int_desc_7_wuser_14_wuser = int_desc_n_wuser_14_wuser[7];
assign int_desc_7_wuser_15_wuser = int_desc_n_wuser_15_wuser[7];
assign int_desc_8_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[8];
assign int_desc_8_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[8];
assign int_desc_8_attr_axregion = int_desc_n_attr_axregion[8];
assign int_desc_8_attr_axqos = int_desc_n_attr_axqos[8];
assign int_desc_8_attr_axprot = int_desc_n_attr_axprot[8];
assign int_desc_8_attr_axcache = int_desc_n_attr_axcache[8];
assign int_desc_8_attr_axlock = int_desc_n_attr_axlock[8];
assign int_desc_8_attr_axburst = int_desc_n_attr_axburst[8];
assign int_desc_8_axid_0_axid = int_desc_n_axid_0_axid[8];
assign int_desc_8_axid_1_axid = int_desc_n_axid_1_axid[8];
assign int_desc_8_axid_2_axid = int_desc_n_axid_2_axid[8];
assign int_desc_8_axid_3_axid = int_desc_n_axid_3_axid[8];
assign int_desc_8_axuser_0_axuser = int_desc_n_axuser_0_axuser[8];
assign int_desc_8_axuser_1_axuser = int_desc_n_axuser_1_axuser[8];
assign int_desc_8_axuser_2_axuser = int_desc_n_axuser_2_axuser[8];
assign int_desc_8_axuser_3_axuser = int_desc_n_axuser_3_axuser[8];
assign int_desc_8_axuser_4_axuser = int_desc_n_axuser_4_axuser[8];
assign int_desc_8_axuser_5_axuser = int_desc_n_axuser_5_axuser[8];
assign int_desc_8_axuser_6_axuser = int_desc_n_axuser_6_axuser[8];
assign int_desc_8_axuser_7_axuser = int_desc_n_axuser_7_axuser[8];
assign int_desc_8_axuser_8_axuser = int_desc_n_axuser_8_axuser[8];
assign int_desc_8_axuser_9_axuser = int_desc_n_axuser_9_axuser[8];
assign int_desc_8_axuser_10_axuser = int_desc_n_axuser_10_axuser[8];
assign int_desc_8_axuser_11_axuser = int_desc_n_axuser_11_axuser[8];
assign int_desc_8_axuser_12_axuser = int_desc_n_axuser_12_axuser[8];
assign int_desc_8_axuser_13_axuser = int_desc_n_axuser_13_axuser[8];
assign int_desc_8_axuser_14_axuser = int_desc_n_axuser_14_axuser[8];
assign int_desc_8_axuser_15_axuser = int_desc_n_axuser_15_axuser[8];
assign int_desc_8_size_txn_size = int_desc_n_size_txn_size[8];
assign int_desc_8_axsize_axsize = int_desc_n_axsize_axsize[8];
assign int_desc_8_axaddr_0_addr = int_desc_n_axaddr_0_addr[8];
assign int_desc_8_axaddr_1_addr = int_desc_n_axaddr_1_addr[8];
assign int_desc_8_axaddr_2_addr = int_desc_n_axaddr_2_addr[8];
assign int_desc_8_axaddr_3_addr = int_desc_n_axaddr_3_addr[8];
assign int_desc_8_data_offset_addr = int_desc_n_data_offset_addr[8];
assign int_desc_8_wuser_0_wuser = int_desc_n_wuser_0_wuser[8];
assign int_desc_8_wuser_1_wuser = int_desc_n_wuser_1_wuser[8];
assign int_desc_8_wuser_2_wuser = int_desc_n_wuser_2_wuser[8];
assign int_desc_8_wuser_3_wuser = int_desc_n_wuser_3_wuser[8];
assign int_desc_8_wuser_4_wuser = int_desc_n_wuser_4_wuser[8];
assign int_desc_8_wuser_5_wuser = int_desc_n_wuser_5_wuser[8];
assign int_desc_8_wuser_6_wuser = int_desc_n_wuser_6_wuser[8];
assign int_desc_8_wuser_7_wuser = int_desc_n_wuser_7_wuser[8];
assign int_desc_8_wuser_8_wuser = int_desc_n_wuser_8_wuser[8];
assign int_desc_8_wuser_9_wuser = int_desc_n_wuser_9_wuser[8];
assign int_desc_8_wuser_10_wuser = int_desc_n_wuser_10_wuser[8];
assign int_desc_8_wuser_11_wuser = int_desc_n_wuser_11_wuser[8];
assign int_desc_8_wuser_12_wuser = int_desc_n_wuser_12_wuser[8];
assign int_desc_8_wuser_13_wuser = int_desc_n_wuser_13_wuser[8];
assign int_desc_8_wuser_14_wuser = int_desc_n_wuser_14_wuser[8];
assign int_desc_8_wuser_15_wuser = int_desc_n_wuser_15_wuser[8];
assign int_desc_9_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[9];
assign int_desc_9_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[9];
assign int_desc_9_attr_axregion = int_desc_n_attr_axregion[9];
assign int_desc_9_attr_axqos = int_desc_n_attr_axqos[9];
assign int_desc_9_attr_axprot = int_desc_n_attr_axprot[9];
assign int_desc_9_attr_axcache = int_desc_n_attr_axcache[9];
assign int_desc_9_attr_axlock = int_desc_n_attr_axlock[9];
assign int_desc_9_attr_axburst = int_desc_n_attr_axburst[9];
assign int_desc_9_axid_0_axid = int_desc_n_axid_0_axid[9];
assign int_desc_9_axid_1_axid = int_desc_n_axid_1_axid[9];
assign int_desc_9_axid_2_axid = int_desc_n_axid_2_axid[9];
assign int_desc_9_axid_3_axid = int_desc_n_axid_3_axid[9];
assign int_desc_9_axuser_0_axuser = int_desc_n_axuser_0_axuser[9];
assign int_desc_9_axuser_1_axuser = int_desc_n_axuser_1_axuser[9];
assign int_desc_9_axuser_2_axuser = int_desc_n_axuser_2_axuser[9];
assign int_desc_9_axuser_3_axuser = int_desc_n_axuser_3_axuser[9];
assign int_desc_9_axuser_4_axuser = int_desc_n_axuser_4_axuser[9];
assign int_desc_9_axuser_5_axuser = int_desc_n_axuser_5_axuser[9];
assign int_desc_9_axuser_6_axuser = int_desc_n_axuser_6_axuser[9];
assign int_desc_9_axuser_7_axuser = int_desc_n_axuser_7_axuser[9];
assign int_desc_9_axuser_8_axuser = int_desc_n_axuser_8_axuser[9];
assign int_desc_9_axuser_9_axuser = int_desc_n_axuser_9_axuser[9];
assign int_desc_9_axuser_10_axuser = int_desc_n_axuser_10_axuser[9];
assign int_desc_9_axuser_11_axuser = int_desc_n_axuser_11_axuser[9];
assign int_desc_9_axuser_12_axuser = int_desc_n_axuser_12_axuser[9];
assign int_desc_9_axuser_13_axuser = int_desc_n_axuser_13_axuser[9];
assign int_desc_9_axuser_14_axuser = int_desc_n_axuser_14_axuser[9];
assign int_desc_9_axuser_15_axuser = int_desc_n_axuser_15_axuser[9];
assign int_desc_9_size_txn_size = int_desc_n_size_txn_size[9];
assign int_desc_9_axsize_axsize = int_desc_n_axsize_axsize[9];
assign int_desc_9_axaddr_0_addr = int_desc_n_axaddr_0_addr[9];
assign int_desc_9_axaddr_1_addr = int_desc_n_axaddr_1_addr[9];
assign int_desc_9_axaddr_2_addr = int_desc_n_axaddr_2_addr[9];
assign int_desc_9_axaddr_3_addr = int_desc_n_axaddr_3_addr[9];
assign int_desc_9_data_offset_addr = int_desc_n_data_offset_addr[9];
assign int_desc_9_wuser_0_wuser = int_desc_n_wuser_0_wuser[9];
assign int_desc_9_wuser_1_wuser = int_desc_n_wuser_1_wuser[9];
assign int_desc_9_wuser_2_wuser = int_desc_n_wuser_2_wuser[9];
assign int_desc_9_wuser_3_wuser = int_desc_n_wuser_3_wuser[9];
assign int_desc_9_wuser_4_wuser = int_desc_n_wuser_4_wuser[9];
assign int_desc_9_wuser_5_wuser = int_desc_n_wuser_5_wuser[9];
assign int_desc_9_wuser_6_wuser = int_desc_n_wuser_6_wuser[9];
assign int_desc_9_wuser_7_wuser = int_desc_n_wuser_7_wuser[9];
assign int_desc_9_wuser_8_wuser = int_desc_n_wuser_8_wuser[9];
assign int_desc_9_wuser_9_wuser = int_desc_n_wuser_9_wuser[9];
assign int_desc_9_wuser_10_wuser = int_desc_n_wuser_10_wuser[9];
assign int_desc_9_wuser_11_wuser = int_desc_n_wuser_11_wuser[9];
assign int_desc_9_wuser_12_wuser = int_desc_n_wuser_12_wuser[9];
assign int_desc_9_wuser_13_wuser = int_desc_n_wuser_13_wuser[9];
assign int_desc_9_wuser_14_wuser = int_desc_n_wuser_14_wuser[9];
assign int_desc_9_wuser_15_wuser = int_desc_n_wuser_15_wuser[9];
assign int_desc_10_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[10];
assign int_desc_10_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[10];
assign int_desc_10_attr_axregion = int_desc_n_attr_axregion[10];
assign int_desc_10_attr_axqos = int_desc_n_attr_axqos[10];
assign int_desc_10_attr_axprot = int_desc_n_attr_axprot[10];
assign int_desc_10_attr_axcache = int_desc_n_attr_axcache[10];
assign int_desc_10_attr_axlock = int_desc_n_attr_axlock[10];
assign int_desc_10_attr_axburst = int_desc_n_attr_axburst[10];
assign int_desc_10_axid_0_axid = int_desc_n_axid_0_axid[10];
assign int_desc_10_axid_1_axid = int_desc_n_axid_1_axid[10];
assign int_desc_10_axid_2_axid = int_desc_n_axid_2_axid[10];
assign int_desc_10_axid_3_axid = int_desc_n_axid_3_axid[10];
assign int_desc_10_axuser_0_axuser = int_desc_n_axuser_0_axuser[10];
assign int_desc_10_axuser_1_axuser = int_desc_n_axuser_1_axuser[10];
assign int_desc_10_axuser_2_axuser = int_desc_n_axuser_2_axuser[10];
assign int_desc_10_axuser_3_axuser = int_desc_n_axuser_3_axuser[10];
assign int_desc_10_axuser_4_axuser = int_desc_n_axuser_4_axuser[10];
assign int_desc_10_axuser_5_axuser = int_desc_n_axuser_5_axuser[10];
assign int_desc_10_axuser_6_axuser = int_desc_n_axuser_6_axuser[10];
assign int_desc_10_axuser_7_axuser = int_desc_n_axuser_7_axuser[10];
assign int_desc_10_axuser_8_axuser = int_desc_n_axuser_8_axuser[10];
assign int_desc_10_axuser_9_axuser = int_desc_n_axuser_9_axuser[10];
assign int_desc_10_axuser_10_axuser = int_desc_n_axuser_10_axuser[10];
assign int_desc_10_axuser_11_axuser = int_desc_n_axuser_11_axuser[10];
assign int_desc_10_axuser_12_axuser = int_desc_n_axuser_12_axuser[10];
assign int_desc_10_axuser_13_axuser = int_desc_n_axuser_13_axuser[10];
assign int_desc_10_axuser_14_axuser = int_desc_n_axuser_14_axuser[10];
assign int_desc_10_axuser_15_axuser = int_desc_n_axuser_15_axuser[10];
assign int_desc_10_size_txn_size = int_desc_n_size_txn_size[10];
assign int_desc_10_axsize_axsize = int_desc_n_axsize_axsize[10];
assign int_desc_10_axaddr_0_addr = int_desc_n_axaddr_0_addr[10];
assign int_desc_10_axaddr_1_addr = int_desc_n_axaddr_1_addr[10];
assign int_desc_10_axaddr_2_addr = int_desc_n_axaddr_2_addr[10];
assign int_desc_10_axaddr_3_addr = int_desc_n_axaddr_3_addr[10];
assign int_desc_10_data_offset_addr = int_desc_n_data_offset_addr[10];
assign int_desc_10_wuser_0_wuser = int_desc_n_wuser_0_wuser[10];
assign int_desc_10_wuser_1_wuser = int_desc_n_wuser_1_wuser[10];
assign int_desc_10_wuser_2_wuser = int_desc_n_wuser_2_wuser[10];
assign int_desc_10_wuser_3_wuser = int_desc_n_wuser_3_wuser[10];
assign int_desc_10_wuser_4_wuser = int_desc_n_wuser_4_wuser[10];
assign int_desc_10_wuser_5_wuser = int_desc_n_wuser_5_wuser[10];
assign int_desc_10_wuser_6_wuser = int_desc_n_wuser_6_wuser[10];
assign int_desc_10_wuser_7_wuser = int_desc_n_wuser_7_wuser[10];
assign int_desc_10_wuser_8_wuser = int_desc_n_wuser_8_wuser[10];
assign int_desc_10_wuser_9_wuser = int_desc_n_wuser_9_wuser[10];
assign int_desc_10_wuser_10_wuser = int_desc_n_wuser_10_wuser[10];
assign int_desc_10_wuser_11_wuser = int_desc_n_wuser_11_wuser[10];
assign int_desc_10_wuser_12_wuser = int_desc_n_wuser_12_wuser[10];
assign int_desc_10_wuser_13_wuser = int_desc_n_wuser_13_wuser[10];
assign int_desc_10_wuser_14_wuser = int_desc_n_wuser_14_wuser[10];
assign int_desc_10_wuser_15_wuser = int_desc_n_wuser_15_wuser[10];
assign int_desc_11_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[11];
assign int_desc_11_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[11];
assign int_desc_11_attr_axregion = int_desc_n_attr_axregion[11];
assign int_desc_11_attr_axqos = int_desc_n_attr_axqos[11];
assign int_desc_11_attr_axprot = int_desc_n_attr_axprot[11];
assign int_desc_11_attr_axcache = int_desc_n_attr_axcache[11];
assign int_desc_11_attr_axlock = int_desc_n_attr_axlock[11];
assign int_desc_11_attr_axburst = int_desc_n_attr_axburst[11];
assign int_desc_11_axid_0_axid = int_desc_n_axid_0_axid[11];
assign int_desc_11_axid_1_axid = int_desc_n_axid_1_axid[11];
assign int_desc_11_axid_2_axid = int_desc_n_axid_2_axid[11];
assign int_desc_11_axid_3_axid = int_desc_n_axid_3_axid[11];
assign int_desc_11_axuser_0_axuser = int_desc_n_axuser_0_axuser[11];
assign int_desc_11_axuser_1_axuser = int_desc_n_axuser_1_axuser[11];
assign int_desc_11_axuser_2_axuser = int_desc_n_axuser_2_axuser[11];
assign int_desc_11_axuser_3_axuser = int_desc_n_axuser_3_axuser[11];
assign int_desc_11_axuser_4_axuser = int_desc_n_axuser_4_axuser[11];
assign int_desc_11_axuser_5_axuser = int_desc_n_axuser_5_axuser[11];
assign int_desc_11_axuser_6_axuser = int_desc_n_axuser_6_axuser[11];
assign int_desc_11_axuser_7_axuser = int_desc_n_axuser_7_axuser[11];
assign int_desc_11_axuser_8_axuser = int_desc_n_axuser_8_axuser[11];
assign int_desc_11_axuser_9_axuser = int_desc_n_axuser_9_axuser[11];
assign int_desc_11_axuser_10_axuser = int_desc_n_axuser_10_axuser[11];
assign int_desc_11_axuser_11_axuser = int_desc_n_axuser_11_axuser[11];
assign int_desc_11_axuser_12_axuser = int_desc_n_axuser_12_axuser[11];
assign int_desc_11_axuser_13_axuser = int_desc_n_axuser_13_axuser[11];
assign int_desc_11_axuser_14_axuser = int_desc_n_axuser_14_axuser[11];
assign int_desc_11_axuser_15_axuser = int_desc_n_axuser_15_axuser[11];
assign int_desc_11_size_txn_size = int_desc_n_size_txn_size[11];
assign int_desc_11_axsize_axsize = int_desc_n_axsize_axsize[11];
assign int_desc_11_axaddr_0_addr = int_desc_n_axaddr_0_addr[11];
assign int_desc_11_axaddr_1_addr = int_desc_n_axaddr_1_addr[11];
assign int_desc_11_axaddr_2_addr = int_desc_n_axaddr_2_addr[11];
assign int_desc_11_axaddr_3_addr = int_desc_n_axaddr_3_addr[11];
assign int_desc_11_data_offset_addr = int_desc_n_data_offset_addr[11];
assign int_desc_11_wuser_0_wuser = int_desc_n_wuser_0_wuser[11];
assign int_desc_11_wuser_1_wuser = int_desc_n_wuser_1_wuser[11];
assign int_desc_11_wuser_2_wuser = int_desc_n_wuser_2_wuser[11];
assign int_desc_11_wuser_3_wuser = int_desc_n_wuser_3_wuser[11];
assign int_desc_11_wuser_4_wuser = int_desc_n_wuser_4_wuser[11];
assign int_desc_11_wuser_5_wuser = int_desc_n_wuser_5_wuser[11];
assign int_desc_11_wuser_6_wuser = int_desc_n_wuser_6_wuser[11];
assign int_desc_11_wuser_7_wuser = int_desc_n_wuser_7_wuser[11];
assign int_desc_11_wuser_8_wuser = int_desc_n_wuser_8_wuser[11];
assign int_desc_11_wuser_9_wuser = int_desc_n_wuser_9_wuser[11];
assign int_desc_11_wuser_10_wuser = int_desc_n_wuser_10_wuser[11];
assign int_desc_11_wuser_11_wuser = int_desc_n_wuser_11_wuser[11];
assign int_desc_11_wuser_12_wuser = int_desc_n_wuser_12_wuser[11];
assign int_desc_11_wuser_13_wuser = int_desc_n_wuser_13_wuser[11];
assign int_desc_11_wuser_14_wuser = int_desc_n_wuser_14_wuser[11];
assign int_desc_11_wuser_15_wuser = int_desc_n_wuser_15_wuser[11];
assign int_desc_12_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[12];
assign int_desc_12_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[12];
assign int_desc_12_attr_axregion = int_desc_n_attr_axregion[12];
assign int_desc_12_attr_axqos = int_desc_n_attr_axqos[12];
assign int_desc_12_attr_axprot = int_desc_n_attr_axprot[12];
assign int_desc_12_attr_axcache = int_desc_n_attr_axcache[12];
assign int_desc_12_attr_axlock = int_desc_n_attr_axlock[12];
assign int_desc_12_attr_axburst = int_desc_n_attr_axburst[12];
assign int_desc_12_axid_0_axid = int_desc_n_axid_0_axid[12];
assign int_desc_12_axid_1_axid = int_desc_n_axid_1_axid[12];
assign int_desc_12_axid_2_axid = int_desc_n_axid_2_axid[12];
assign int_desc_12_axid_3_axid = int_desc_n_axid_3_axid[12];
assign int_desc_12_axuser_0_axuser = int_desc_n_axuser_0_axuser[12];
assign int_desc_12_axuser_1_axuser = int_desc_n_axuser_1_axuser[12];
assign int_desc_12_axuser_2_axuser = int_desc_n_axuser_2_axuser[12];
assign int_desc_12_axuser_3_axuser = int_desc_n_axuser_3_axuser[12];
assign int_desc_12_axuser_4_axuser = int_desc_n_axuser_4_axuser[12];
assign int_desc_12_axuser_5_axuser = int_desc_n_axuser_5_axuser[12];
assign int_desc_12_axuser_6_axuser = int_desc_n_axuser_6_axuser[12];
assign int_desc_12_axuser_7_axuser = int_desc_n_axuser_7_axuser[12];
assign int_desc_12_axuser_8_axuser = int_desc_n_axuser_8_axuser[12];
assign int_desc_12_axuser_9_axuser = int_desc_n_axuser_9_axuser[12];
assign int_desc_12_axuser_10_axuser = int_desc_n_axuser_10_axuser[12];
assign int_desc_12_axuser_11_axuser = int_desc_n_axuser_11_axuser[12];
assign int_desc_12_axuser_12_axuser = int_desc_n_axuser_12_axuser[12];
assign int_desc_12_axuser_13_axuser = int_desc_n_axuser_13_axuser[12];
assign int_desc_12_axuser_14_axuser = int_desc_n_axuser_14_axuser[12];
assign int_desc_12_axuser_15_axuser = int_desc_n_axuser_15_axuser[12];
assign int_desc_12_size_txn_size = int_desc_n_size_txn_size[12];
assign int_desc_12_axsize_axsize = int_desc_n_axsize_axsize[12];
assign int_desc_12_axaddr_0_addr = int_desc_n_axaddr_0_addr[12];
assign int_desc_12_axaddr_1_addr = int_desc_n_axaddr_1_addr[12];
assign int_desc_12_axaddr_2_addr = int_desc_n_axaddr_2_addr[12];
assign int_desc_12_axaddr_3_addr = int_desc_n_axaddr_3_addr[12];
assign int_desc_12_data_offset_addr = int_desc_n_data_offset_addr[12];
assign int_desc_12_wuser_0_wuser = int_desc_n_wuser_0_wuser[12];
assign int_desc_12_wuser_1_wuser = int_desc_n_wuser_1_wuser[12];
assign int_desc_12_wuser_2_wuser = int_desc_n_wuser_2_wuser[12];
assign int_desc_12_wuser_3_wuser = int_desc_n_wuser_3_wuser[12];
assign int_desc_12_wuser_4_wuser = int_desc_n_wuser_4_wuser[12];
assign int_desc_12_wuser_5_wuser = int_desc_n_wuser_5_wuser[12];
assign int_desc_12_wuser_6_wuser = int_desc_n_wuser_6_wuser[12];
assign int_desc_12_wuser_7_wuser = int_desc_n_wuser_7_wuser[12];
assign int_desc_12_wuser_8_wuser = int_desc_n_wuser_8_wuser[12];
assign int_desc_12_wuser_9_wuser = int_desc_n_wuser_9_wuser[12];
assign int_desc_12_wuser_10_wuser = int_desc_n_wuser_10_wuser[12];
assign int_desc_12_wuser_11_wuser = int_desc_n_wuser_11_wuser[12];
assign int_desc_12_wuser_12_wuser = int_desc_n_wuser_12_wuser[12];
assign int_desc_12_wuser_13_wuser = int_desc_n_wuser_13_wuser[12];
assign int_desc_12_wuser_14_wuser = int_desc_n_wuser_14_wuser[12];
assign int_desc_12_wuser_15_wuser = int_desc_n_wuser_15_wuser[12];
assign int_desc_13_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[13];
assign int_desc_13_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[13];
assign int_desc_13_attr_axregion = int_desc_n_attr_axregion[13];
assign int_desc_13_attr_axqos = int_desc_n_attr_axqos[13];
assign int_desc_13_attr_axprot = int_desc_n_attr_axprot[13];
assign int_desc_13_attr_axcache = int_desc_n_attr_axcache[13];
assign int_desc_13_attr_axlock = int_desc_n_attr_axlock[13];
assign int_desc_13_attr_axburst = int_desc_n_attr_axburst[13];
assign int_desc_13_axid_0_axid = int_desc_n_axid_0_axid[13];
assign int_desc_13_axid_1_axid = int_desc_n_axid_1_axid[13];
assign int_desc_13_axid_2_axid = int_desc_n_axid_2_axid[13];
assign int_desc_13_axid_3_axid = int_desc_n_axid_3_axid[13];
assign int_desc_13_axuser_0_axuser = int_desc_n_axuser_0_axuser[13];
assign int_desc_13_axuser_1_axuser = int_desc_n_axuser_1_axuser[13];
assign int_desc_13_axuser_2_axuser = int_desc_n_axuser_2_axuser[13];
assign int_desc_13_axuser_3_axuser = int_desc_n_axuser_3_axuser[13];
assign int_desc_13_axuser_4_axuser = int_desc_n_axuser_4_axuser[13];
assign int_desc_13_axuser_5_axuser = int_desc_n_axuser_5_axuser[13];
assign int_desc_13_axuser_6_axuser = int_desc_n_axuser_6_axuser[13];
assign int_desc_13_axuser_7_axuser = int_desc_n_axuser_7_axuser[13];
assign int_desc_13_axuser_8_axuser = int_desc_n_axuser_8_axuser[13];
assign int_desc_13_axuser_9_axuser = int_desc_n_axuser_9_axuser[13];
assign int_desc_13_axuser_10_axuser = int_desc_n_axuser_10_axuser[13];
assign int_desc_13_axuser_11_axuser = int_desc_n_axuser_11_axuser[13];
assign int_desc_13_axuser_12_axuser = int_desc_n_axuser_12_axuser[13];
assign int_desc_13_axuser_13_axuser = int_desc_n_axuser_13_axuser[13];
assign int_desc_13_axuser_14_axuser = int_desc_n_axuser_14_axuser[13];
assign int_desc_13_axuser_15_axuser = int_desc_n_axuser_15_axuser[13];
assign int_desc_13_size_txn_size = int_desc_n_size_txn_size[13];
assign int_desc_13_axsize_axsize = int_desc_n_axsize_axsize[13];
assign int_desc_13_axaddr_0_addr = int_desc_n_axaddr_0_addr[13];
assign int_desc_13_axaddr_1_addr = int_desc_n_axaddr_1_addr[13];
assign int_desc_13_axaddr_2_addr = int_desc_n_axaddr_2_addr[13];
assign int_desc_13_axaddr_3_addr = int_desc_n_axaddr_3_addr[13];
assign int_desc_13_data_offset_addr = int_desc_n_data_offset_addr[13];
assign int_desc_13_wuser_0_wuser = int_desc_n_wuser_0_wuser[13];
assign int_desc_13_wuser_1_wuser = int_desc_n_wuser_1_wuser[13];
assign int_desc_13_wuser_2_wuser = int_desc_n_wuser_2_wuser[13];
assign int_desc_13_wuser_3_wuser = int_desc_n_wuser_3_wuser[13];
assign int_desc_13_wuser_4_wuser = int_desc_n_wuser_4_wuser[13];
assign int_desc_13_wuser_5_wuser = int_desc_n_wuser_5_wuser[13];
assign int_desc_13_wuser_6_wuser = int_desc_n_wuser_6_wuser[13];
assign int_desc_13_wuser_7_wuser = int_desc_n_wuser_7_wuser[13];
assign int_desc_13_wuser_8_wuser = int_desc_n_wuser_8_wuser[13];
assign int_desc_13_wuser_9_wuser = int_desc_n_wuser_9_wuser[13];
assign int_desc_13_wuser_10_wuser = int_desc_n_wuser_10_wuser[13];
assign int_desc_13_wuser_11_wuser = int_desc_n_wuser_11_wuser[13];
assign int_desc_13_wuser_12_wuser = int_desc_n_wuser_12_wuser[13];
assign int_desc_13_wuser_13_wuser = int_desc_n_wuser_13_wuser[13];
assign int_desc_13_wuser_14_wuser = int_desc_n_wuser_14_wuser[13];
assign int_desc_13_wuser_15_wuser = int_desc_n_wuser_15_wuser[13];
assign int_desc_14_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[14];
assign int_desc_14_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[14];
assign int_desc_14_attr_axregion = int_desc_n_attr_axregion[14];
assign int_desc_14_attr_axqos = int_desc_n_attr_axqos[14];
assign int_desc_14_attr_axprot = int_desc_n_attr_axprot[14];
assign int_desc_14_attr_axcache = int_desc_n_attr_axcache[14];
assign int_desc_14_attr_axlock = int_desc_n_attr_axlock[14];
assign int_desc_14_attr_axburst = int_desc_n_attr_axburst[14];
assign int_desc_14_axid_0_axid = int_desc_n_axid_0_axid[14];
assign int_desc_14_axid_1_axid = int_desc_n_axid_1_axid[14];
assign int_desc_14_axid_2_axid = int_desc_n_axid_2_axid[14];
assign int_desc_14_axid_3_axid = int_desc_n_axid_3_axid[14];
assign int_desc_14_axuser_0_axuser = int_desc_n_axuser_0_axuser[14];
assign int_desc_14_axuser_1_axuser = int_desc_n_axuser_1_axuser[14];
assign int_desc_14_axuser_2_axuser = int_desc_n_axuser_2_axuser[14];
assign int_desc_14_axuser_3_axuser = int_desc_n_axuser_3_axuser[14];
assign int_desc_14_axuser_4_axuser = int_desc_n_axuser_4_axuser[14];
assign int_desc_14_axuser_5_axuser = int_desc_n_axuser_5_axuser[14];
assign int_desc_14_axuser_6_axuser = int_desc_n_axuser_6_axuser[14];
assign int_desc_14_axuser_7_axuser = int_desc_n_axuser_7_axuser[14];
assign int_desc_14_axuser_8_axuser = int_desc_n_axuser_8_axuser[14];
assign int_desc_14_axuser_9_axuser = int_desc_n_axuser_9_axuser[14];
assign int_desc_14_axuser_10_axuser = int_desc_n_axuser_10_axuser[14];
assign int_desc_14_axuser_11_axuser = int_desc_n_axuser_11_axuser[14];
assign int_desc_14_axuser_12_axuser = int_desc_n_axuser_12_axuser[14];
assign int_desc_14_axuser_13_axuser = int_desc_n_axuser_13_axuser[14];
assign int_desc_14_axuser_14_axuser = int_desc_n_axuser_14_axuser[14];
assign int_desc_14_axuser_15_axuser = int_desc_n_axuser_15_axuser[14];
assign int_desc_14_size_txn_size = int_desc_n_size_txn_size[14];
assign int_desc_14_axsize_axsize = int_desc_n_axsize_axsize[14];
assign int_desc_14_axaddr_0_addr = int_desc_n_axaddr_0_addr[14];
assign int_desc_14_axaddr_1_addr = int_desc_n_axaddr_1_addr[14];
assign int_desc_14_axaddr_2_addr = int_desc_n_axaddr_2_addr[14];
assign int_desc_14_axaddr_3_addr = int_desc_n_axaddr_3_addr[14];
assign int_desc_14_data_offset_addr = int_desc_n_data_offset_addr[14];
assign int_desc_14_wuser_0_wuser = int_desc_n_wuser_0_wuser[14];
assign int_desc_14_wuser_1_wuser = int_desc_n_wuser_1_wuser[14];
assign int_desc_14_wuser_2_wuser = int_desc_n_wuser_2_wuser[14];
assign int_desc_14_wuser_3_wuser = int_desc_n_wuser_3_wuser[14];
assign int_desc_14_wuser_4_wuser = int_desc_n_wuser_4_wuser[14];
assign int_desc_14_wuser_5_wuser = int_desc_n_wuser_5_wuser[14];
assign int_desc_14_wuser_6_wuser = int_desc_n_wuser_6_wuser[14];
assign int_desc_14_wuser_7_wuser = int_desc_n_wuser_7_wuser[14];
assign int_desc_14_wuser_8_wuser = int_desc_n_wuser_8_wuser[14];
assign int_desc_14_wuser_9_wuser = int_desc_n_wuser_9_wuser[14];
assign int_desc_14_wuser_10_wuser = int_desc_n_wuser_10_wuser[14];
assign int_desc_14_wuser_11_wuser = int_desc_n_wuser_11_wuser[14];
assign int_desc_14_wuser_12_wuser = int_desc_n_wuser_12_wuser[14];
assign int_desc_14_wuser_13_wuser = int_desc_n_wuser_13_wuser[14];
assign int_desc_14_wuser_14_wuser = int_desc_n_wuser_14_wuser[14];
assign int_desc_14_wuser_15_wuser = int_desc_n_wuser_15_wuser[14];
assign int_desc_15_txn_type_wr_strb = int_desc_n_txn_type_wr_strb[15];
assign int_desc_15_txn_type_wr_rd = int_desc_n_txn_type_wr_rd[15];
assign int_desc_15_attr_axregion = int_desc_n_attr_axregion[15];
assign int_desc_15_attr_axqos = int_desc_n_attr_axqos[15];
assign int_desc_15_attr_axprot = int_desc_n_attr_axprot[15];
assign int_desc_15_attr_axcache = int_desc_n_attr_axcache[15];
assign int_desc_15_attr_axlock = int_desc_n_attr_axlock[15];
assign int_desc_15_attr_axburst = int_desc_n_attr_axburst[15];
assign int_desc_15_axid_0_axid = int_desc_n_axid_0_axid[15];
assign int_desc_15_axid_1_axid = int_desc_n_axid_1_axid[15];
assign int_desc_15_axid_2_axid = int_desc_n_axid_2_axid[15];
assign int_desc_15_axid_3_axid = int_desc_n_axid_3_axid[15];
assign int_desc_15_axuser_0_axuser = int_desc_n_axuser_0_axuser[15];
assign int_desc_15_axuser_1_axuser = int_desc_n_axuser_1_axuser[15];
assign int_desc_15_axuser_2_axuser = int_desc_n_axuser_2_axuser[15];
assign int_desc_15_axuser_3_axuser = int_desc_n_axuser_3_axuser[15];
assign int_desc_15_axuser_4_axuser = int_desc_n_axuser_4_axuser[15];
assign int_desc_15_axuser_5_axuser = int_desc_n_axuser_5_axuser[15];
assign int_desc_15_axuser_6_axuser = int_desc_n_axuser_6_axuser[15];
assign int_desc_15_axuser_7_axuser = int_desc_n_axuser_7_axuser[15];
assign int_desc_15_axuser_8_axuser = int_desc_n_axuser_8_axuser[15];
assign int_desc_15_axuser_9_axuser = int_desc_n_axuser_9_axuser[15];
assign int_desc_15_axuser_10_axuser = int_desc_n_axuser_10_axuser[15];
assign int_desc_15_axuser_11_axuser = int_desc_n_axuser_11_axuser[15];
assign int_desc_15_axuser_12_axuser = int_desc_n_axuser_12_axuser[15];
assign int_desc_15_axuser_13_axuser = int_desc_n_axuser_13_axuser[15];
assign int_desc_15_axuser_14_axuser = int_desc_n_axuser_14_axuser[15];
assign int_desc_15_axuser_15_axuser = int_desc_n_axuser_15_axuser[15];
assign int_desc_15_size_txn_size = int_desc_n_size_txn_size[15];
assign int_desc_15_axsize_axsize = int_desc_n_axsize_axsize[15];
assign int_desc_15_axaddr_0_addr = int_desc_n_axaddr_0_addr[15];
assign int_desc_15_axaddr_1_addr = int_desc_n_axaddr_1_addr[15];
assign int_desc_15_axaddr_2_addr = int_desc_n_axaddr_2_addr[15];
assign int_desc_15_axaddr_3_addr = int_desc_n_axaddr_3_addr[15];
assign int_desc_15_data_offset_addr = int_desc_n_data_offset_addr[15];
assign int_desc_15_wuser_0_wuser = int_desc_n_wuser_0_wuser[15];
assign int_desc_15_wuser_1_wuser = int_desc_n_wuser_1_wuser[15];
assign int_desc_15_wuser_2_wuser = int_desc_n_wuser_2_wuser[15];
assign int_desc_15_wuser_3_wuser = int_desc_n_wuser_3_wuser[15];
assign int_desc_15_wuser_4_wuser = int_desc_n_wuser_4_wuser[15];
assign int_desc_15_wuser_5_wuser = int_desc_n_wuser_5_wuser[15];
assign int_desc_15_wuser_6_wuser = int_desc_n_wuser_6_wuser[15];
assign int_desc_15_wuser_7_wuser = int_desc_n_wuser_7_wuser[15];
assign int_desc_15_wuser_8_wuser = int_desc_n_wuser_8_wuser[15];
assign int_desc_15_wuser_9_wuser = int_desc_n_wuser_9_wuser[15];
assign int_desc_15_wuser_10_wuser = int_desc_n_wuser_10_wuser[15];
assign int_desc_15_wuser_11_wuser = int_desc_n_wuser_11_wuser[15];
assign int_desc_15_wuser_12_wuser = int_desc_n_wuser_12_wuser[15];
assign int_desc_15_wuser_13_wuser = int_desc_n_wuser_13_wuser[15];
assign int_desc_15_wuser_14_wuser = int_desc_n_wuser_14_wuser[15];
assign int_desc_15_wuser_15_wuser = int_desc_n_wuser_15_wuser[15];


assign	int_desc_n_data_host_addr_0_addr[0] = int_desc_0_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[0] = int_desc_0_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[0] = int_desc_0_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[0] = int_desc_0_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[0] = int_desc_0_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[0] = int_desc_0_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[0] = int_desc_0_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[0] = int_desc_0_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[1] = int_desc_1_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[1] = int_desc_1_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[1] = int_desc_1_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[1] = int_desc_1_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[1] = int_desc_1_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[1] = int_desc_1_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[1] = int_desc_1_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[1] = int_desc_1_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[2] = int_desc_2_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[2] = int_desc_2_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[2] = int_desc_2_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[2] = int_desc_2_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[2] = int_desc_2_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[2] = int_desc_2_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[2] = int_desc_2_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[2] = int_desc_2_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[3] = int_desc_3_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[3] = int_desc_3_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[3] = int_desc_3_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[3] = int_desc_3_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[3] = int_desc_3_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[3] = int_desc_3_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[3] = int_desc_3_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[3] = int_desc_3_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[4] = int_desc_4_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[4] = int_desc_4_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[4] = int_desc_4_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[4] = int_desc_4_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[4] = int_desc_4_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[4] = int_desc_4_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[4] = int_desc_4_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[4] = int_desc_4_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[5] = int_desc_5_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[5] = int_desc_5_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[5] = int_desc_5_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[5] = int_desc_5_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[5] = int_desc_5_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[5] = int_desc_5_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[5] = int_desc_5_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[5] = int_desc_5_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[6] = int_desc_6_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[6] = int_desc_6_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[6] = int_desc_6_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[6] = int_desc_6_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[6] = int_desc_6_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[6] = int_desc_6_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[6] = int_desc_6_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[6] = int_desc_6_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[7] = int_desc_7_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[7] = int_desc_7_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[7] = int_desc_7_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[7] = int_desc_7_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[7] = int_desc_7_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[7] = int_desc_7_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[7] = int_desc_7_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[7] = int_desc_7_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[8] = int_desc_8_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[8] = int_desc_8_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[8] = int_desc_8_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[8] = int_desc_8_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[8] = int_desc_8_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[8] = int_desc_8_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[8] = int_desc_8_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[8] = int_desc_8_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[9] = int_desc_9_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[9] = int_desc_9_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[9] = int_desc_9_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[9] = int_desc_9_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[9] = int_desc_9_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[9] = int_desc_9_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[9] = int_desc_9_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[9] = int_desc_9_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[10] = int_desc_10_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[10] = int_desc_10_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[10] = int_desc_10_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[10] = int_desc_10_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[10] = int_desc_10_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[10] = int_desc_10_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[10] = int_desc_10_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[10] = int_desc_10_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[11] = int_desc_11_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[11] = int_desc_11_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[11] = int_desc_11_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[11] = int_desc_11_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[11] = int_desc_11_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[11] = int_desc_11_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[11] = int_desc_11_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[11] = int_desc_11_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[12] = int_desc_12_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[12] = int_desc_12_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[12] = int_desc_12_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[12] = int_desc_12_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[12] = int_desc_12_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[12] = int_desc_12_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[12] = int_desc_12_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[12] = int_desc_12_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[13] = int_desc_13_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[13] = int_desc_13_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[13] = int_desc_13_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[13] = int_desc_13_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[13] = int_desc_13_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[13] = int_desc_13_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[13] = int_desc_13_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[13] = int_desc_13_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[14] = int_desc_14_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[14] = int_desc_14_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[14] = int_desc_14_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[14] = int_desc_14_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[14] = int_desc_14_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[14] = int_desc_14_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[14] = int_desc_14_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[14] = int_desc_14_wstrb_host_addr_3_addr;
assign	int_desc_n_data_host_addr_0_addr[15] = int_desc_15_data_host_addr_0_addr;
assign	int_desc_n_data_host_addr_1_addr[15] = int_desc_15_data_host_addr_1_addr;
assign	int_desc_n_data_host_addr_2_addr[15] = int_desc_15_data_host_addr_2_addr;
assign	int_desc_n_data_host_addr_3_addr[15] = int_desc_15_data_host_addr_3_addr;
assign	int_desc_n_wstrb_host_addr_0_addr[15] = int_desc_15_wstrb_host_addr_0_addr;
assign	int_desc_n_wstrb_host_addr_1_addr[15] = int_desc_15_wstrb_host_addr_1_addr;
assign	int_desc_n_wstrb_host_addr_2_addr[15] = int_desc_15_wstrb_host_addr_2_addr;
assign	int_desc_n_wstrb_host_addr_3_addr[15] = int_desc_15_wstrb_host_addr_3_addr;
assign	int_desc_n_xuser_0_xuser[0] = int_desc_0_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[0] = int_desc_0_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[0] = int_desc_0_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[0] = int_desc_0_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[0] = int_desc_0_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[0] = int_desc_0_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[0] = int_desc_0_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[0] = int_desc_0_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[0] = int_desc_0_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[0] = int_desc_0_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[0] = int_desc_0_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[0] = int_desc_0_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[0] = int_desc_0_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[0] = int_desc_0_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[0] = int_desc_0_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[0] = int_desc_0_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[1] = int_desc_1_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[1] = int_desc_1_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[1] = int_desc_1_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[1] = int_desc_1_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[1] = int_desc_1_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[1] = int_desc_1_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[1] = int_desc_1_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[1] = int_desc_1_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[1] = int_desc_1_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[1] = int_desc_1_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[1] = int_desc_1_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[1] = int_desc_1_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[1] = int_desc_1_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[1] = int_desc_1_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[1] = int_desc_1_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[1] = int_desc_1_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[2] = int_desc_2_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[2] = int_desc_2_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[2] = int_desc_2_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[2] = int_desc_2_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[2] = int_desc_2_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[2] = int_desc_2_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[2] = int_desc_2_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[2] = int_desc_2_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[2] = int_desc_2_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[2] = int_desc_2_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[2] = int_desc_2_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[2] = int_desc_2_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[2] = int_desc_2_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[2] = int_desc_2_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[2] = int_desc_2_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[2] = int_desc_2_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[3] = int_desc_3_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[3] = int_desc_3_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[3] = int_desc_3_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[3] = int_desc_3_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[3] = int_desc_3_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[3] = int_desc_3_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[3] = int_desc_3_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[3] = int_desc_3_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[3] = int_desc_3_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[3] = int_desc_3_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[3] = int_desc_3_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[3] = int_desc_3_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[3] = int_desc_3_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[3] = int_desc_3_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[3] = int_desc_3_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[3] = int_desc_3_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[4] = int_desc_4_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[4] = int_desc_4_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[4] = int_desc_4_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[4] = int_desc_4_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[4] = int_desc_4_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[4] = int_desc_4_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[4] = int_desc_4_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[4] = int_desc_4_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[4] = int_desc_4_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[4] = int_desc_4_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[4] = int_desc_4_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[4] = int_desc_4_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[4] = int_desc_4_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[4] = int_desc_4_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[4] = int_desc_4_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[4] = int_desc_4_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[5] = int_desc_5_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[5] = int_desc_5_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[5] = int_desc_5_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[5] = int_desc_5_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[5] = int_desc_5_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[5] = int_desc_5_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[5] = int_desc_5_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[5] = int_desc_5_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[5] = int_desc_5_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[5] = int_desc_5_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[5] = int_desc_5_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[5] = int_desc_5_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[5] = int_desc_5_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[5] = int_desc_5_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[5] = int_desc_5_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[5] = int_desc_5_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[6] = int_desc_6_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[6] = int_desc_6_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[6] = int_desc_6_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[6] = int_desc_6_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[6] = int_desc_6_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[6] = int_desc_6_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[6] = int_desc_6_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[6] = int_desc_6_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[6] = int_desc_6_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[6] = int_desc_6_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[6] = int_desc_6_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[6] = int_desc_6_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[6] = int_desc_6_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[6] = int_desc_6_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[6] = int_desc_6_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[6] = int_desc_6_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[7] = int_desc_7_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[7] = int_desc_7_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[7] = int_desc_7_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[7] = int_desc_7_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[7] = int_desc_7_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[7] = int_desc_7_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[7] = int_desc_7_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[7] = int_desc_7_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[7] = int_desc_7_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[7] = int_desc_7_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[7] = int_desc_7_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[7] = int_desc_7_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[7] = int_desc_7_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[7] = int_desc_7_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[7] = int_desc_7_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[7] = int_desc_7_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[8] = int_desc_8_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[8] = int_desc_8_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[8] = int_desc_8_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[8] = int_desc_8_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[8] = int_desc_8_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[8] = int_desc_8_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[8] = int_desc_8_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[8] = int_desc_8_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[8] = int_desc_8_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[8] = int_desc_8_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[8] = int_desc_8_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[8] = int_desc_8_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[8] = int_desc_8_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[8] = int_desc_8_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[8] = int_desc_8_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[8] = int_desc_8_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[9] = int_desc_9_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[9] = int_desc_9_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[9] = int_desc_9_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[9] = int_desc_9_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[9] = int_desc_9_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[9] = int_desc_9_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[9] = int_desc_9_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[9] = int_desc_9_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[9] = int_desc_9_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[9] = int_desc_9_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[9] = int_desc_9_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[9] = int_desc_9_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[9] = int_desc_9_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[9] = int_desc_9_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[9] = int_desc_9_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[9] = int_desc_9_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[10] = int_desc_10_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[10] = int_desc_10_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[10] = int_desc_10_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[10] = int_desc_10_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[10] = int_desc_10_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[10] = int_desc_10_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[10] = int_desc_10_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[10] = int_desc_10_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[10] = int_desc_10_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[10] = int_desc_10_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[10] = int_desc_10_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[10] = int_desc_10_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[10] = int_desc_10_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[10] = int_desc_10_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[10] = int_desc_10_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[10] = int_desc_10_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[11] = int_desc_11_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[11] = int_desc_11_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[11] = int_desc_11_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[11] = int_desc_11_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[11] = int_desc_11_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[11] = int_desc_11_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[11] = int_desc_11_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[11] = int_desc_11_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[11] = int_desc_11_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[11] = int_desc_11_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[11] = int_desc_11_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[11] = int_desc_11_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[11] = int_desc_11_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[11] = int_desc_11_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[11] = int_desc_11_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[11] = int_desc_11_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[12] = int_desc_12_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[12] = int_desc_12_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[12] = int_desc_12_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[12] = int_desc_12_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[12] = int_desc_12_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[12] = int_desc_12_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[12] = int_desc_12_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[12] = int_desc_12_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[12] = int_desc_12_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[12] = int_desc_12_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[12] = int_desc_12_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[12] = int_desc_12_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[12] = int_desc_12_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[12] = int_desc_12_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[12] = int_desc_12_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[12] = int_desc_12_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[13] = int_desc_13_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[13] = int_desc_13_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[13] = int_desc_13_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[13] = int_desc_13_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[13] = int_desc_13_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[13] = int_desc_13_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[13] = int_desc_13_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[13] = int_desc_13_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[13] = int_desc_13_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[13] = int_desc_13_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[13] = int_desc_13_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[13] = int_desc_13_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[13] = int_desc_13_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[13] = int_desc_13_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[13] = int_desc_13_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[13] = int_desc_13_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[14] = int_desc_14_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[14] = int_desc_14_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[14] = int_desc_14_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[14] = int_desc_14_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[14] = int_desc_14_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[14] = int_desc_14_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[14] = int_desc_14_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[14] = int_desc_14_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[14] = int_desc_14_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[14] = int_desc_14_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[14] = int_desc_14_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[14] = int_desc_14_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[14] = int_desc_14_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[14] = int_desc_14_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[14] = int_desc_14_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[14] = int_desc_14_xuser_15_xuser;
assign	int_desc_n_xuser_0_xuser[15] = int_desc_15_xuser_0_xuser;
assign	int_desc_n_xuser_1_xuser[15] = int_desc_15_xuser_1_xuser;
assign	int_desc_n_xuser_2_xuser[15] = int_desc_15_xuser_2_xuser;
assign	int_desc_n_xuser_3_xuser[15] = int_desc_15_xuser_3_xuser;
assign	int_desc_n_xuser_4_xuser[15] = int_desc_15_xuser_4_xuser;
assign	int_desc_n_xuser_5_xuser[15] = int_desc_15_xuser_5_xuser;
assign	int_desc_n_xuser_6_xuser[15] = int_desc_15_xuser_6_xuser;
assign	int_desc_n_xuser_7_xuser[15] = int_desc_15_xuser_7_xuser;
assign	int_desc_n_xuser_8_xuser[15] = int_desc_15_xuser_8_xuser;
assign	int_desc_n_xuser_9_xuser[15] = int_desc_15_xuser_9_xuser;
assign	int_desc_n_xuser_10_xuser[15] = int_desc_15_xuser_10_xuser;
assign	int_desc_n_xuser_11_xuser[15] = int_desc_15_xuser_11_xuser;
assign	int_desc_n_xuser_12_xuser[15] = int_desc_15_xuser_12_xuser;
assign	int_desc_n_xuser_13_xuser[15] = int_desc_15_xuser_13_xuser;
assign	int_desc_n_xuser_14_xuser[15] = int_desc_15_xuser_14_xuser;
assign	int_desc_n_xuser_15_xuser[15] = int_desc_15_xuser_15_xuser;
