/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */

 // Inputs
		 ,.int_desc_0_data_host_addr_0_addr(int_desc_0_data_host_addr_0_addr[31:0])
		 ,.int_desc_0_data_host_addr_1_addr(int_desc_0_data_host_addr_1_addr[31:0])
		 ,.int_desc_0_data_host_addr_2_addr(int_desc_0_data_host_addr_2_addr[31:0])
		 ,.int_desc_0_data_host_addr_3_addr(int_desc_0_data_host_addr_3_addr[31:0])
		 ,.int_desc_0_wstrb_host_addr_0_addr(int_desc_0_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_0_wstrb_host_addr_1_addr(int_desc_0_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_0_wstrb_host_addr_2_addr(int_desc_0_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_0_wstrb_host_addr_3_addr(int_desc_0_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_1_data_host_addr_0_addr(int_desc_1_data_host_addr_0_addr[31:0])
		 ,.int_desc_1_data_host_addr_1_addr(int_desc_1_data_host_addr_1_addr[31:0])
		 ,.int_desc_1_data_host_addr_2_addr(int_desc_1_data_host_addr_2_addr[31:0])
		 ,.int_desc_1_data_host_addr_3_addr(int_desc_1_data_host_addr_3_addr[31:0])
		 ,.int_desc_1_wstrb_host_addr_0_addr(int_desc_1_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_1_wstrb_host_addr_1_addr(int_desc_1_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_1_wstrb_host_addr_2_addr(int_desc_1_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_1_wstrb_host_addr_3_addr(int_desc_1_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_2_data_host_addr_0_addr(int_desc_2_data_host_addr_0_addr[31:0])
		 ,.int_desc_2_data_host_addr_1_addr(int_desc_2_data_host_addr_1_addr[31:0])
		 ,.int_desc_2_data_host_addr_2_addr(int_desc_2_data_host_addr_2_addr[31:0])
		 ,.int_desc_2_data_host_addr_3_addr(int_desc_2_data_host_addr_3_addr[31:0])
		 ,.int_desc_2_wstrb_host_addr_0_addr(int_desc_2_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_2_wstrb_host_addr_1_addr(int_desc_2_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_2_wstrb_host_addr_2_addr(int_desc_2_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_2_wstrb_host_addr_3_addr(int_desc_2_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_3_data_host_addr_0_addr(int_desc_3_data_host_addr_0_addr[31:0])
		 ,.int_desc_3_data_host_addr_1_addr(int_desc_3_data_host_addr_1_addr[31:0])
		 ,.int_desc_3_data_host_addr_2_addr(int_desc_3_data_host_addr_2_addr[31:0])
		 ,.int_desc_3_data_host_addr_3_addr(int_desc_3_data_host_addr_3_addr[31:0])
		 ,.int_desc_3_wstrb_host_addr_0_addr(int_desc_3_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_3_wstrb_host_addr_1_addr(int_desc_3_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_3_wstrb_host_addr_2_addr(int_desc_3_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_3_wstrb_host_addr_3_addr(int_desc_3_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_4_data_host_addr_0_addr(int_desc_4_data_host_addr_0_addr[31:0])
		 ,.int_desc_4_data_host_addr_1_addr(int_desc_4_data_host_addr_1_addr[31:0])
		 ,.int_desc_4_data_host_addr_2_addr(int_desc_4_data_host_addr_2_addr[31:0])
		 ,.int_desc_4_data_host_addr_3_addr(int_desc_4_data_host_addr_3_addr[31:0])
		 ,.int_desc_4_wstrb_host_addr_0_addr(int_desc_4_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_4_wstrb_host_addr_1_addr(int_desc_4_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_4_wstrb_host_addr_2_addr(int_desc_4_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_4_wstrb_host_addr_3_addr(int_desc_4_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_5_data_host_addr_0_addr(int_desc_5_data_host_addr_0_addr[31:0])
		 ,.int_desc_5_data_host_addr_1_addr(int_desc_5_data_host_addr_1_addr[31:0])
		 ,.int_desc_5_data_host_addr_2_addr(int_desc_5_data_host_addr_2_addr[31:0])
		 ,.int_desc_5_data_host_addr_3_addr(int_desc_5_data_host_addr_3_addr[31:0])
		 ,.int_desc_5_wstrb_host_addr_0_addr(int_desc_5_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_5_wstrb_host_addr_1_addr(int_desc_5_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_5_wstrb_host_addr_2_addr(int_desc_5_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_5_wstrb_host_addr_3_addr(int_desc_5_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_6_data_host_addr_0_addr(int_desc_6_data_host_addr_0_addr[31:0])
		 ,.int_desc_6_data_host_addr_1_addr(int_desc_6_data_host_addr_1_addr[31:0])
		 ,.int_desc_6_data_host_addr_2_addr(int_desc_6_data_host_addr_2_addr[31:0])
		 ,.int_desc_6_data_host_addr_3_addr(int_desc_6_data_host_addr_3_addr[31:0])
		 ,.int_desc_6_wstrb_host_addr_0_addr(int_desc_6_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_6_wstrb_host_addr_1_addr(int_desc_6_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_6_wstrb_host_addr_2_addr(int_desc_6_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_6_wstrb_host_addr_3_addr(int_desc_6_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_7_data_host_addr_0_addr(int_desc_7_data_host_addr_0_addr[31:0])
		 ,.int_desc_7_data_host_addr_1_addr(int_desc_7_data_host_addr_1_addr[31:0])
		 ,.int_desc_7_data_host_addr_2_addr(int_desc_7_data_host_addr_2_addr[31:0])
		 ,.int_desc_7_data_host_addr_3_addr(int_desc_7_data_host_addr_3_addr[31:0])
		 ,.int_desc_7_wstrb_host_addr_0_addr(int_desc_7_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_7_wstrb_host_addr_1_addr(int_desc_7_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_7_wstrb_host_addr_2_addr(int_desc_7_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_7_wstrb_host_addr_3_addr(int_desc_7_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_8_data_host_addr_0_addr(int_desc_8_data_host_addr_0_addr[31:0])
		 ,.int_desc_8_data_host_addr_1_addr(int_desc_8_data_host_addr_1_addr[31:0])
		 ,.int_desc_8_data_host_addr_2_addr(int_desc_8_data_host_addr_2_addr[31:0])
		 ,.int_desc_8_data_host_addr_3_addr(int_desc_8_data_host_addr_3_addr[31:0])
		 ,.int_desc_8_wstrb_host_addr_0_addr(int_desc_8_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_8_wstrb_host_addr_1_addr(int_desc_8_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_8_wstrb_host_addr_2_addr(int_desc_8_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_8_wstrb_host_addr_3_addr(int_desc_8_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_9_data_host_addr_0_addr(int_desc_9_data_host_addr_0_addr[31:0])
		 ,.int_desc_9_data_host_addr_1_addr(int_desc_9_data_host_addr_1_addr[31:0])
		 ,.int_desc_9_data_host_addr_2_addr(int_desc_9_data_host_addr_2_addr[31:0])
		 ,.int_desc_9_data_host_addr_3_addr(int_desc_9_data_host_addr_3_addr[31:0])
		 ,.int_desc_9_wstrb_host_addr_0_addr(int_desc_9_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_9_wstrb_host_addr_1_addr(int_desc_9_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_9_wstrb_host_addr_2_addr(int_desc_9_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_9_wstrb_host_addr_3_addr(int_desc_9_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_10_data_host_addr_0_addr(int_desc_10_data_host_addr_0_addr[31:0])
		 ,.int_desc_10_data_host_addr_1_addr(int_desc_10_data_host_addr_1_addr[31:0])
		 ,.int_desc_10_data_host_addr_2_addr(int_desc_10_data_host_addr_2_addr[31:0])
		 ,.int_desc_10_data_host_addr_3_addr(int_desc_10_data_host_addr_3_addr[31:0])
		 ,.int_desc_10_wstrb_host_addr_0_addr(int_desc_10_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_10_wstrb_host_addr_1_addr(int_desc_10_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_10_wstrb_host_addr_2_addr(int_desc_10_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_10_wstrb_host_addr_3_addr(int_desc_10_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_11_data_host_addr_0_addr(int_desc_11_data_host_addr_0_addr[31:0])
		 ,.int_desc_11_data_host_addr_1_addr(int_desc_11_data_host_addr_1_addr[31:0])
		 ,.int_desc_11_data_host_addr_2_addr(int_desc_11_data_host_addr_2_addr[31:0])
		 ,.int_desc_11_data_host_addr_3_addr(int_desc_11_data_host_addr_3_addr[31:0])
		 ,.int_desc_11_wstrb_host_addr_0_addr(int_desc_11_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_11_wstrb_host_addr_1_addr(int_desc_11_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_11_wstrb_host_addr_2_addr(int_desc_11_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_11_wstrb_host_addr_3_addr(int_desc_11_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_12_data_host_addr_0_addr(int_desc_12_data_host_addr_0_addr[31:0])
		 ,.int_desc_12_data_host_addr_1_addr(int_desc_12_data_host_addr_1_addr[31:0])
		 ,.int_desc_12_data_host_addr_2_addr(int_desc_12_data_host_addr_2_addr[31:0])
		 ,.int_desc_12_data_host_addr_3_addr(int_desc_12_data_host_addr_3_addr[31:0])
		 ,.int_desc_12_wstrb_host_addr_0_addr(int_desc_12_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_12_wstrb_host_addr_1_addr(int_desc_12_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_12_wstrb_host_addr_2_addr(int_desc_12_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_12_wstrb_host_addr_3_addr(int_desc_12_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_13_data_host_addr_0_addr(int_desc_13_data_host_addr_0_addr[31:0])
		 ,.int_desc_13_data_host_addr_1_addr(int_desc_13_data_host_addr_1_addr[31:0])
		 ,.int_desc_13_data_host_addr_2_addr(int_desc_13_data_host_addr_2_addr[31:0])
		 ,.int_desc_13_data_host_addr_3_addr(int_desc_13_data_host_addr_3_addr[31:0])
		 ,.int_desc_13_wstrb_host_addr_0_addr(int_desc_13_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_13_wstrb_host_addr_1_addr(int_desc_13_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_13_wstrb_host_addr_2_addr(int_desc_13_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_13_wstrb_host_addr_3_addr(int_desc_13_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_14_data_host_addr_0_addr(int_desc_14_data_host_addr_0_addr[31:0])
		 ,.int_desc_14_data_host_addr_1_addr(int_desc_14_data_host_addr_1_addr[31:0])
		 ,.int_desc_14_data_host_addr_2_addr(int_desc_14_data_host_addr_2_addr[31:0])
		 ,.int_desc_14_data_host_addr_3_addr(int_desc_14_data_host_addr_3_addr[31:0])
		 ,.int_desc_14_wstrb_host_addr_0_addr(int_desc_14_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_14_wstrb_host_addr_1_addr(int_desc_14_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_14_wstrb_host_addr_2_addr(int_desc_14_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_14_wstrb_host_addr_3_addr(int_desc_14_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_15_data_host_addr_0_addr(int_desc_15_data_host_addr_0_addr[31:0])
		 ,.int_desc_15_data_host_addr_1_addr(int_desc_15_data_host_addr_1_addr[31:0])
		 ,.int_desc_15_data_host_addr_2_addr(int_desc_15_data_host_addr_2_addr[31:0])
		 ,.int_desc_15_data_host_addr_3_addr(int_desc_15_data_host_addr_3_addr[31:0])
		 ,.int_desc_15_wstrb_host_addr_0_addr(int_desc_15_wstrb_host_addr_0_addr[31:0])
		 ,.int_desc_15_wstrb_host_addr_1_addr(int_desc_15_wstrb_host_addr_1_addr[31:0])
		 ,.int_desc_15_wstrb_host_addr_2_addr(int_desc_15_wstrb_host_addr_2_addr[31:0])
		 ,.int_desc_15_wstrb_host_addr_3_addr(int_desc_15_wstrb_host_addr_3_addr[31:0])
		 ,.int_desc_0_xuser_0_xuser(int_desc_0_xuser_0_xuser[31:0])
		 ,.int_desc_0_xuser_1_xuser(int_desc_0_xuser_1_xuser[31:0])
		 ,.int_desc_0_xuser_2_xuser(int_desc_0_xuser_2_xuser[31:0])
		 ,.int_desc_0_xuser_3_xuser(int_desc_0_xuser_3_xuser[31:0])
		 ,.int_desc_0_xuser_4_xuser(int_desc_0_xuser_4_xuser[31:0])
		 ,.int_desc_0_xuser_5_xuser(int_desc_0_xuser_5_xuser[31:0])
		 ,.int_desc_0_xuser_6_xuser(int_desc_0_xuser_6_xuser[31:0])
		 ,.int_desc_0_xuser_7_xuser(int_desc_0_xuser_7_xuser[31:0])
		 ,.int_desc_0_xuser_8_xuser(int_desc_0_xuser_8_xuser[31:0])
		 ,.int_desc_0_xuser_9_xuser(int_desc_0_xuser_9_xuser[31:0])
		 ,.int_desc_0_xuser_10_xuser(int_desc_0_xuser_10_xuser[31:0])
		 ,.int_desc_0_xuser_11_xuser(int_desc_0_xuser_11_xuser[31:0])
		 ,.int_desc_0_xuser_12_xuser(int_desc_0_xuser_12_xuser[31:0])
		 ,.int_desc_0_xuser_13_xuser(int_desc_0_xuser_13_xuser[31:0])
		 ,.int_desc_0_xuser_14_xuser(int_desc_0_xuser_14_xuser[31:0])
		 ,.int_desc_0_xuser_15_xuser(int_desc_0_xuser_15_xuser[31:0])
		 ,.int_desc_1_xuser_0_xuser(int_desc_1_xuser_0_xuser[31:0])
		 ,.int_desc_1_xuser_1_xuser(int_desc_1_xuser_1_xuser[31:0])
		 ,.int_desc_1_xuser_2_xuser(int_desc_1_xuser_2_xuser[31:0])
		 ,.int_desc_1_xuser_3_xuser(int_desc_1_xuser_3_xuser[31:0])
		 ,.int_desc_1_xuser_4_xuser(int_desc_1_xuser_4_xuser[31:0])
		 ,.int_desc_1_xuser_5_xuser(int_desc_1_xuser_5_xuser[31:0])
		 ,.int_desc_1_xuser_6_xuser(int_desc_1_xuser_6_xuser[31:0])
		 ,.int_desc_1_xuser_7_xuser(int_desc_1_xuser_7_xuser[31:0])
		 ,.int_desc_1_xuser_8_xuser(int_desc_1_xuser_8_xuser[31:0])
		 ,.int_desc_1_xuser_9_xuser(int_desc_1_xuser_9_xuser[31:0])
		 ,.int_desc_1_xuser_10_xuser(int_desc_1_xuser_10_xuser[31:0])
		 ,.int_desc_1_xuser_11_xuser(int_desc_1_xuser_11_xuser[31:0])
		 ,.int_desc_1_xuser_12_xuser(int_desc_1_xuser_12_xuser[31:0])
		 ,.int_desc_1_xuser_13_xuser(int_desc_1_xuser_13_xuser[31:0])
		 ,.int_desc_1_xuser_14_xuser(int_desc_1_xuser_14_xuser[31:0])
		 ,.int_desc_1_xuser_15_xuser(int_desc_1_xuser_15_xuser[31:0])
		 ,.int_desc_2_xuser_0_xuser(int_desc_2_xuser_0_xuser[31:0])
		 ,.int_desc_2_xuser_1_xuser(int_desc_2_xuser_1_xuser[31:0])
		 ,.int_desc_2_xuser_2_xuser(int_desc_2_xuser_2_xuser[31:0])
		 ,.int_desc_2_xuser_3_xuser(int_desc_2_xuser_3_xuser[31:0])
		 ,.int_desc_2_xuser_4_xuser(int_desc_2_xuser_4_xuser[31:0])
		 ,.int_desc_2_xuser_5_xuser(int_desc_2_xuser_5_xuser[31:0])
		 ,.int_desc_2_xuser_6_xuser(int_desc_2_xuser_6_xuser[31:0])
		 ,.int_desc_2_xuser_7_xuser(int_desc_2_xuser_7_xuser[31:0])
		 ,.int_desc_2_xuser_8_xuser(int_desc_2_xuser_8_xuser[31:0])
		 ,.int_desc_2_xuser_9_xuser(int_desc_2_xuser_9_xuser[31:0])
		 ,.int_desc_2_xuser_10_xuser(int_desc_2_xuser_10_xuser[31:0])
		 ,.int_desc_2_xuser_11_xuser(int_desc_2_xuser_11_xuser[31:0])
		 ,.int_desc_2_xuser_12_xuser(int_desc_2_xuser_12_xuser[31:0])
		 ,.int_desc_2_xuser_13_xuser(int_desc_2_xuser_13_xuser[31:0])
		 ,.int_desc_2_xuser_14_xuser(int_desc_2_xuser_14_xuser[31:0])
		 ,.int_desc_2_xuser_15_xuser(int_desc_2_xuser_15_xuser[31:0])
		 ,.int_desc_3_xuser_0_xuser(int_desc_3_xuser_0_xuser[31:0])
		 ,.int_desc_3_xuser_1_xuser(int_desc_3_xuser_1_xuser[31:0])
		 ,.int_desc_3_xuser_2_xuser(int_desc_3_xuser_2_xuser[31:0])
		 ,.int_desc_3_xuser_3_xuser(int_desc_3_xuser_3_xuser[31:0])
		 ,.int_desc_3_xuser_4_xuser(int_desc_3_xuser_4_xuser[31:0])
		 ,.int_desc_3_xuser_5_xuser(int_desc_3_xuser_5_xuser[31:0])
		 ,.int_desc_3_xuser_6_xuser(int_desc_3_xuser_6_xuser[31:0])
		 ,.int_desc_3_xuser_7_xuser(int_desc_3_xuser_7_xuser[31:0])
		 ,.int_desc_3_xuser_8_xuser(int_desc_3_xuser_8_xuser[31:0])
		 ,.int_desc_3_xuser_9_xuser(int_desc_3_xuser_9_xuser[31:0])
		 ,.int_desc_3_xuser_10_xuser(int_desc_3_xuser_10_xuser[31:0])
		 ,.int_desc_3_xuser_11_xuser(int_desc_3_xuser_11_xuser[31:0])
		 ,.int_desc_3_xuser_12_xuser(int_desc_3_xuser_12_xuser[31:0])
		 ,.int_desc_3_xuser_13_xuser(int_desc_3_xuser_13_xuser[31:0])
		 ,.int_desc_3_xuser_14_xuser(int_desc_3_xuser_14_xuser[31:0])
		 ,.int_desc_3_xuser_15_xuser(int_desc_3_xuser_15_xuser[31:0])
		 ,.int_desc_4_xuser_0_xuser(int_desc_4_xuser_0_xuser[31:0])
		 ,.int_desc_4_xuser_1_xuser(int_desc_4_xuser_1_xuser[31:0])
		 ,.int_desc_4_xuser_2_xuser(int_desc_4_xuser_2_xuser[31:0])
		 ,.int_desc_4_xuser_3_xuser(int_desc_4_xuser_3_xuser[31:0])
		 ,.int_desc_4_xuser_4_xuser(int_desc_4_xuser_4_xuser[31:0])
		 ,.int_desc_4_xuser_5_xuser(int_desc_4_xuser_5_xuser[31:0])
		 ,.int_desc_4_xuser_6_xuser(int_desc_4_xuser_6_xuser[31:0])
		 ,.int_desc_4_xuser_7_xuser(int_desc_4_xuser_7_xuser[31:0])
		 ,.int_desc_4_xuser_8_xuser(int_desc_4_xuser_8_xuser[31:0])
		 ,.int_desc_4_xuser_9_xuser(int_desc_4_xuser_9_xuser[31:0])
		 ,.int_desc_4_xuser_10_xuser(int_desc_4_xuser_10_xuser[31:0])
		 ,.int_desc_4_xuser_11_xuser(int_desc_4_xuser_11_xuser[31:0])
		 ,.int_desc_4_xuser_12_xuser(int_desc_4_xuser_12_xuser[31:0])
		 ,.int_desc_4_xuser_13_xuser(int_desc_4_xuser_13_xuser[31:0])
		 ,.int_desc_4_xuser_14_xuser(int_desc_4_xuser_14_xuser[31:0])
		 ,.int_desc_4_xuser_15_xuser(int_desc_4_xuser_15_xuser[31:0])
		 ,.int_desc_5_xuser_0_xuser(int_desc_5_xuser_0_xuser[31:0])
		 ,.int_desc_5_xuser_1_xuser(int_desc_5_xuser_1_xuser[31:0])
		 ,.int_desc_5_xuser_2_xuser(int_desc_5_xuser_2_xuser[31:0])
		 ,.int_desc_5_xuser_3_xuser(int_desc_5_xuser_3_xuser[31:0])
		 ,.int_desc_5_xuser_4_xuser(int_desc_5_xuser_4_xuser[31:0])
		 ,.int_desc_5_xuser_5_xuser(int_desc_5_xuser_5_xuser[31:0])
		 ,.int_desc_5_xuser_6_xuser(int_desc_5_xuser_6_xuser[31:0])
		 ,.int_desc_5_xuser_7_xuser(int_desc_5_xuser_7_xuser[31:0])
		 ,.int_desc_5_xuser_8_xuser(int_desc_5_xuser_8_xuser[31:0])
		 ,.int_desc_5_xuser_9_xuser(int_desc_5_xuser_9_xuser[31:0])
		 ,.int_desc_5_xuser_10_xuser(int_desc_5_xuser_10_xuser[31:0])
		 ,.int_desc_5_xuser_11_xuser(int_desc_5_xuser_11_xuser[31:0])
		 ,.int_desc_5_xuser_12_xuser(int_desc_5_xuser_12_xuser[31:0])
		 ,.int_desc_5_xuser_13_xuser(int_desc_5_xuser_13_xuser[31:0])
		 ,.int_desc_5_xuser_14_xuser(int_desc_5_xuser_14_xuser[31:0])
		 ,.int_desc_5_xuser_15_xuser(int_desc_5_xuser_15_xuser[31:0])
		 ,.int_desc_6_xuser_0_xuser(int_desc_6_xuser_0_xuser[31:0])
		 ,.int_desc_6_xuser_1_xuser(int_desc_6_xuser_1_xuser[31:0])
		 ,.int_desc_6_xuser_2_xuser(int_desc_6_xuser_2_xuser[31:0])
		 ,.int_desc_6_xuser_3_xuser(int_desc_6_xuser_3_xuser[31:0])
		 ,.int_desc_6_xuser_4_xuser(int_desc_6_xuser_4_xuser[31:0])
		 ,.int_desc_6_xuser_5_xuser(int_desc_6_xuser_5_xuser[31:0])
		 ,.int_desc_6_xuser_6_xuser(int_desc_6_xuser_6_xuser[31:0])
		 ,.int_desc_6_xuser_7_xuser(int_desc_6_xuser_7_xuser[31:0])
		 ,.int_desc_6_xuser_8_xuser(int_desc_6_xuser_8_xuser[31:0])
		 ,.int_desc_6_xuser_9_xuser(int_desc_6_xuser_9_xuser[31:0])
		 ,.int_desc_6_xuser_10_xuser(int_desc_6_xuser_10_xuser[31:0])
		 ,.int_desc_6_xuser_11_xuser(int_desc_6_xuser_11_xuser[31:0])
		 ,.int_desc_6_xuser_12_xuser(int_desc_6_xuser_12_xuser[31:0])
		 ,.int_desc_6_xuser_13_xuser(int_desc_6_xuser_13_xuser[31:0])
		 ,.int_desc_6_xuser_14_xuser(int_desc_6_xuser_14_xuser[31:0])
		 ,.int_desc_6_xuser_15_xuser(int_desc_6_xuser_15_xuser[31:0])
		 ,.int_desc_7_xuser_0_xuser(int_desc_7_xuser_0_xuser[31:0])
		 ,.int_desc_7_xuser_1_xuser(int_desc_7_xuser_1_xuser[31:0])
		 ,.int_desc_7_xuser_2_xuser(int_desc_7_xuser_2_xuser[31:0])
		 ,.int_desc_7_xuser_3_xuser(int_desc_7_xuser_3_xuser[31:0])
		 ,.int_desc_7_xuser_4_xuser(int_desc_7_xuser_4_xuser[31:0])
		 ,.int_desc_7_xuser_5_xuser(int_desc_7_xuser_5_xuser[31:0])
		 ,.int_desc_7_xuser_6_xuser(int_desc_7_xuser_6_xuser[31:0])
		 ,.int_desc_7_xuser_7_xuser(int_desc_7_xuser_7_xuser[31:0])
		 ,.int_desc_7_xuser_8_xuser(int_desc_7_xuser_8_xuser[31:0])
		 ,.int_desc_7_xuser_9_xuser(int_desc_7_xuser_9_xuser[31:0])
		 ,.int_desc_7_xuser_10_xuser(int_desc_7_xuser_10_xuser[31:0])
		 ,.int_desc_7_xuser_11_xuser(int_desc_7_xuser_11_xuser[31:0])
		 ,.int_desc_7_xuser_12_xuser(int_desc_7_xuser_12_xuser[31:0])
		 ,.int_desc_7_xuser_13_xuser(int_desc_7_xuser_13_xuser[31:0])
		 ,.int_desc_7_xuser_14_xuser(int_desc_7_xuser_14_xuser[31:0])
		 ,.int_desc_7_xuser_15_xuser(int_desc_7_xuser_15_xuser[31:0])
		 ,.int_desc_8_xuser_0_xuser(int_desc_8_xuser_0_xuser[31:0])
		 ,.int_desc_8_xuser_1_xuser(int_desc_8_xuser_1_xuser[31:0])
		 ,.int_desc_8_xuser_2_xuser(int_desc_8_xuser_2_xuser[31:0])
		 ,.int_desc_8_xuser_3_xuser(int_desc_8_xuser_3_xuser[31:0])
		 ,.int_desc_8_xuser_4_xuser(int_desc_8_xuser_4_xuser[31:0])
		 ,.int_desc_8_xuser_5_xuser(int_desc_8_xuser_5_xuser[31:0])
		 ,.int_desc_8_xuser_6_xuser(int_desc_8_xuser_6_xuser[31:0])
		 ,.int_desc_8_xuser_7_xuser(int_desc_8_xuser_7_xuser[31:0])
		 ,.int_desc_8_xuser_8_xuser(int_desc_8_xuser_8_xuser[31:0])
		 ,.int_desc_8_xuser_9_xuser(int_desc_8_xuser_9_xuser[31:0])
		 ,.int_desc_8_xuser_10_xuser(int_desc_8_xuser_10_xuser[31:0])
		 ,.int_desc_8_xuser_11_xuser(int_desc_8_xuser_11_xuser[31:0])
		 ,.int_desc_8_xuser_12_xuser(int_desc_8_xuser_12_xuser[31:0])
		 ,.int_desc_8_xuser_13_xuser(int_desc_8_xuser_13_xuser[31:0])
		 ,.int_desc_8_xuser_14_xuser(int_desc_8_xuser_14_xuser[31:0])
		 ,.int_desc_8_xuser_15_xuser(int_desc_8_xuser_15_xuser[31:0])
		 ,.int_desc_9_xuser_0_xuser(int_desc_9_xuser_0_xuser[31:0])
		 ,.int_desc_9_xuser_1_xuser(int_desc_9_xuser_1_xuser[31:0])
		 ,.int_desc_9_xuser_2_xuser(int_desc_9_xuser_2_xuser[31:0])
		 ,.int_desc_9_xuser_3_xuser(int_desc_9_xuser_3_xuser[31:0])
		 ,.int_desc_9_xuser_4_xuser(int_desc_9_xuser_4_xuser[31:0])
		 ,.int_desc_9_xuser_5_xuser(int_desc_9_xuser_5_xuser[31:0])
		 ,.int_desc_9_xuser_6_xuser(int_desc_9_xuser_6_xuser[31:0])
		 ,.int_desc_9_xuser_7_xuser(int_desc_9_xuser_7_xuser[31:0])
		 ,.int_desc_9_xuser_8_xuser(int_desc_9_xuser_8_xuser[31:0])
		 ,.int_desc_9_xuser_9_xuser(int_desc_9_xuser_9_xuser[31:0])
		 ,.int_desc_9_xuser_10_xuser(int_desc_9_xuser_10_xuser[31:0])
		 ,.int_desc_9_xuser_11_xuser(int_desc_9_xuser_11_xuser[31:0])
		 ,.int_desc_9_xuser_12_xuser(int_desc_9_xuser_12_xuser[31:0])
		 ,.int_desc_9_xuser_13_xuser(int_desc_9_xuser_13_xuser[31:0])
		 ,.int_desc_9_xuser_14_xuser(int_desc_9_xuser_14_xuser[31:0])
		 ,.int_desc_9_xuser_15_xuser(int_desc_9_xuser_15_xuser[31:0])
		 ,.int_desc_10_xuser_0_xuser(int_desc_10_xuser_0_xuser[31:0])
		 ,.int_desc_10_xuser_1_xuser(int_desc_10_xuser_1_xuser[31:0])
		 ,.int_desc_10_xuser_2_xuser(int_desc_10_xuser_2_xuser[31:0])
		 ,.int_desc_10_xuser_3_xuser(int_desc_10_xuser_3_xuser[31:0])
		 ,.int_desc_10_xuser_4_xuser(int_desc_10_xuser_4_xuser[31:0])
		 ,.int_desc_10_xuser_5_xuser(int_desc_10_xuser_5_xuser[31:0])
		 ,.int_desc_10_xuser_6_xuser(int_desc_10_xuser_6_xuser[31:0])
		 ,.int_desc_10_xuser_7_xuser(int_desc_10_xuser_7_xuser[31:0])
		 ,.int_desc_10_xuser_8_xuser(int_desc_10_xuser_8_xuser[31:0])
		 ,.int_desc_10_xuser_9_xuser(int_desc_10_xuser_9_xuser[31:0])
		 ,.int_desc_10_xuser_10_xuser(int_desc_10_xuser_10_xuser[31:0])
		 ,.int_desc_10_xuser_11_xuser(int_desc_10_xuser_11_xuser[31:0])
		 ,.int_desc_10_xuser_12_xuser(int_desc_10_xuser_12_xuser[31:0])
		 ,.int_desc_10_xuser_13_xuser(int_desc_10_xuser_13_xuser[31:0])
		 ,.int_desc_10_xuser_14_xuser(int_desc_10_xuser_14_xuser[31:0])
		 ,.int_desc_10_xuser_15_xuser(int_desc_10_xuser_15_xuser[31:0])
		 ,.int_desc_11_xuser_0_xuser(int_desc_11_xuser_0_xuser[31:0])
		 ,.int_desc_11_xuser_1_xuser(int_desc_11_xuser_1_xuser[31:0])
		 ,.int_desc_11_xuser_2_xuser(int_desc_11_xuser_2_xuser[31:0])
		 ,.int_desc_11_xuser_3_xuser(int_desc_11_xuser_3_xuser[31:0])
		 ,.int_desc_11_xuser_4_xuser(int_desc_11_xuser_4_xuser[31:0])
		 ,.int_desc_11_xuser_5_xuser(int_desc_11_xuser_5_xuser[31:0])
		 ,.int_desc_11_xuser_6_xuser(int_desc_11_xuser_6_xuser[31:0])
		 ,.int_desc_11_xuser_7_xuser(int_desc_11_xuser_7_xuser[31:0])
		 ,.int_desc_11_xuser_8_xuser(int_desc_11_xuser_8_xuser[31:0])
		 ,.int_desc_11_xuser_9_xuser(int_desc_11_xuser_9_xuser[31:0])
		 ,.int_desc_11_xuser_10_xuser(int_desc_11_xuser_10_xuser[31:0])
		 ,.int_desc_11_xuser_11_xuser(int_desc_11_xuser_11_xuser[31:0])
		 ,.int_desc_11_xuser_12_xuser(int_desc_11_xuser_12_xuser[31:0])
		 ,.int_desc_11_xuser_13_xuser(int_desc_11_xuser_13_xuser[31:0])
		 ,.int_desc_11_xuser_14_xuser(int_desc_11_xuser_14_xuser[31:0])
		 ,.int_desc_11_xuser_15_xuser(int_desc_11_xuser_15_xuser[31:0])
		 ,.int_desc_12_xuser_0_xuser(int_desc_12_xuser_0_xuser[31:0])
		 ,.int_desc_12_xuser_1_xuser(int_desc_12_xuser_1_xuser[31:0])
		 ,.int_desc_12_xuser_2_xuser(int_desc_12_xuser_2_xuser[31:0])
		 ,.int_desc_12_xuser_3_xuser(int_desc_12_xuser_3_xuser[31:0])
		 ,.int_desc_12_xuser_4_xuser(int_desc_12_xuser_4_xuser[31:0])
		 ,.int_desc_12_xuser_5_xuser(int_desc_12_xuser_5_xuser[31:0])
		 ,.int_desc_12_xuser_6_xuser(int_desc_12_xuser_6_xuser[31:0])
		 ,.int_desc_12_xuser_7_xuser(int_desc_12_xuser_7_xuser[31:0])
		 ,.int_desc_12_xuser_8_xuser(int_desc_12_xuser_8_xuser[31:0])
		 ,.int_desc_12_xuser_9_xuser(int_desc_12_xuser_9_xuser[31:0])
		 ,.int_desc_12_xuser_10_xuser(int_desc_12_xuser_10_xuser[31:0])
		 ,.int_desc_12_xuser_11_xuser(int_desc_12_xuser_11_xuser[31:0])
		 ,.int_desc_12_xuser_12_xuser(int_desc_12_xuser_12_xuser[31:0])
		 ,.int_desc_12_xuser_13_xuser(int_desc_12_xuser_13_xuser[31:0])
		 ,.int_desc_12_xuser_14_xuser(int_desc_12_xuser_14_xuser[31:0])
		 ,.int_desc_12_xuser_15_xuser(int_desc_12_xuser_15_xuser[31:0])
		 ,.int_desc_13_xuser_0_xuser(int_desc_13_xuser_0_xuser[31:0])
		 ,.int_desc_13_xuser_1_xuser(int_desc_13_xuser_1_xuser[31:0])
		 ,.int_desc_13_xuser_2_xuser(int_desc_13_xuser_2_xuser[31:0])
		 ,.int_desc_13_xuser_3_xuser(int_desc_13_xuser_3_xuser[31:0])
		 ,.int_desc_13_xuser_4_xuser(int_desc_13_xuser_4_xuser[31:0])
		 ,.int_desc_13_xuser_5_xuser(int_desc_13_xuser_5_xuser[31:0])
		 ,.int_desc_13_xuser_6_xuser(int_desc_13_xuser_6_xuser[31:0])
		 ,.int_desc_13_xuser_7_xuser(int_desc_13_xuser_7_xuser[31:0])
		 ,.int_desc_13_xuser_8_xuser(int_desc_13_xuser_8_xuser[31:0])
		 ,.int_desc_13_xuser_9_xuser(int_desc_13_xuser_9_xuser[31:0])
		 ,.int_desc_13_xuser_10_xuser(int_desc_13_xuser_10_xuser[31:0])
		 ,.int_desc_13_xuser_11_xuser(int_desc_13_xuser_11_xuser[31:0])
		 ,.int_desc_13_xuser_12_xuser(int_desc_13_xuser_12_xuser[31:0])
		 ,.int_desc_13_xuser_13_xuser(int_desc_13_xuser_13_xuser[31:0])
		 ,.int_desc_13_xuser_14_xuser(int_desc_13_xuser_14_xuser[31:0])
		 ,.int_desc_13_xuser_15_xuser(int_desc_13_xuser_15_xuser[31:0])
		 ,.int_desc_14_xuser_0_xuser(int_desc_14_xuser_0_xuser[31:0])
		 ,.int_desc_14_xuser_1_xuser(int_desc_14_xuser_1_xuser[31:0])
		 ,.int_desc_14_xuser_2_xuser(int_desc_14_xuser_2_xuser[31:0])
		 ,.int_desc_14_xuser_3_xuser(int_desc_14_xuser_3_xuser[31:0])
		 ,.int_desc_14_xuser_4_xuser(int_desc_14_xuser_4_xuser[31:0])
		 ,.int_desc_14_xuser_5_xuser(int_desc_14_xuser_5_xuser[31:0])
		 ,.int_desc_14_xuser_6_xuser(int_desc_14_xuser_6_xuser[31:0])
		 ,.int_desc_14_xuser_7_xuser(int_desc_14_xuser_7_xuser[31:0])
		 ,.int_desc_14_xuser_8_xuser(int_desc_14_xuser_8_xuser[31:0])
		 ,.int_desc_14_xuser_9_xuser(int_desc_14_xuser_9_xuser[31:0])
		 ,.int_desc_14_xuser_10_xuser(int_desc_14_xuser_10_xuser[31:0])
		 ,.int_desc_14_xuser_11_xuser(int_desc_14_xuser_11_xuser[31:0])
		 ,.int_desc_14_xuser_12_xuser(int_desc_14_xuser_12_xuser[31:0])
		 ,.int_desc_14_xuser_13_xuser(int_desc_14_xuser_13_xuser[31:0])
		 ,.int_desc_14_xuser_14_xuser(int_desc_14_xuser_14_xuser[31:0])
		 ,.int_desc_14_xuser_15_xuser(int_desc_14_xuser_15_xuser[31:0])
		 ,.int_desc_15_xuser_0_xuser(int_desc_15_xuser_0_xuser[31:0])
		 ,.int_desc_15_xuser_1_xuser(int_desc_15_xuser_1_xuser[31:0])
		 ,.int_desc_15_xuser_2_xuser(int_desc_15_xuser_2_xuser[31:0])
		 ,.int_desc_15_xuser_3_xuser(int_desc_15_xuser_3_xuser[31:0])
		 ,.int_desc_15_xuser_4_xuser(int_desc_15_xuser_4_xuser[31:0])
		 ,.int_desc_15_xuser_5_xuser(int_desc_15_xuser_5_xuser[31:0])
		 ,.int_desc_15_xuser_6_xuser(int_desc_15_xuser_6_xuser[31:0])
		 ,.int_desc_15_xuser_7_xuser(int_desc_15_xuser_7_xuser[31:0])
		 ,.int_desc_15_xuser_8_xuser(int_desc_15_xuser_8_xuser[31:0])
		 ,.int_desc_15_xuser_9_xuser(int_desc_15_xuser_9_xuser[31:0])
		 ,.int_desc_15_xuser_10_xuser(int_desc_15_xuser_10_xuser[31:0])
		 ,.int_desc_15_xuser_11_xuser(int_desc_15_xuser_11_xuser[31:0])
		 ,.int_desc_15_xuser_12_xuser(int_desc_15_xuser_12_xuser[31:0])
		 ,.int_desc_15_xuser_13_xuser(int_desc_15_xuser_13_xuser[31:0])
		 ,.int_desc_15_xuser_14_xuser(int_desc_15_xuser_14_xuser[31:0])
		 ,.int_desc_15_xuser_15_xuser(int_desc_15_xuser_15_xuser[31:0])
		  
   
