/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */

        ,input [0:0]	int_desc_0_txn_type_wr_strb
        ,input [0:0]	int_desc_0_txn_type_wr_rd
        ,input [3:0]	int_desc_0_attr_axregion
        ,input [3:0]	int_desc_0_attr_axqos
        ,input [2:0]	int_desc_0_attr_axprot
        ,input [3:0]	int_desc_0_attr_axcache
        ,input [1:0]	int_desc_0_attr_axlock
        ,input [1:0]	int_desc_0_attr_axburst
        ,input [31:0]	int_desc_0_axid_0_axid
        ,input [31:0]	int_desc_0_axid_1_axid
        ,input [31:0]	int_desc_0_axid_2_axid
        ,input [31:0]	int_desc_0_axid_3_axid
        ,input [31:0]	int_desc_0_axuser_0_axuser
        ,input [31:0]	int_desc_0_axuser_1_axuser
        ,input [31:0]	int_desc_0_axuser_2_axuser
        ,input [31:0]	int_desc_0_axuser_3_axuser
        ,input [31:0]	int_desc_0_axuser_4_axuser
        ,input [31:0]	int_desc_0_axuser_5_axuser
        ,input [31:0]	int_desc_0_axuser_6_axuser
        ,input [31:0]	int_desc_0_axuser_7_axuser
        ,input [31:0]	int_desc_0_axuser_8_axuser
        ,input [31:0]	int_desc_0_axuser_9_axuser
        ,input [31:0]	int_desc_0_axuser_10_axuser
        ,input [31:0]	int_desc_0_axuser_11_axuser
        ,input [31:0]	int_desc_0_axuser_12_axuser
        ,input [31:0]	int_desc_0_axuser_13_axuser
        ,input [31:0]	int_desc_0_axuser_14_axuser
        ,input [31:0]	int_desc_0_axuser_15_axuser
        ,input [31:0]	int_desc_0_size_txn_size
        ,input [2:0]	int_desc_0_axsize_axsize
        ,input [31:0]	int_desc_0_axaddr_0_addr
        ,input [31:0]	int_desc_0_axaddr_1_addr
        ,input [31:0]	int_desc_0_axaddr_2_addr
        ,input [31:0]	int_desc_0_axaddr_3_addr
        ,input [31:0]	int_desc_0_data_offset_addr
        ,input [31:0]	int_desc_0_wuser_0_wuser
        ,input [31:0]	int_desc_0_wuser_1_wuser
        ,input [31:0]	int_desc_0_wuser_2_wuser
        ,input [31:0]	int_desc_0_wuser_3_wuser
        ,input [31:0]	int_desc_0_wuser_4_wuser
        ,input [31:0]	int_desc_0_wuser_5_wuser
        ,input [31:0]	int_desc_0_wuser_6_wuser
        ,input [31:0]	int_desc_0_wuser_7_wuser
        ,input [31:0]	int_desc_0_wuser_8_wuser
        ,input [31:0]	int_desc_0_wuser_9_wuser
        ,input [31:0]	int_desc_0_wuser_10_wuser
        ,input [31:0]	int_desc_0_wuser_11_wuser
        ,input [31:0]	int_desc_0_wuser_12_wuser
        ,input [31:0]	int_desc_0_wuser_13_wuser
        ,input [31:0]	int_desc_0_wuser_14_wuser
        ,input [31:0]	int_desc_0_wuser_15_wuser
        ,input [0:0]	int_desc_1_txn_type_wr_strb
        ,input [0:0]	int_desc_1_txn_type_wr_rd
        ,input [3:0]	int_desc_1_attr_axregion
        ,input [3:0]	int_desc_1_attr_axqos
        ,input [2:0]	int_desc_1_attr_axprot
        ,input [3:0]	int_desc_1_attr_axcache
        ,input [1:0]	int_desc_1_attr_axlock
        ,input [1:0]	int_desc_1_attr_axburst
        ,input [31:0]	int_desc_1_axid_0_axid
        ,input [31:0]	int_desc_1_axid_1_axid
        ,input [31:0]	int_desc_1_axid_2_axid
        ,input [31:0]	int_desc_1_axid_3_axid
        ,input [31:0]	int_desc_1_axuser_0_axuser
        ,input [31:0]	int_desc_1_axuser_1_axuser
        ,input [31:0]	int_desc_1_axuser_2_axuser
        ,input [31:0]	int_desc_1_axuser_3_axuser
        ,input [31:0]	int_desc_1_axuser_4_axuser
        ,input [31:0]	int_desc_1_axuser_5_axuser
        ,input [31:0]	int_desc_1_axuser_6_axuser
        ,input [31:0]	int_desc_1_axuser_7_axuser
        ,input [31:0]	int_desc_1_axuser_8_axuser
        ,input [31:0]	int_desc_1_axuser_9_axuser
        ,input [31:0]	int_desc_1_axuser_10_axuser
        ,input [31:0]	int_desc_1_axuser_11_axuser
        ,input [31:0]	int_desc_1_axuser_12_axuser
        ,input [31:0]	int_desc_1_axuser_13_axuser
        ,input [31:0]	int_desc_1_axuser_14_axuser
        ,input [31:0]	int_desc_1_axuser_15_axuser
        ,input [31:0]	int_desc_1_size_txn_size
        ,input [2:0]	int_desc_1_axsize_axsize
        ,input [31:0]	int_desc_1_axaddr_0_addr
        ,input [31:0]	int_desc_1_axaddr_1_addr
        ,input [31:0]	int_desc_1_axaddr_2_addr
        ,input [31:0]	int_desc_1_axaddr_3_addr
        ,input [31:0]	int_desc_1_data_offset_addr
        ,input [31:0]	int_desc_1_wuser_0_wuser
        ,input [31:0]	int_desc_1_wuser_1_wuser
        ,input [31:0]	int_desc_1_wuser_2_wuser
        ,input [31:0]	int_desc_1_wuser_3_wuser
        ,input [31:0]	int_desc_1_wuser_4_wuser
        ,input [31:0]	int_desc_1_wuser_5_wuser
        ,input [31:0]	int_desc_1_wuser_6_wuser
        ,input [31:0]	int_desc_1_wuser_7_wuser
        ,input [31:0]	int_desc_1_wuser_8_wuser
        ,input [31:0]	int_desc_1_wuser_9_wuser
        ,input [31:0]	int_desc_1_wuser_10_wuser
        ,input [31:0]	int_desc_1_wuser_11_wuser
        ,input [31:0]	int_desc_1_wuser_12_wuser
        ,input [31:0]	int_desc_1_wuser_13_wuser
        ,input [31:0]	int_desc_1_wuser_14_wuser
        ,input [31:0]	int_desc_1_wuser_15_wuser
        ,input [0:0]	int_desc_2_txn_type_wr_strb
        ,input [0:0]	int_desc_2_txn_type_wr_rd
        ,input [3:0]	int_desc_2_attr_axregion
        ,input [3:0]	int_desc_2_attr_axqos
        ,input [2:0]	int_desc_2_attr_axprot
        ,input [3:0]	int_desc_2_attr_axcache
        ,input [1:0]	int_desc_2_attr_axlock
        ,input [1:0]	int_desc_2_attr_axburst
        ,input [31:0]	int_desc_2_axid_0_axid
        ,input [31:0]	int_desc_2_axid_1_axid
        ,input [31:0]	int_desc_2_axid_2_axid
        ,input [31:0]	int_desc_2_axid_3_axid
        ,input [31:0]	int_desc_2_axuser_0_axuser
        ,input [31:0]	int_desc_2_axuser_1_axuser
        ,input [31:0]	int_desc_2_axuser_2_axuser
        ,input [31:0]	int_desc_2_axuser_3_axuser
        ,input [31:0]	int_desc_2_axuser_4_axuser
        ,input [31:0]	int_desc_2_axuser_5_axuser
        ,input [31:0]	int_desc_2_axuser_6_axuser
        ,input [31:0]	int_desc_2_axuser_7_axuser
        ,input [31:0]	int_desc_2_axuser_8_axuser
        ,input [31:0]	int_desc_2_axuser_9_axuser
        ,input [31:0]	int_desc_2_axuser_10_axuser
        ,input [31:0]	int_desc_2_axuser_11_axuser
        ,input [31:0]	int_desc_2_axuser_12_axuser
        ,input [31:0]	int_desc_2_axuser_13_axuser
        ,input [31:0]	int_desc_2_axuser_14_axuser
        ,input [31:0]	int_desc_2_axuser_15_axuser
        ,input [31:0]	int_desc_2_size_txn_size
        ,input [2:0]	int_desc_2_axsize_axsize
        ,input [31:0]	int_desc_2_axaddr_0_addr
        ,input [31:0]	int_desc_2_axaddr_1_addr
        ,input [31:0]	int_desc_2_axaddr_2_addr
        ,input [31:0]	int_desc_2_axaddr_3_addr
        ,input [31:0]	int_desc_2_data_offset_addr
        ,input [31:0]	int_desc_2_wuser_0_wuser
        ,input [31:0]	int_desc_2_wuser_1_wuser
        ,input [31:0]	int_desc_2_wuser_2_wuser
        ,input [31:0]	int_desc_2_wuser_3_wuser
        ,input [31:0]	int_desc_2_wuser_4_wuser
        ,input [31:0]	int_desc_2_wuser_5_wuser
        ,input [31:0]	int_desc_2_wuser_6_wuser
        ,input [31:0]	int_desc_2_wuser_7_wuser
        ,input [31:0]	int_desc_2_wuser_8_wuser
        ,input [31:0]	int_desc_2_wuser_9_wuser
        ,input [31:0]	int_desc_2_wuser_10_wuser
        ,input [31:0]	int_desc_2_wuser_11_wuser
        ,input [31:0]	int_desc_2_wuser_12_wuser
        ,input [31:0]	int_desc_2_wuser_13_wuser
        ,input [31:0]	int_desc_2_wuser_14_wuser
        ,input [31:0]	int_desc_2_wuser_15_wuser
        ,input [0:0]	int_desc_3_txn_type_wr_strb
        ,input [0:0]	int_desc_3_txn_type_wr_rd
        ,input [3:0]	int_desc_3_attr_axregion
        ,input [3:0]	int_desc_3_attr_axqos
        ,input [2:0]	int_desc_3_attr_axprot
        ,input [3:0]	int_desc_3_attr_axcache
        ,input [1:0]	int_desc_3_attr_axlock
        ,input [1:0]	int_desc_3_attr_axburst
        ,input [31:0]	int_desc_3_axid_0_axid
        ,input [31:0]	int_desc_3_axid_1_axid
        ,input [31:0]	int_desc_3_axid_2_axid
        ,input [31:0]	int_desc_3_axid_3_axid
        ,input [31:0]	int_desc_3_axuser_0_axuser
        ,input [31:0]	int_desc_3_axuser_1_axuser
        ,input [31:0]	int_desc_3_axuser_2_axuser
        ,input [31:0]	int_desc_3_axuser_3_axuser
        ,input [31:0]	int_desc_3_axuser_4_axuser
        ,input [31:0]	int_desc_3_axuser_5_axuser
        ,input [31:0]	int_desc_3_axuser_6_axuser
        ,input [31:0]	int_desc_3_axuser_7_axuser
        ,input [31:0]	int_desc_3_axuser_8_axuser
        ,input [31:0]	int_desc_3_axuser_9_axuser
        ,input [31:0]	int_desc_3_axuser_10_axuser
        ,input [31:0]	int_desc_3_axuser_11_axuser
        ,input [31:0]	int_desc_3_axuser_12_axuser
        ,input [31:0]	int_desc_3_axuser_13_axuser
        ,input [31:0]	int_desc_3_axuser_14_axuser
        ,input [31:0]	int_desc_3_axuser_15_axuser
        ,input [31:0]	int_desc_3_size_txn_size
        ,input [2:0]	int_desc_3_axsize_axsize
        ,input [31:0]	int_desc_3_axaddr_0_addr
        ,input [31:0]	int_desc_3_axaddr_1_addr
        ,input [31:0]	int_desc_3_axaddr_2_addr
        ,input [31:0]	int_desc_3_axaddr_3_addr
        ,input [31:0]	int_desc_3_data_offset_addr
        ,input [31:0]	int_desc_3_wuser_0_wuser
        ,input [31:0]	int_desc_3_wuser_1_wuser
        ,input [31:0]	int_desc_3_wuser_2_wuser
        ,input [31:0]	int_desc_3_wuser_3_wuser
        ,input [31:0]	int_desc_3_wuser_4_wuser
        ,input [31:0]	int_desc_3_wuser_5_wuser
        ,input [31:0]	int_desc_3_wuser_6_wuser
        ,input [31:0]	int_desc_3_wuser_7_wuser
        ,input [31:0]	int_desc_3_wuser_8_wuser
        ,input [31:0]	int_desc_3_wuser_9_wuser
        ,input [31:0]	int_desc_3_wuser_10_wuser
        ,input [31:0]	int_desc_3_wuser_11_wuser
        ,input [31:0]	int_desc_3_wuser_12_wuser
        ,input [31:0]	int_desc_3_wuser_13_wuser
        ,input [31:0]	int_desc_3_wuser_14_wuser
        ,input [31:0]	int_desc_3_wuser_15_wuser
        ,input [0:0]	int_desc_4_txn_type_wr_strb
        ,input [0:0]	int_desc_4_txn_type_wr_rd
        ,input [3:0]	int_desc_4_attr_axregion
        ,input [3:0]	int_desc_4_attr_axqos
        ,input [2:0]	int_desc_4_attr_axprot
        ,input [3:0]	int_desc_4_attr_axcache
        ,input [1:0]	int_desc_4_attr_axlock
        ,input [1:0]	int_desc_4_attr_axburst
        ,input [31:0]	int_desc_4_axid_0_axid
        ,input [31:0]	int_desc_4_axid_1_axid
        ,input [31:0]	int_desc_4_axid_2_axid
        ,input [31:0]	int_desc_4_axid_3_axid
        ,input [31:0]	int_desc_4_axuser_0_axuser
        ,input [31:0]	int_desc_4_axuser_1_axuser
        ,input [31:0]	int_desc_4_axuser_2_axuser
        ,input [31:0]	int_desc_4_axuser_3_axuser
        ,input [31:0]	int_desc_4_axuser_4_axuser
        ,input [31:0]	int_desc_4_axuser_5_axuser
        ,input [31:0]	int_desc_4_axuser_6_axuser
        ,input [31:0]	int_desc_4_axuser_7_axuser
        ,input [31:0]	int_desc_4_axuser_8_axuser
        ,input [31:0]	int_desc_4_axuser_9_axuser
        ,input [31:0]	int_desc_4_axuser_10_axuser
        ,input [31:0]	int_desc_4_axuser_11_axuser
        ,input [31:0]	int_desc_4_axuser_12_axuser
        ,input [31:0]	int_desc_4_axuser_13_axuser
        ,input [31:0]	int_desc_4_axuser_14_axuser
        ,input [31:0]	int_desc_4_axuser_15_axuser
        ,input [31:0]	int_desc_4_size_txn_size
        ,input [2:0]	int_desc_4_axsize_axsize
        ,input [31:0]	int_desc_4_axaddr_0_addr
        ,input [31:0]	int_desc_4_axaddr_1_addr
        ,input [31:0]	int_desc_4_axaddr_2_addr
        ,input [31:0]	int_desc_4_axaddr_3_addr
        ,input [31:0]	int_desc_4_data_offset_addr
        ,input [31:0]	int_desc_4_wuser_0_wuser
        ,input [31:0]	int_desc_4_wuser_1_wuser
        ,input [31:0]	int_desc_4_wuser_2_wuser
        ,input [31:0]	int_desc_4_wuser_3_wuser
        ,input [31:0]	int_desc_4_wuser_4_wuser
        ,input [31:0]	int_desc_4_wuser_5_wuser
        ,input [31:0]	int_desc_4_wuser_6_wuser
        ,input [31:0]	int_desc_4_wuser_7_wuser
        ,input [31:0]	int_desc_4_wuser_8_wuser
        ,input [31:0]	int_desc_4_wuser_9_wuser
        ,input [31:0]	int_desc_4_wuser_10_wuser
        ,input [31:0]	int_desc_4_wuser_11_wuser
        ,input [31:0]	int_desc_4_wuser_12_wuser
        ,input [31:0]	int_desc_4_wuser_13_wuser
        ,input [31:0]	int_desc_4_wuser_14_wuser
        ,input [31:0]	int_desc_4_wuser_15_wuser
        ,input [0:0]	int_desc_5_txn_type_wr_strb
        ,input [0:0]	int_desc_5_txn_type_wr_rd
        ,input [3:0]	int_desc_5_attr_axregion
        ,input [3:0]	int_desc_5_attr_axqos
        ,input [2:0]	int_desc_5_attr_axprot
        ,input [3:0]	int_desc_5_attr_axcache
        ,input [1:0]	int_desc_5_attr_axlock
        ,input [1:0]	int_desc_5_attr_axburst
        ,input [31:0]	int_desc_5_axid_0_axid
        ,input [31:0]	int_desc_5_axid_1_axid
        ,input [31:0]	int_desc_5_axid_2_axid
        ,input [31:0]	int_desc_5_axid_3_axid
        ,input [31:0]	int_desc_5_axuser_0_axuser
        ,input [31:0]	int_desc_5_axuser_1_axuser
        ,input [31:0]	int_desc_5_axuser_2_axuser
        ,input [31:0]	int_desc_5_axuser_3_axuser
        ,input [31:0]	int_desc_5_axuser_4_axuser
        ,input [31:0]	int_desc_5_axuser_5_axuser
        ,input [31:0]	int_desc_5_axuser_6_axuser
        ,input [31:0]	int_desc_5_axuser_7_axuser
        ,input [31:0]	int_desc_5_axuser_8_axuser
        ,input [31:0]	int_desc_5_axuser_9_axuser
        ,input [31:0]	int_desc_5_axuser_10_axuser
        ,input [31:0]	int_desc_5_axuser_11_axuser
        ,input [31:0]	int_desc_5_axuser_12_axuser
        ,input [31:0]	int_desc_5_axuser_13_axuser
        ,input [31:0]	int_desc_5_axuser_14_axuser
        ,input [31:0]	int_desc_5_axuser_15_axuser
        ,input [31:0]	int_desc_5_size_txn_size
        ,input [2:0]	int_desc_5_axsize_axsize
        ,input [31:0]	int_desc_5_axaddr_0_addr
        ,input [31:0]	int_desc_5_axaddr_1_addr
        ,input [31:0]	int_desc_5_axaddr_2_addr
        ,input [31:0]	int_desc_5_axaddr_3_addr
        ,input [31:0]	int_desc_5_data_offset_addr
        ,input [31:0]	int_desc_5_wuser_0_wuser
        ,input [31:0]	int_desc_5_wuser_1_wuser
        ,input [31:0]	int_desc_5_wuser_2_wuser
        ,input [31:0]	int_desc_5_wuser_3_wuser
        ,input [31:0]	int_desc_5_wuser_4_wuser
        ,input [31:0]	int_desc_5_wuser_5_wuser
        ,input [31:0]	int_desc_5_wuser_6_wuser
        ,input [31:0]	int_desc_5_wuser_7_wuser
        ,input [31:0]	int_desc_5_wuser_8_wuser
        ,input [31:0]	int_desc_5_wuser_9_wuser
        ,input [31:0]	int_desc_5_wuser_10_wuser
        ,input [31:0]	int_desc_5_wuser_11_wuser
        ,input [31:0]	int_desc_5_wuser_12_wuser
        ,input [31:0]	int_desc_5_wuser_13_wuser
        ,input [31:0]	int_desc_5_wuser_14_wuser
        ,input [31:0]	int_desc_5_wuser_15_wuser
        ,input [0:0]	int_desc_6_txn_type_wr_strb
        ,input [0:0]	int_desc_6_txn_type_wr_rd
        ,input [3:0]	int_desc_6_attr_axregion
        ,input [3:0]	int_desc_6_attr_axqos
        ,input [2:0]	int_desc_6_attr_axprot
        ,input [3:0]	int_desc_6_attr_axcache
        ,input [1:0]	int_desc_6_attr_axlock
        ,input [1:0]	int_desc_6_attr_axburst
        ,input [31:0]	int_desc_6_axid_0_axid
        ,input [31:0]	int_desc_6_axid_1_axid
        ,input [31:0]	int_desc_6_axid_2_axid
        ,input [31:0]	int_desc_6_axid_3_axid
        ,input [31:0]	int_desc_6_axuser_0_axuser
        ,input [31:0]	int_desc_6_axuser_1_axuser
        ,input [31:0]	int_desc_6_axuser_2_axuser
        ,input [31:0]	int_desc_6_axuser_3_axuser
        ,input [31:0]	int_desc_6_axuser_4_axuser
        ,input [31:0]	int_desc_6_axuser_5_axuser
        ,input [31:0]	int_desc_6_axuser_6_axuser
        ,input [31:0]	int_desc_6_axuser_7_axuser
        ,input [31:0]	int_desc_6_axuser_8_axuser
        ,input [31:0]	int_desc_6_axuser_9_axuser
        ,input [31:0]	int_desc_6_axuser_10_axuser
        ,input [31:0]	int_desc_6_axuser_11_axuser
        ,input [31:0]	int_desc_6_axuser_12_axuser
        ,input [31:0]	int_desc_6_axuser_13_axuser
        ,input [31:0]	int_desc_6_axuser_14_axuser
        ,input [31:0]	int_desc_6_axuser_15_axuser
        ,input [31:0]	int_desc_6_size_txn_size
        ,input [2:0]	int_desc_6_axsize_axsize
        ,input [31:0]	int_desc_6_axaddr_0_addr
        ,input [31:0]	int_desc_6_axaddr_1_addr
        ,input [31:0]	int_desc_6_axaddr_2_addr
        ,input [31:0]	int_desc_6_axaddr_3_addr
        ,input [31:0]	int_desc_6_data_offset_addr
        ,input [31:0]	int_desc_6_wuser_0_wuser
        ,input [31:0]	int_desc_6_wuser_1_wuser
        ,input [31:0]	int_desc_6_wuser_2_wuser
        ,input [31:0]	int_desc_6_wuser_3_wuser
        ,input [31:0]	int_desc_6_wuser_4_wuser
        ,input [31:0]	int_desc_6_wuser_5_wuser
        ,input [31:0]	int_desc_6_wuser_6_wuser
        ,input [31:0]	int_desc_6_wuser_7_wuser
        ,input [31:0]	int_desc_6_wuser_8_wuser
        ,input [31:0]	int_desc_6_wuser_9_wuser
        ,input [31:0]	int_desc_6_wuser_10_wuser
        ,input [31:0]	int_desc_6_wuser_11_wuser
        ,input [31:0]	int_desc_6_wuser_12_wuser
        ,input [31:0]	int_desc_6_wuser_13_wuser
        ,input [31:0]	int_desc_6_wuser_14_wuser
        ,input [31:0]	int_desc_6_wuser_15_wuser
        ,input [0:0]	int_desc_7_txn_type_wr_strb
        ,input [0:0]	int_desc_7_txn_type_wr_rd
        ,input [3:0]	int_desc_7_attr_axregion
        ,input [3:0]	int_desc_7_attr_axqos
        ,input [2:0]	int_desc_7_attr_axprot
        ,input [3:0]	int_desc_7_attr_axcache
        ,input [1:0]	int_desc_7_attr_axlock
        ,input [1:0]	int_desc_7_attr_axburst
        ,input [31:0]	int_desc_7_axid_0_axid
        ,input [31:0]	int_desc_7_axid_1_axid
        ,input [31:0]	int_desc_7_axid_2_axid
        ,input [31:0]	int_desc_7_axid_3_axid
        ,input [31:0]	int_desc_7_axuser_0_axuser
        ,input [31:0]	int_desc_7_axuser_1_axuser
        ,input [31:0]	int_desc_7_axuser_2_axuser
        ,input [31:0]	int_desc_7_axuser_3_axuser
        ,input [31:0]	int_desc_7_axuser_4_axuser
        ,input [31:0]	int_desc_7_axuser_5_axuser
        ,input [31:0]	int_desc_7_axuser_6_axuser
        ,input [31:0]	int_desc_7_axuser_7_axuser
        ,input [31:0]	int_desc_7_axuser_8_axuser
        ,input [31:0]	int_desc_7_axuser_9_axuser
        ,input [31:0]	int_desc_7_axuser_10_axuser
        ,input [31:0]	int_desc_7_axuser_11_axuser
        ,input [31:0]	int_desc_7_axuser_12_axuser
        ,input [31:0]	int_desc_7_axuser_13_axuser
        ,input [31:0]	int_desc_7_axuser_14_axuser
        ,input [31:0]	int_desc_7_axuser_15_axuser
        ,input [31:0]	int_desc_7_size_txn_size
        ,input [2:0]	int_desc_7_axsize_axsize
        ,input [31:0]	int_desc_7_axaddr_0_addr
        ,input [31:0]	int_desc_7_axaddr_1_addr
        ,input [31:0]	int_desc_7_axaddr_2_addr
        ,input [31:0]	int_desc_7_axaddr_3_addr
        ,input [31:0]	int_desc_7_data_offset_addr
        ,input [31:0]	int_desc_7_wuser_0_wuser
        ,input [31:0]	int_desc_7_wuser_1_wuser
        ,input [31:0]	int_desc_7_wuser_2_wuser
        ,input [31:0]	int_desc_7_wuser_3_wuser
        ,input [31:0]	int_desc_7_wuser_4_wuser
        ,input [31:0]	int_desc_7_wuser_5_wuser
        ,input [31:0]	int_desc_7_wuser_6_wuser
        ,input [31:0]	int_desc_7_wuser_7_wuser
        ,input [31:0]	int_desc_7_wuser_8_wuser
        ,input [31:0]	int_desc_7_wuser_9_wuser
        ,input [31:0]	int_desc_7_wuser_10_wuser
        ,input [31:0]	int_desc_7_wuser_11_wuser
        ,input [31:0]	int_desc_7_wuser_12_wuser
        ,input [31:0]	int_desc_7_wuser_13_wuser
        ,input [31:0]	int_desc_7_wuser_14_wuser
        ,input [31:0]	int_desc_7_wuser_15_wuser
        ,input [0:0]	int_desc_8_txn_type_wr_strb
        ,input [0:0]	int_desc_8_txn_type_wr_rd
        ,input [3:0]	int_desc_8_attr_axregion
        ,input [3:0]	int_desc_8_attr_axqos
        ,input [2:0]	int_desc_8_attr_axprot
        ,input [3:0]	int_desc_8_attr_axcache
        ,input [1:0]	int_desc_8_attr_axlock
        ,input [1:0]	int_desc_8_attr_axburst
        ,input [31:0]	int_desc_8_axid_0_axid
        ,input [31:0]	int_desc_8_axid_1_axid
        ,input [31:0]	int_desc_8_axid_2_axid
        ,input [31:0]	int_desc_8_axid_3_axid
        ,input [31:0]	int_desc_8_axuser_0_axuser
        ,input [31:0]	int_desc_8_axuser_1_axuser
        ,input [31:0]	int_desc_8_axuser_2_axuser
        ,input [31:0]	int_desc_8_axuser_3_axuser
        ,input [31:0]	int_desc_8_axuser_4_axuser
        ,input [31:0]	int_desc_8_axuser_5_axuser
        ,input [31:0]	int_desc_8_axuser_6_axuser
        ,input [31:0]	int_desc_8_axuser_7_axuser
        ,input [31:0]	int_desc_8_axuser_8_axuser
        ,input [31:0]	int_desc_8_axuser_9_axuser
        ,input [31:0]	int_desc_8_axuser_10_axuser
        ,input [31:0]	int_desc_8_axuser_11_axuser
        ,input [31:0]	int_desc_8_axuser_12_axuser
        ,input [31:0]	int_desc_8_axuser_13_axuser
        ,input [31:0]	int_desc_8_axuser_14_axuser
        ,input [31:0]	int_desc_8_axuser_15_axuser
        ,input [31:0]	int_desc_8_size_txn_size
        ,input [2:0]	int_desc_8_axsize_axsize
        ,input [31:0]	int_desc_8_axaddr_0_addr
        ,input [31:0]	int_desc_8_axaddr_1_addr
        ,input [31:0]	int_desc_8_axaddr_2_addr
        ,input [31:0]	int_desc_8_axaddr_3_addr
        ,input [31:0]	int_desc_8_data_offset_addr
        ,input [31:0]	int_desc_8_wuser_0_wuser
        ,input [31:0]	int_desc_8_wuser_1_wuser
        ,input [31:0]	int_desc_8_wuser_2_wuser
        ,input [31:0]	int_desc_8_wuser_3_wuser
        ,input [31:0]	int_desc_8_wuser_4_wuser
        ,input [31:0]	int_desc_8_wuser_5_wuser
        ,input [31:0]	int_desc_8_wuser_6_wuser
        ,input [31:0]	int_desc_8_wuser_7_wuser
        ,input [31:0]	int_desc_8_wuser_8_wuser
        ,input [31:0]	int_desc_8_wuser_9_wuser
        ,input [31:0]	int_desc_8_wuser_10_wuser
        ,input [31:0]	int_desc_8_wuser_11_wuser
        ,input [31:0]	int_desc_8_wuser_12_wuser
        ,input [31:0]	int_desc_8_wuser_13_wuser
        ,input [31:0]	int_desc_8_wuser_14_wuser
        ,input [31:0]	int_desc_8_wuser_15_wuser
        ,input [0:0]	int_desc_9_txn_type_wr_strb
        ,input [0:0]	int_desc_9_txn_type_wr_rd
        ,input [3:0]	int_desc_9_attr_axregion
        ,input [3:0]	int_desc_9_attr_axqos
        ,input [2:0]	int_desc_9_attr_axprot
        ,input [3:0]	int_desc_9_attr_axcache
        ,input [1:0]	int_desc_9_attr_axlock
        ,input [1:0]	int_desc_9_attr_axburst
        ,input [31:0]	int_desc_9_axid_0_axid
        ,input [31:0]	int_desc_9_axid_1_axid
        ,input [31:0]	int_desc_9_axid_2_axid
        ,input [31:0]	int_desc_9_axid_3_axid
        ,input [31:0]	int_desc_9_axuser_0_axuser
        ,input [31:0]	int_desc_9_axuser_1_axuser
        ,input [31:0]	int_desc_9_axuser_2_axuser
        ,input [31:0]	int_desc_9_axuser_3_axuser
        ,input [31:0]	int_desc_9_axuser_4_axuser
        ,input [31:0]	int_desc_9_axuser_5_axuser
        ,input [31:0]	int_desc_9_axuser_6_axuser
        ,input [31:0]	int_desc_9_axuser_7_axuser
        ,input [31:0]	int_desc_9_axuser_8_axuser
        ,input [31:0]	int_desc_9_axuser_9_axuser
        ,input [31:0]	int_desc_9_axuser_10_axuser
        ,input [31:0]	int_desc_9_axuser_11_axuser
        ,input [31:0]	int_desc_9_axuser_12_axuser
        ,input [31:0]	int_desc_9_axuser_13_axuser
        ,input [31:0]	int_desc_9_axuser_14_axuser
        ,input [31:0]	int_desc_9_axuser_15_axuser
        ,input [31:0]	int_desc_9_size_txn_size
        ,input [2:0]	int_desc_9_axsize_axsize
        ,input [31:0]	int_desc_9_axaddr_0_addr
        ,input [31:0]	int_desc_9_axaddr_1_addr
        ,input [31:0]	int_desc_9_axaddr_2_addr
        ,input [31:0]	int_desc_9_axaddr_3_addr
        ,input [31:0]	int_desc_9_data_offset_addr
        ,input [31:0]	int_desc_9_wuser_0_wuser
        ,input [31:0]	int_desc_9_wuser_1_wuser
        ,input [31:0]	int_desc_9_wuser_2_wuser
        ,input [31:0]	int_desc_9_wuser_3_wuser
        ,input [31:0]	int_desc_9_wuser_4_wuser
        ,input [31:0]	int_desc_9_wuser_5_wuser
        ,input [31:0]	int_desc_9_wuser_6_wuser
        ,input [31:0]	int_desc_9_wuser_7_wuser
        ,input [31:0]	int_desc_9_wuser_8_wuser
        ,input [31:0]	int_desc_9_wuser_9_wuser
        ,input [31:0]	int_desc_9_wuser_10_wuser
        ,input [31:0]	int_desc_9_wuser_11_wuser
        ,input [31:0]	int_desc_9_wuser_12_wuser
        ,input [31:0]	int_desc_9_wuser_13_wuser
        ,input [31:0]	int_desc_9_wuser_14_wuser
        ,input [31:0]	int_desc_9_wuser_15_wuser
        ,input [0:0]	int_desc_10_txn_type_wr_strb
        ,input [0:0]	int_desc_10_txn_type_wr_rd
        ,input [3:0]	int_desc_10_attr_axregion
        ,input [3:0]	int_desc_10_attr_axqos
        ,input [2:0]	int_desc_10_attr_axprot
        ,input [3:0]	int_desc_10_attr_axcache
        ,input [1:0]	int_desc_10_attr_axlock
        ,input [1:0]	int_desc_10_attr_axburst
        ,input [31:0]	int_desc_10_axid_0_axid
        ,input [31:0]	int_desc_10_axid_1_axid
        ,input [31:0]	int_desc_10_axid_2_axid
        ,input [31:0]	int_desc_10_axid_3_axid
        ,input [31:0]	int_desc_10_axuser_0_axuser
        ,input [31:0]	int_desc_10_axuser_1_axuser
        ,input [31:0]	int_desc_10_axuser_2_axuser
        ,input [31:0]	int_desc_10_axuser_3_axuser
        ,input [31:0]	int_desc_10_axuser_4_axuser
        ,input [31:0]	int_desc_10_axuser_5_axuser
        ,input [31:0]	int_desc_10_axuser_6_axuser
        ,input [31:0]	int_desc_10_axuser_7_axuser
        ,input [31:0]	int_desc_10_axuser_8_axuser
        ,input [31:0]	int_desc_10_axuser_9_axuser
        ,input [31:0]	int_desc_10_axuser_10_axuser
        ,input [31:0]	int_desc_10_axuser_11_axuser
        ,input [31:0]	int_desc_10_axuser_12_axuser
        ,input [31:0]	int_desc_10_axuser_13_axuser
        ,input [31:0]	int_desc_10_axuser_14_axuser
        ,input [31:0]	int_desc_10_axuser_15_axuser
        ,input [31:0]	int_desc_10_size_txn_size
        ,input [2:0]	int_desc_10_axsize_axsize
        ,input [31:0]	int_desc_10_axaddr_0_addr
        ,input [31:0]	int_desc_10_axaddr_1_addr
        ,input [31:0]	int_desc_10_axaddr_2_addr
        ,input [31:0]	int_desc_10_axaddr_3_addr
        ,input [31:0]	int_desc_10_data_offset_addr
        ,input [31:0]	int_desc_10_wuser_0_wuser
        ,input [31:0]	int_desc_10_wuser_1_wuser
        ,input [31:0]	int_desc_10_wuser_2_wuser
        ,input [31:0]	int_desc_10_wuser_3_wuser
        ,input [31:0]	int_desc_10_wuser_4_wuser
        ,input [31:0]	int_desc_10_wuser_5_wuser
        ,input [31:0]	int_desc_10_wuser_6_wuser
        ,input [31:0]	int_desc_10_wuser_7_wuser
        ,input [31:0]	int_desc_10_wuser_8_wuser
        ,input [31:0]	int_desc_10_wuser_9_wuser
        ,input [31:0]	int_desc_10_wuser_10_wuser
        ,input [31:0]	int_desc_10_wuser_11_wuser
        ,input [31:0]	int_desc_10_wuser_12_wuser
        ,input [31:0]	int_desc_10_wuser_13_wuser
        ,input [31:0]	int_desc_10_wuser_14_wuser
        ,input [31:0]	int_desc_10_wuser_15_wuser
        ,input [0:0]	int_desc_11_txn_type_wr_strb
        ,input [0:0]	int_desc_11_txn_type_wr_rd
        ,input [3:0]	int_desc_11_attr_axregion
        ,input [3:0]	int_desc_11_attr_axqos
        ,input [2:0]	int_desc_11_attr_axprot
        ,input [3:0]	int_desc_11_attr_axcache
        ,input [1:0]	int_desc_11_attr_axlock
        ,input [1:0]	int_desc_11_attr_axburst
        ,input [31:0]	int_desc_11_axid_0_axid
        ,input [31:0]	int_desc_11_axid_1_axid
        ,input [31:0]	int_desc_11_axid_2_axid
        ,input [31:0]	int_desc_11_axid_3_axid
        ,input [31:0]	int_desc_11_axuser_0_axuser
        ,input [31:0]	int_desc_11_axuser_1_axuser
        ,input [31:0]	int_desc_11_axuser_2_axuser
        ,input [31:0]	int_desc_11_axuser_3_axuser
        ,input [31:0]	int_desc_11_axuser_4_axuser
        ,input [31:0]	int_desc_11_axuser_5_axuser
        ,input [31:0]	int_desc_11_axuser_6_axuser
        ,input [31:0]	int_desc_11_axuser_7_axuser
        ,input [31:0]	int_desc_11_axuser_8_axuser
        ,input [31:0]	int_desc_11_axuser_9_axuser
        ,input [31:0]	int_desc_11_axuser_10_axuser
        ,input [31:0]	int_desc_11_axuser_11_axuser
        ,input [31:0]	int_desc_11_axuser_12_axuser
        ,input [31:0]	int_desc_11_axuser_13_axuser
        ,input [31:0]	int_desc_11_axuser_14_axuser
        ,input [31:0]	int_desc_11_axuser_15_axuser
        ,input [31:0]	int_desc_11_size_txn_size
        ,input [2:0]	int_desc_11_axsize_axsize
        ,input [31:0]	int_desc_11_axaddr_0_addr
        ,input [31:0]	int_desc_11_axaddr_1_addr
        ,input [31:0]	int_desc_11_axaddr_2_addr
        ,input [31:0]	int_desc_11_axaddr_3_addr
        ,input [31:0]	int_desc_11_data_offset_addr
        ,input [31:0]	int_desc_11_wuser_0_wuser
        ,input [31:0]	int_desc_11_wuser_1_wuser
        ,input [31:0]	int_desc_11_wuser_2_wuser
        ,input [31:0]	int_desc_11_wuser_3_wuser
        ,input [31:0]	int_desc_11_wuser_4_wuser
        ,input [31:0]	int_desc_11_wuser_5_wuser
        ,input [31:0]	int_desc_11_wuser_6_wuser
        ,input [31:0]	int_desc_11_wuser_7_wuser
        ,input [31:0]	int_desc_11_wuser_8_wuser
        ,input [31:0]	int_desc_11_wuser_9_wuser
        ,input [31:0]	int_desc_11_wuser_10_wuser
        ,input [31:0]	int_desc_11_wuser_11_wuser
        ,input [31:0]	int_desc_11_wuser_12_wuser
        ,input [31:0]	int_desc_11_wuser_13_wuser
        ,input [31:0]	int_desc_11_wuser_14_wuser
        ,input [31:0]	int_desc_11_wuser_15_wuser
        ,input [0:0]	int_desc_12_txn_type_wr_strb
        ,input [0:0]	int_desc_12_txn_type_wr_rd
        ,input [3:0]	int_desc_12_attr_axregion
        ,input [3:0]	int_desc_12_attr_axqos
        ,input [2:0]	int_desc_12_attr_axprot
        ,input [3:0]	int_desc_12_attr_axcache
        ,input [1:0]	int_desc_12_attr_axlock
        ,input [1:0]	int_desc_12_attr_axburst
        ,input [31:0]	int_desc_12_axid_0_axid
        ,input [31:0]	int_desc_12_axid_1_axid
        ,input [31:0]	int_desc_12_axid_2_axid
        ,input [31:0]	int_desc_12_axid_3_axid
        ,input [31:0]	int_desc_12_axuser_0_axuser
        ,input [31:0]	int_desc_12_axuser_1_axuser
        ,input [31:0]	int_desc_12_axuser_2_axuser
        ,input [31:0]	int_desc_12_axuser_3_axuser
        ,input [31:0]	int_desc_12_axuser_4_axuser
        ,input [31:0]	int_desc_12_axuser_5_axuser
        ,input [31:0]	int_desc_12_axuser_6_axuser
        ,input [31:0]	int_desc_12_axuser_7_axuser
        ,input [31:0]	int_desc_12_axuser_8_axuser
        ,input [31:0]	int_desc_12_axuser_9_axuser
        ,input [31:0]	int_desc_12_axuser_10_axuser
        ,input [31:0]	int_desc_12_axuser_11_axuser
        ,input [31:0]	int_desc_12_axuser_12_axuser
        ,input [31:0]	int_desc_12_axuser_13_axuser
        ,input [31:0]	int_desc_12_axuser_14_axuser
        ,input [31:0]	int_desc_12_axuser_15_axuser
        ,input [31:0]	int_desc_12_size_txn_size
        ,input [2:0]	int_desc_12_axsize_axsize
        ,input [31:0]	int_desc_12_axaddr_0_addr
        ,input [31:0]	int_desc_12_axaddr_1_addr
        ,input [31:0]	int_desc_12_axaddr_2_addr
        ,input [31:0]	int_desc_12_axaddr_3_addr
        ,input [31:0]	int_desc_12_data_offset_addr
        ,input [31:0]	int_desc_12_wuser_0_wuser
        ,input [31:0]	int_desc_12_wuser_1_wuser
        ,input [31:0]	int_desc_12_wuser_2_wuser
        ,input [31:0]	int_desc_12_wuser_3_wuser
        ,input [31:0]	int_desc_12_wuser_4_wuser
        ,input [31:0]	int_desc_12_wuser_5_wuser
        ,input [31:0]	int_desc_12_wuser_6_wuser
        ,input [31:0]	int_desc_12_wuser_7_wuser
        ,input [31:0]	int_desc_12_wuser_8_wuser
        ,input [31:0]	int_desc_12_wuser_9_wuser
        ,input [31:0]	int_desc_12_wuser_10_wuser
        ,input [31:0]	int_desc_12_wuser_11_wuser
        ,input [31:0]	int_desc_12_wuser_12_wuser
        ,input [31:0]	int_desc_12_wuser_13_wuser
        ,input [31:0]	int_desc_12_wuser_14_wuser
        ,input [31:0]	int_desc_12_wuser_15_wuser
        ,input [0:0]	int_desc_13_txn_type_wr_strb
        ,input [0:0]	int_desc_13_txn_type_wr_rd
        ,input [3:0]	int_desc_13_attr_axregion
        ,input [3:0]	int_desc_13_attr_axqos
        ,input [2:0]	int_desc_13_attr_axprot
        ,input [3:0]	int_desc_13_attr_axcache
        ,input [1:0]	int_desc_13_attr_axlock
        ,input [1:0]	int_desc_13_attr_axburst
        ,input [31:0]	int_desc_13_axid_0_axid
        ,input [31:0]	int_desc_13_axid_1_axid
        ,input [31:0]	int_desc_13_axid_2_axid
        ,input [31:0]	int_desc_13_axid_3_axid
        ,input [31:0]	int_desc_13_axuser_0_axuser
        ,input [31:0]	int_desc_13_axuser_1_axuser
        ,input [31:0]	int_desc_13_axuser_2_axuser
        ,input [31:0]	int_desc_13_axuser_3_axuser
        ,input [31:0]	int_desc_13_axuser_4_axuser
        ,input [31:0]	int_desc_13_axuser_5_axuser
        ,input [31:0]	int_desc_13_axuser_6_axuser
        ,input [31:0]	int_desc_13_axuser_7_axuser
        ,input [31:0]	int_desc_13_axuser_8_axuser
        ,input [31:0]	int_desc_13_axuser_9_axuser
        ,input [31:0]	int_desc_13_axuser_10_axuser
        ,input [31:0]	int_desc_13_axuser_11_axuser
        ,input [31:0]	int_desc_13_axuser_12_axuser
        ,input [31:0]	int_desc_13_axuser_13_axuser
        ,input [31:0]	int_desc_13_axuser_14_axuser
        ,input [31:0]	int_desc_13_axuser_15_axuser
        ,input [31:0]	int_desc_13_size_txn_size
        ,input [2:0]	int_desc_13_axsize_axsize
        ,input [31:0]	int_desc_13_axaddr_0_addr
        ,input [31:0]	int_desc_13_axaddr_1_addr
        ,input [31:0]	int_desc_13_axaddr_2_addr
        ,input [31:0]	int_desc_13_axaddr_3_addr
        ,input [31:0]	int_desc_13_data_offset_addr
        ,input [31:0]	int_desc_13_wuser_0_wuser
        ,input [31:0]	int_desc_13_wuser_1_wuser
        ,input [31:0]	int_desc_13_wuser_2_wuser
        ,input [31:0]	int_desc_13_wuser_3_wuser
        ,input [31:0]	int_desc_13_wuser_4_wuser
        ,input [31:0]	int_desc_13_wuser_5_wuser
        ,input [31:0]	int_desc_13_wuser_6_wuser
        ,input [31:0]	int_desc_13_wuser_7_wuser
        ,input [31:0]	int_desc_13_wuser_8_wuser
        ,input [31:0]	int_desc_13_wuser_9_wuser
        ,input [31:0]	int_desc_13_wuser_10_wuser
        ,input [31:0]	int_desc_13_wuser_11_wuser
        ,input [31:0]	int_desc_13_wuser_12_wuser
        ,input [31:0]	int_desc_13_wuser_13_wuser
        ,input [31:0]	int_desc_13_wuser_14_wuser
        ,input [31:0]	int_desc_13_wuser_15_wuser
        ,input [0:0]	int_desc_14_txn_type_wr_strb
        ,input [0:0]	int_desc_14_txn_type_wr_rd
        ,input [3:0]	int_desc_14_attr_axregion
        ,input [3:0]	int_desc_14_attr_axqos
        ,input [2:0]	int_desc_14_attr_axprot
        ,input [3:0]	int_desc_14_attr_axcache
        ,input [1:0]	int_desc_14_attr_axlock
        ,input [1:0]	int_desc_14_attr_axburst
        ,input [31:0]	int_desc_14_axid_0_axid
        ,input [31:0]	int_desc_14_axid_1_axid
        ,input [31:0]	int_desc_14_axid_2_axid
        ,input [31:0]	int_desc_14_axid_3_axid
        ,input [31:0]	int_desc_14_axuser_0_axuser
        ,input [31:0]	int_desc_14_axuser_1_axuser
        ,input [31:0]	int_desc_14_axuser_2_axuser
        ,input [31:0]	int_desc_14_axuser_3_axuser
        ,input [31:0]	int_desc_14_axuser_4_axuser
        ,input [31:0]	int_desc_14_axuser_5_axuser
        ,input [31:0]	int_desc_14_axuser_6_axuser
        ,input [31:0]	int_desc_14_axuser_7_axuser
        ,input [31:0]	int_desc_14_axuser_8_axuser
        ,input [31:0]	int_desc_14_axuser_9_axuser
        ,input [31:0]	int_desc_14_axuser_10_axuser
        ,input [31:0]	int_desc_14_axuser_11_axuser
        ,input [31:0]	int_desc_14_axuser_12_axuser
        ,input [31:0]	int_desc_14_axuser_13_axuser
        ,input [31:0]	int_desc_14_axuser_14_axuser
        ,input [31:0]	int_desc_14_axuser_15_axuser
        ,input [31:0]	int_desc_14_size_txn_size
        ,input [2:0]	int_desc_14_axsize_axsize
        ,input [31:0]	int_desc_14_axaddr_0_addr
        ,input [31:0]	int_desc_14_axaddr_1_addr
        ,input [31:0]	int_desc_14_axaddr_2_addr
        ,input [31:0]	int_desc_14_axaddr_3_addr
        ,input [31:0]	int_desc_14_data_offset_addr
        ,input [31:0]	int_desc_14_wuser_0_wuser
        ,input [31:0]	int_desc_14_wuser_1_wuser
        ,input [31:0]	int_desc_14_wuser_2_wuser
        ,input [31:0]	int_desc_14_wuser_3_wuser
        ,input [31:0]	int_desc_14_wuser_4_wuser
        ,input [31:0]	int_desc_14_wuser_5_wuser
        ,input [31:0]	int_desc_14_wuser_6_wuser
        ,input [31:0]	int_desc_14_wuser_7_wuser
        ,input [31:0]	int_desc_14_wuser_8_wuser
        ,input [31:0]	int_desc_14_wuser_9_wuser
        ,input [31:0]	int_desc_14_wuser_10_wuser
        ,input [31:0]	int_desc_14_wuser_11_wuser
        ,input [31:0]	int_desc_14_wuser_12_wuser
        ,input [31:0]	int_desc_14_wuser_13_wuser
        ,input [31:0]	int_desc_14_wuser_14_wuser
        ,input [31:0]	int_desc_14_wuser_15_wuser
        ,input [0:0]	int_desc_15_txn_type_wr_strb
        ,input [0:0]	int_desc_15_txn_type_wr_rd
        ,input [3:0]	int_desc_15_attr_axregion
        ,input [3:0]	int_desc_15_attr_axqos
        ,input [2:0]	int_desc_15_attr_axprot
        ,input [3:0]	int_desc_15_attr_axcache
        ,input [1:0]	int_desc_15_attr_axlock
        ,input [1:0]	int_desc_15_attr_axburst
        ,input [31:0]	int_desc_15_axid_0_axid
        ,input [31:0]	int_desc_15_axid_1_axid
        ,input [31:0]	int_desc_15_axid_2_axid
        ,input [31:0]	int_desc_15_axid_3_axid
        ,input [31:0]	int_desc_15_axuser_0_axuser
        ,input [31:0]	int_desc_15_axuser_1_axuser
        ,input [31:0]	int_desc_15_axuser_2_axuser
        ,input [31:0]	int_desc_15_axuser_3_axuser
        ,input [31:0]	int_desc_15_axuser_4_axuser
        ,input [31:0]	int_desc_15_axuser_5_axuser
        ,input [31:0]	int_desc_15_axuser_6_axuser
        ,input [31:0]	int_desc_15_axuser_7_axuser
        ,input [31:0]	int_desc_15_axuser_8_axuser
        ,input [31:0]	int_desc_15_axuser_9_axuser
        ,input [31:0]	int_desc_15_axuser_10_axuser
        ,input [31:0]	int_desc_15_axuser_11_axuser
        ,input [31:0]	int_desc_15_axuser_12_axuser
        ,input [31:0]	int_desc_15_axuser_13_axuser
        ,input [31:0]	int_desc_15_axuser_14_axuser
        ,input [31:0]	int_desc_15_axuser_15_axuser
        ,input [31:0]	int_desc_15_size_txn_size
        ,input [2:0]	int_desc_15_axsize_axsize
        ,input [31:0]	int_desc_15_axaddr_0_addr
        ,input [31:0]	int_desc_15_axaddr_1_addr
        ,input [31:0]	int_desc_15_axaddr_2_addr
        ,input [31:0]	int_desc_15_axaddr_3_addr
        ,input [31:0]	int_desc_15_data_offset_addr
        ,input [31:0]	int_desc_15_wuser_0_wuser
        ,input [31:0]	int_desc_15_wuser_1_wuser
        ,input [31:0]	int_desc_15_wuser_2_wuser
        ,input [31:0]	int_desc_15_wuser_3_wuser
        ,input [31:0]	int_desc_15_wuser_4_wuser
        ,input [31:0]	int_desc_15_wuser_5_wuser
        ,input [31:0]	int_desc_15_wuser_6_wuser
        ,input [31:0]	int_desc_15_wuser_7_wuser
        ,input [31:0]	int_desc_15_wuser_8_wuser
        ,input [31:0]	int_desc_15_wuser_9_wuser
        ,input [31:0]	int_desc_15_wuser_10_wuser
        ,input [31:0]	int_desc_15_wuser_11_wuser
        ,input [31:0]	int_desc_15_wuser_12_wuser
        ,input [31:0]	int_desc_15_wuser_13_wuser
        ,input [31:0]	int_desc_15_wuser_14_wuser
        ,input [31:0]	int_desc_15_wuser_15_wuser

        ,input  [31:0]	int_desc_0_data_host_addr_0_addr
        ,input  [31:0]	int_desc_0_data_host_addr_1_addr
        ,input  [31:0]	int_desc_0_data_host_addr_2_addr
        ,input  [31:0]	int_desc_0_data_host_addr_3_addr
        ,input  [31:0]	int_desc_0_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_0_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_0_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_0_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_1_data_host_addr_0_addr
        ,input  [31:0]	int_desc_1_data_host_addr_1_addr
        ,input  [31:0]	int_desc_1_data_host_addr_2_addr
        ,input  [31:0]	int_desc_1_data_host_addr_3_addr
        ,input  [31:0]	int_desc_1_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_1_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_1_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_1_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_2_data_host_addr_0_addr
        ,input  [31:0]	int_desc_2_data_host_addr_1_addr
        ,input  [31:0]	int_desc_2_data_host_addr_2_addr
        ,input  [31:0]	int_desc_2_data_host_addr_3_addr
        ,input  [31:0]	int_desc_2_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_2_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_2_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_2_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_3_data_host_addr_0_addr
        ,input  [31:0]	int_desc_3_data_host_addr_1_addr
        ,input  [31:0]	int_desc_3_data_host_addr_2_addr
        ,input  [31:0]	int_desc_3_data_host_addr_3_addr
        ,input  [31:0]	int_desc_3_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_3_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_3_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_3_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_4_data_host_addr_0_addr
        ,input  [31:0]	int_desc_4_data_host_addr_1_addr
        ,input  [31:0]	int_desc_4_data_host_addr_2_addr
        ,input  [31:0]	int_desc_4_data_host_addr_3_addr
        ,input  [31:0]	int_desc_4_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_4_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_4_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_4_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_5_data_host_addr_0_addr
        ,input  [31:0]	int_desc_5_data_host_addr_1_addr
        ,input  [31:0]	int_desc_5_data_host_addr_2_addr
        ,input  [31:0]	int_desc_5_data_host_addr_3_addr
        ,input  [31:0]	int_desc_5_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_5_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_5_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_5_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_6_data_host_addr_0_addr
        ,input  [31:0]	int_desc_6_data_host_addr_1_addr
        ,input  [31:0]	int_desc_6_data_host_addr_2_addr
        ,input  [31:0]	int_desc_6_data_host_addr_3_addr
        ,input  [31:0]	int_desc_6_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_6_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_6_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_6_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_7_data_host_addr_0_addr
        ,input  [31:0]	int_desc_7_data_host_addr_1_addr
        ,input  [31:0]	int_desc_7_data_host_addr_2_addr
        ,input  [31:0]	int_desc_7_data_host_addr_3_addr
        ,input  [31:0]	int_desc_7_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_7_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_7_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_7_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_8_data_host_addr_0_addr
        ,input  [31:0]	int_desc_8_data_host_addr_1_addr
        ,input  [31:0]	int_desc_8_data_host_addr_2_addr
        ,input  [31:0]	int_desc_8_data_host_addr_3_addr
        ,input  [31:0]	int_desc_8_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_8_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_8_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_8_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_9_data_host_addr_0_addr
        ,input  [31:0]	int_desc_9_data_host_addr_1_addr
        ,input  [31:0]	int_desc_9_data_host_addr_2_addr
        ,input  [31:0]	int_desc_9_data_host_addr_3_addr
        ,input  [31:0]	int_desc_9_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_9_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_9_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_9_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_10_data_host_addr_0_addr
        ,input  [31:0]	int_desc_10_data_host_addr_1_addr
        ,input  [31:0]	int_desc_10_data_host_addr_2_addr
        ,input  [31:0]	int_desc_10_data_host_addr_3_addr
        ,input  [31:0]	int_desc_10_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_10_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_10_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_10_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_11_data_host_addr_0_addr
        ,input  [31:0]	int_desc_11_data_host_addr_1_addr
        ,input  [31:0]	int_desc_11_data_host_addr_2_addr
        ,input  [31:0]	int_desc_11_data_host_addr_3_addr
        ,input  [31:0]	int_desc_11_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_11_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_11_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_11_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_12_data_host_addr_0_addr
        ,input  [31:0]	int_desc_12_data_host_addr_1_addr
        ,input  [31:0]	int_desc_12_data_host_addr_2_addr
        ,input  [31:0]	int_desc_12_data_host_addr_3_addr
        ,input  [31:0]	int_desc_12_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_12_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_12_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_12_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_13_data_host_addr_0_addr
        ,input  [31:0]	int_desc_13_data_host_addr_1_addr
        ,input  [31:0]	int_desc_13_data_host_addr_2_addr
        ,input  [31:0]	int_desc_13_data_host_addr_3_addr
        ,input  [31:0]	int_desc_13_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_13_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_13_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_13_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_14_data_host_addr_0_addr
        ,input  [31:0]	int_desc_14_data_host_addr_1_addr
        ,input  [31:0]	int_desc_14_data_host_addr_2_addr
        ,input  [31:0]	int_desc_14_data_host_addr_3_addr
        ,input  [31:0]	int_desc_14_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_14_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_14_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_14_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_15_data_host_addr_0_addr
        ,input  [31:0]	int_desc_15_data_host_addr_1_addr
        ,input  [31:0]	int_desc_15_data_host_addr_2_addr
        ,input  [31:0]	int_desc_15_data_host_addr_3_addr
        ,input  [31:0]	int_desc_15_wstrb_host_addr_0_addr
        ,input  [31:0]	int_desc_15_wstrb_host_addr_1_addr
        ,input  [31:0]	int_desc_15_wstrb_host_addr_2_addr
        ,input  [31:0]	int_desc_15_wstrb_host_addr_3_addr
        ,input  [31:0]	int_desc_0_xuser_0_xuser
        ,input  [31:0]	int_desc_0_xuser_1_xuser
        ,input  [31:0]	int_desc_0_xuser_2_xuser
        ,input  [31:0]	int_desc_0_xuser_3_xuser
        ,input  [31:0]	int_desc_0_xuser_4_xuser
        ,input  [31:0]	int_desc_0_xuser_5_xuser
        ,input  [31:0]	int_desc_0_xuser_6_xuser
        ,input  [31:0]	int_desc_0_xuser_7_xuser
        ,input  [31:0]	int_desc_0_xuser_8_xuser
        ,input  [31:0]	int_desc_0_xuser_9_xuser
        ,input  [31:0]	int_desc_0_xuser_10_xuser
        ,input  [31:0]	int_desc_0_xuser_11_xuser
        ,input  [31:0]	int_desc_0_xuser_12_xuser
        ,input  [31:0]	int_desc_0_xuser_13_xuser
        ,input  [31:0]	int_desc_0_xuser_14_xuser
        ,input  [31:0]	int_desc_0_xuser_15_xuser
        ,input  [31:0]	int_desc_1_xuser_0_xuser
        ,input  [31:0]	int_desc_1_xuser_1_xuser
        ,input  [31:0]	int_desc_1_xuser_2_xuser
        ,input  [31:0]	int_desc_1_xuser_3_xuser
        ,input  [31:0]	int_desc_1_xuser_4_xuser
        ,input  [31:0]	int_desc_1_xuser_5_xuser
        ,input  [31:0]	int_desc_1_xuser_6_xuser
        ,input  [31:0]	int_desc_1_xuser_7_xuser
        ,input  [31:0]	int_desc_1_xuser_8_xuser
        ,input  [31:0]	int_desc_1_xuser_9_xuser
        ,input  [31:0]	int_desc_1_xuser_10_xuser
        ,input  [31:0]	int_desc_1_xuser_11_xuser
        ,input  [31:0]	int_desc_1_xuser_12_xuser
        ,input  [31:0]	int_desc_1_xuser_13_xuser
        ,input  [31:0]	int_desc_1_xuser_14_xuser
        ,input  [31:0]	int_desc_1_xuser_15_xuser
        ,input  [31:0]	int_desc_2_xuser_0_xuser
        ,input  [31:0]	int_desc_2_xuser_1_xuser
        ,input  [31:0]	int_desc_2_xuser_2_xuser
        ,input  [31:0]	int_desc_2_xuser_3_xuser
        ,input  [31:0]	int_desc_2_xuser_4_xuser
        ,input  [31:0]	int_desc_2_xuser_5_xuser
        ,input  [31:0]	int_desc_2_xuser_6_xuser
        ,input  [31:0]	int_desc_2_xuser_7_xuser
        ,input  [31:0]	int_desc_2_xuser_8_xuser
        ,input  [31:0]	int_desc_2_xuser_9_xuser
        ,input  [31:0]	int_desc_2_xuser_10_xuser
        ,input  [31:0]	int_desc_2_xuser_11_xuser
        ,input  [31:0]	int_desc_2_xuser_12_xuser
        ,input  [31:0]	int_desc_2_xuser_13_xuser
        ,input  [31:0]	int_desc_2_xuser_14_xuser
        ,input  [31:0]	int_desc_2_xuser_15_xuser
        ,input  [31:0]	int_desc_3_xuser_0_xuser
        ,input  [31:0]	int_desc_3_xuser_1_xuser
        ,input  [31:0]	int_desc_3_xuser_2_xuser
        ,input  [31:0]	int_desc_3_xuser_3_xuser
        ,input  [31:0]	int_desc_3_xuser_4_xuser
        ,input  [31:0]	int_desc_3_xuser_5_xuser
        ,input  [31:0]	int_desc_3_xuser_6_xuser
        ,input  [31:0]	int_desc_3_xuser_7_xuser
        ,input  [31:0]	int_desc_3_xuser_8_xuser
        ,input  [31:0]	int_desc_3_xuser_9_xuser
        ,input  [31:0]	int_desc_3_xuser_10_xuser
        ,input  [31:0]	int_desc_3_xuser_11_xuser
        ,input  [31:0]	int_desc_3_xuser_12_xuser
        ,input  [31:0]	int_desc_3_xuser_13_xuser
        ,input  [31:0]	int_desc_3_xuser_14_xuser
        ,input  [31:0]	int_desc_3_xuser_15_xuser
        ,input  [31:0]	int_desc_4_xuser_0_xuser
        ,input  [31:0]	int_desc_4_xuser_1_xuser
        ,input  [31:0]	int_desc_4_xuser_2_xuser
        ,input  [31:0]	int_desc_4_xuser_3_xuser
        ,input  [31:0]	int_desc_4_xuser_4_xuser
        ,input  [31:0]	int_desc_4_xuser_5_xuser
        ,input  [31:0]	int_desc_4_xuser_6_xuser
        ,input  [31:0]	int_desc_4_xuser_7_xuser
        ,input  [31:0]	int_desc_4_xuser_8_xuser
        ,input  [31:0]	int_desc_4_xuser_9_xuser
        ,input  [31:0]	int_desc_4_xuser_10_xuser
        ,input  [31:0]	int_desc_4_xuser_11_xuser
        ,input  [31:0]	int_desc_4_xuser_12_xuser
        ,input  [31:0]	int_desc_4_xuser_13_xuser
        ,input  [31:0]	int_desc_4_xuser_14_xuser
        ,input  [31:0]	int_desc_4_xuser_15_xuser
        ,input  [31:0]	int_desc_5_xuser_0_xuser
        ,input  [31:0]	int_desc_5_xuser_1_xuser
        ,input  [31:0]	int_desc_5_xuser_2_xuser
        ,input  [31:0]	int_desc_5_xuser_3_xuser
        ,input  [31:0]	int_desc_5_xuser_4_xuser
        ,input  [31:0]	int_desc_5_xuser_5_xuser
        ,input  [31:0]	int_desc_5_xuser_6_xuser
        ,input  [31:0]	int_desc_5_xuser_7_xuser
        ,input  [31:0]	int_desc_5_xuser_8_xuser
        ,input  [31:0]	int_desc_5_xuser_9_xuser
        ,input  [31:0]	int_desc_5_xuser_10_xuser
        ,input  [31:0]	int_desc_5_xuser_11_xuser
        ,input  [31:0]	int_desc_5_xuser_12_xuser
        ,input  [31:0]	int_desc_5_xuser_13_xuser
        ,input  [31:0]	int_desc_5_xuser_14_xuser
        ,input  [31:0]	int_desc_5_xuser_15_xuser
        ,input  [31:0]	int_desc_6_xuser_0_xuser
        ,input  [31:0]	int_desc_6_xuser_1_xuser
        ,input  [31:0]	int_desc_6_xuser_2_xuser
        ,input  [31:0]	int_desc_6_xuser_3_xuser
        ,input  [31:0]	int_desc_6_xuser_4_xuser
        ,input  [31:0]	int_desc_6_xuser_5_xuser
        ,input  [31:0]	int_desc_6_xuser_6_xuser
        ,input  [31:0]	int_desc_6_xuser_7_xuser
        ,input  [31:0]	int_desc_6_xuser_8_xuser
        ,input  [31:0]	int_desc_6_xuser_9_xuser
        ,input  [31:0]	int_desc_6_xuser_10_xuser
        ,input  [31:0]	int_desc_6_xuser_11_xuser
        ,input  [31:0]	int_desc_6_xuser_12_xuser
        ,input  [31:0]	int_desc_6_xuser_13_xuser
        ,input  [31:0]	int_desc_6_xuser_14_xuser
        ,input  [31:0]	int_desc_6_xuser_15_xuser
        ,input  [31:0]	int_desc_7_xuser_0_xuser
        ,input  [31:0]	int_desc_7_xuser_1_xuser
        ,input  [31:0]	int_desc_7_xuser_2_xuser
        ,input  [31:0]	int_desc_7_xuser_3_xuser
        ,input  [31:0]	int_desc_7_xuser_4_xuser
        ,input  [31:0]	int_desc_7_xuser_5_xuser
        ,input  [31:0]	int_desc_7_xuser_6_xuser
        ,input  [31:0]	int_desc_7_xuser_7_xuser
        ,input  [31:0]	int_desc_7_xuser_8_xuser
        ,input  [31:0]	int_desc_7_xuser_9_xuser
        ,input  [31:0]	int_desc_7_xuser_10_xuser
        ,input  [31:0]	int_desc_7_xuser_11_xuser
        ,input  [31:0]	int_desc_7_xuser_12_xuser
        ,input  [31:0]	int_desc_7_xuser_13_xuser
        ,input  [31:0]	int_desc_7_xuser_14_xuser
        ,input  [31:0]	int_desc_7_xuser_15_xuser
        ,input  [31:0]	int_desc_8_xuser_0_xuser
        ,input  [31:0]	int_desc_8_xuser_1_xuser
        ,input  [31:0]	int_desc_8_xuser_2_xuser
        ,input  [31:0]	int_desc_8_xuser_3_xuser
        ,input  [31:0]	int_desc_8_xuser_4_xuser
        ,input  [31:0]	int_desc_8_xuser_5_xuser
        ,input  [31:0]	int_desc_8_xuser_6_xuser
        ,input  [31:0]	int_desc_8_xuser_7_xuser
        ,input  [31:0]	int_desc_8_xuser_8_xuser
        ,input  [31:0]	int_desc_8_xuser_9_xuser
        ,input  [31:0]	int_desc_8_xuser_10_xuser
        ,input  [31:0]	int_desc_8_xuser_11_xuser
        ,input  [31:0]	int_desc_8_xuser_12_xuser
        ,input  [31:0]	int_desc_8_xuser_13_xuser
        ,input  [31:0]	int_desc_8_xuser_14_xuser
        ,input  [31:0]	int_desc_8_xuser_15_xuser
        ,input  [31:0]	int_desc_9_xuser_0_xuser
        ,input  [31:0]	int_desc_9_xuser_1_xuser
        ,input  [31:0]	int_desc_9_xuser_2_xuser
        ,input  [31:0]	int_desc_9_xuser_3_xuser
        ,input  [31:0]	int_desc_9_xuser_4_xuser
        ,input  [31:0]	int_desc_9_xuser_5_xuser
        ,input  [31:0]	int_desc_9_xuser_6_xuser
        ,input  [31:0]	int_desc_9_xuser_7_xuser
        ,input  [31:0]	int_desc_9_xuser_8_xuser
        ,input  [31:0]	int_desc_9_xuser_9_xuser
        ,input  [31:0]	int_desc_9_xuser_10_xuser
        ,input  [31:0]	int_desc_9_xuser_11_xuser
        ,input  [31:0]	int_desc_9_xuser_12_xuser
        ,input  [31:0]	int_desc_9_xuser_13_xuser
        ,input  [31:0]	int_desc_9_xuser_14_xuser
        ,input  [31:0]	int_desc_9_xuser_15_xuser
        ,input  [31:0]	int_desc_10_xuser_0_xuser
        ,input  [31:0]	int_desc_10_xuser_1_xuser
        ,input  [31:0]	int_desc_10_xuser_2_xuser
        ,input  [31:0]	int_desc_10_xuser_3_xuser
        ,input  [31:0]	int_desc_10_xuser_4_xuser
        ,input  [31:0]	int_desc_10_xuser_5_xuser
        ,input  [31:0]	int_desc_10_xuser_6_xuser
        ,input  [31:0]	int_desc_10_xuser_7_xuser
        ,input  [31:0]	int_desc_10_xuser_8_xuser
        ,input  [31:0]	int_desc_10_xuser_9_xuser
        ,input  [31:0]	int_desc_10_xuser_10_xuser
        ,input  [31:0]	int_desc_10_xuser_11_xuser
        ,input  [31:0]	int_desc_10_xuser_12_xuser
        ,input  [31:0]	int_desc_10_xuser_13_xuser
        ,input  [31:0]	int_desc_10_xuser_14_xuser
        ,input  [31:0]	int_desc_10_xuser_15_xuser
        ,input  [31:0]	int_desc_11_xuser_0_xuser
        ,input  [31:0]	int_desc_11_xuser_1_xuser
        ,input  [31:0]	int_desc_11_xuser_2_xuser
        ,input  [31:0]	int_desc_11_xuser_3_xuser
        ,input  [31:0]	int_desc_11_xuser_4_xuser
        ,input  [31:0]	int_desc_11_xuser_5_xuser
        ,input  [31:0]	int_desc_11_xuser_6_xuser
        ,input  [31:0]	int_desc_11_xuser_7_xuser
        ,input  [31:0]	int_desc_11_xuser_8_xuser
        ,input  [31:0]	int_desc_11_xuser_9_xuser
        ,input  [31:0]	int_desc_11_xuser_10_xuser
        ,input  [31:0]	int_desc_11_xuser_11_xuser
        ,input  [31:0]	int_desc_11_xuser_12_xuser
        ,input  [31:0]	int_desc_11_xuser_13_xuser
        ,input  [31:0]	int_desc_11_xuser_14_xuser
        ,input  [31:0]	int_desc_11_xuser_15_xuser
        ,input  [31:0]	int_desc_12_xuser_0_xuser
        ,input  [31:0]	int_desc_12_xuser_1_xuser
        ,input  [31:0]	int_desc_12_xuser_2_xuser
        ,input  [31:0]	int_desc_12_xuser_3_xuser
        ,input  [31:0]	int_desc_12_xuser_4_xuser
        ,input  [31:0]	int_desc_12_xuser_5_xuser
        ,input  [31:0]	int_desc_12_xuser_6_xuser
        ,input  [31:0]	int_desc_12_xuser_7_xuser
        ,input  [31:0]	int_desc_12_xuser_8_xuser
        ,input  [31:0]	int_desc_12_xuser_9_xuser
        ,input  [31:0]	int_desc_12_xuser_10_xuser
        ,input  [31:0]	int_desc_12_xuser_11_xuser
        ,input  [31:0]	int_desc_12_xuser_12_xuser
        ,input  [31:0]	int_desc_12_xuser_13_xuser
        ,input  [31:0]	int_desc_12_xuser_14_xuser
        ,input  [31:0]	int_desc_12_xuser_15_xuser
        ,input  [31:0]	int_desc_13_xuser_0_xuser
        ,input  [31:0]	int_desc_13_xuser_1_xuser
        ,input  [31:0]	int_desc_13_xuser_2_xuser
        ,input  [31:0]	int_desc_13_xuser_3_xuser
        ,input  [31:0]	int_desc_13_xuser_4_xuser
        ,input  [31:0]	int_desc_13_xuser_5_xuser
        ,input  [31:0]	int_desc_13_xuser_6_xuser
        ,input  [31:0]	int_desc_13_xuser_7_xuser
        ,input  [31:0]	int_desc_13_xuser_8_xuser
        ,input  [31:0]	int_desc_13_xuser_9_xuser
        ,input  [31:0]	int_desc_13_xuser_10_xuser
        ,input  [31:0]	int_desc_13_xuser_11_xuser
        ,input  [31:0]	int_desc_13_xuser_12_xuser
        ,input  [31:0]	int_desc_13_xuser_13_xuser
        ,input  [31:0]	int_desc_13_xuser_14_xuser
        ,input  [31:0]	int_desc_13_xuser_15_xuser
        ,input  [31:0]	int_desc_14_xuser_0_xuser
        ,input  [31:0]	int_desc_14_xuser_1_xuser
        ,input  [31:0]	int_desc_14_xuser_2_xuser
        ,input  [31:0]	int_desc_14_xuser_3_xuser
        ,input  [31:0]	int_desc_14_xuser_4_xuser
        ,input  [31:0]	int_desc_14_xuser_5_xuser
        ,input  [31:0]	int_desc_14_xuser_6_xuser
        ,input  [31:0]	int_desc_14_xuser_7_xuser
        ,input  [31:0]	int_desc_14_xuser_8_xuser
        ,input  [31:0]	int_desc_14_xuser_9_xuser
        ,input  [31:0]	int_desc_14_xuser_10_xuser
        ,input  [31:0]	int_desc_14_xuser_11_xuser
        ,input  [31:0]	int_desc_14_xuser_12_xuser
        ,input  [31:0]	int_desc_14_xuser_13_xuser
        ,input  [31:0]	int_desc_14_xuser_14_xuser
        ,input  [31:0]	int_desc_14_xuser_15_xuser
        ,input  [31:0]	int_desc_15_xuser_0_xuser
        ,input  [31:0]	int_desc_15_xuser_1_xuser
        ,input  [31:0]	int_desc_15_xuser_2_xuser
        ,input  [31:0]	int_desc_15_xuser_3_xuser
        ,input  [31:0]	int_desc_15_xuser_4_xuser
        ,input  [31:0]	int_desc_15_xuser_5_xuser
        ,input  [31:0]	int_desc_15_xuser_6_xuser
        ,input  [31:0]	int_desc_15_xuser_7_xuser
        ,input  [31:0]	int_desc_15_xuser_8_xuser
        ,input  [31:0]	int_desc_15_xuser_9_xuser
        ,input  [31:0]	int_desc_15_xuser_10_xuser
        ,input  [31:0]	int_desc_15_xuser_11_xuser
        ,input  [31:0]	int_desc_15_xuser_12_xuser
        ,input  [31:0]	int_desc_15_xuser_13_xuser
        ,input  [31:0]	int_desc_15_xuser_14_xuser
        ,input  [31:0]	int_desc_15_xuser_15_xuser
