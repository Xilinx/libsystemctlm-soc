`timescale 1ns / 1ps

`include "include/axi.svh"

module axilite_dev_dpi(
	input clk,
	input resetn);

	`AXILITE_NETS(m00, 32, 32);

	axilite_dev axidev(.s00_axi_aclk(clk), .s00_axi_aresetn(resetn),
		`AXILITE_CONNECT_PORT(s00_axi_, m00_));


   initial begin
      if ($test$plusargs("trace") != 0) begin
         $display("[%0t] Tracing to logs/vlt_dump.vcd...\n", $time);
         $dumpfile("logs/vlt_dump.vcd");
         $dumpvars();
      end
      $display("[%0t] Model running...\n", $time);
   end


endmodule
