/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */

// OFFSET ADDR of REGS
`define BRIDGE_IDENTIFICATION_REG_ADDR 'h0
`define LAST_BRIDGE_REG_ADDR 'h4
`define VERSION_REG_ADDR 'h20
`define BRIDGE_TYPE_REG_ADDR 'h24
`define MODE_SELECT_REG_ADDR 'h38
`define RESET_REG_ADDR 'h3C
`define H2C_INTR_0_REG_ADDR 'h40
`define H2C_INTR_1_REG_ADDR 'h44
`define H2C_INTR_2_REG_ADDR 'h48
`define H2C_INTR_3_REG_ADDR 'h4C
`define C2H_INTR_STATUS_0_REG_ADDR 'h60
`define INTR_C2H_TOGGLE_STATUS_0_REG_ADDR 'h64
`define INTR_C2H_TOGGLE_CLEAR_0_REG_ADDR 'h68
`define INTR_C2H_TOGGLE_ENABLE_0_REG_ADDR 'h6C
`define C2H_INTR_STATUS_1_REG_ADDR 'h70
`define INTR_C2H_TOGGLE_STATUS_1_REG_ADDR 'h74
`define INTR_C2H_TOGGLE_CLEAR_1_REG_ADDR 'h78
`define INTR_C2H_TOGGLE_ENABLE_1_REG_ADDR 'h7C
`define C2H_GPIO_0_REG_ADDR 'h80
`define C2H_GPIO_1_REG_ADDR 'h84
`define C2H_GPIO_2_REG_ADDR 'h88
`define C2H_GPIO_3_REG_ADDR 'h8C
`define C2H_GPIO_4_REG_ADDR 'h90
`define C2H_GPIO_5_REG_ADDR 'h94
`define C2H_GPIO_6_REG_ADDR 'h98
`define C2H_GPIO_7_REG_ADDR 'h9C
`define C2H_GPIO_8_REG_ADDR 'hA0
`define C2H_GPIO_9_REG_ADDR 'hA4
`define C2H_GPIO_10_REG_ADDR 'hA8
`define C2H_GPIO_11_REG_ADDR 'hAC
`define C2H_GPIO_12_REG_ADDR 'hB0
`define C2H_GPIO_13_REG_ADDR 'hB4
`define C2H_GPIO_14_REG_ADDR 'hB8
`define C2H_GPIO_15_REG_ADDR 'hBC
`define H2C_GPIO_0_REG_ADDR 'hC0
`define H2C_GPIO_1_REG_ADDR 'hC4
`define H2C_GPIO_2_REG_ADDR 'hC8
`define H2C_GPIO_3_REG_ADDR 'hCC
`define H2C_GPIO_4_REG_ADDR 'hD0
`define H2C_GPIO_5_REG_ADDR 'hD4
`define H2C_GPIO_6_REG_ADDR 'hD8
`define H2C_GPIO_7_REG_ADDR 'hDC
`define H2C_GPIO_8_REG_ADDR 'hE0
`define H2C_GPIO_9_REG_ADDR 'hE4
`define H2C_GPIO_10_REG_ADDR 'hE8
`define H2C_GPIO_11_REG_ADDR 'hEC
`define H2C_GPIO_12_REG_ADDR 'hF0
`define H2C_GPIO_13_REG_ADDR 'hF4
`define H2C_GPIO_14_REG_ADDR 'hF8
`define H2C_GPIO_15_REG_ADDR 'hFC
`define BRIDGE_CONFIG_REG_ADDR 'h200
`define INTR_STATUS_REG_ADDR 'h208
`define INTR_ERROR_STATUS_REG_ADDR 'h20C
`define INTR_ERROR_CLEAR_REG_ADDR 'h210
`define INTR_ERROR_ENABLE_REG_ADDR 'h214
`define BRIDGE_RD_USER_CONFIG_REG_ADDR 'h218
`define BRIDGE_WR_USER_CONFIG_REG_ADDR 'h21C
`define RD_MAX_DESC_REG_ADDR 'h220
`define WR_MAX_DESC_REG_ADDR 'h224
`define SN_MAX_DESC_REG_ADDR 'h228
`define RD_REQ_FIFO_PUSH_DESC_REG_ADDR 'h300
`define RD_REQ_FIFO_FREE_LEVEL_REG_ADDR 'h304
`define RD_REQ_INTR_COMP_STATUS_REG_ADDR 'h308
`define RD_REQ_INTR_COMP_CLEAR_REG_ADDR 'h30C
`define RD_REQ_INTR_COMP_ENABLE_REG_ADDR 'h310
`define RD_RESP_FREE_DESC_REG_ADDR 'h314
`define RD_RESP_FIFO_POP_DESC_REG_ADDR 'h318
`define RD_RESP_FIFO_FILL_LEVEL_REG_ADDR 'h31C
`define WR_REQ_FIFO_PUSH_DESC_REG_ADDR 'h320
`define WR_REQ_FIFO_FREE_LEVEL_REG_ADDR 'h324
`define WR_REQ_INTR_COMP_STATUS_REG_ADDR 'h328
`define WR_REQ_INTR_COMP_CLEAR_REG_ADDR 'h32C
`define WR_REQ_INTR_COMP_ENABLE_REG_ADDR 'h330
`define WR_RESP_FREE_DESC_REG_ADDR 'h334
`define WR_RESP_FIFO_POP_DESC_REG_ADDR 'h338
`define WR_RESP_FIFO_FILL_LEVEL_REG_ADDR 'h33C
`define SN_REQ_FREE_DESC_REG_ADDR 'h340
`define SN_REQ_FIFO_POP_DESC_REG_ADDR 'h344
`define SN_REQ_FIFO_FILL_LEVEL_REG_ADDR 'h348
`define SN_RESP_FIFO_PUSH_DESC_REG_ADDR 'h34C
`define SN_RESP_FIFO_FREE_LEVEL_REG_ADDR 'h350
`define SN_RESP_INTR_COMP_STATUS_REG_ADDR 'h354
`define SN_RESP_INTR_COMP_CLEAR_REG_ADDR 'h358
`define SN_RESP_INTR_COMP_ENABLE_REG_ADDR 'h35C
`define SN_DATA_FIFO_PUSH_DESC_REG_ADDR 'h360
`define SN_DATA_FIFO_FREE_LEVEL_REG_ADDR 'h364
`define SN_DATA_INTR_COMP_STATUS_REG_ADDR 'h368
`define SN_DATA_INTR_COMP_CLEAR_REG_ADDR 'h36C
`define SN_DATA_INTR_COMP_ENABLE_REG_ADDR 'h370
`define INTR_FIFO_ENABLE_REG_ADDR 'h374


`define RD_REQ_DESC_N_BASE_ADDR 'h3000
`define RD_RESP_DESC_N_BASE_ADDR 'h4000
`define WR_REQ_DESC_N_BASE_ADDR 'h5000
`define WR_RESP_DESC_N_BASE_ADDR 'h6000
`define SN_REQ_DESC_N_BASE_ADDR 'h7000
`define SN_RESP_DESC_N_BASE_ADDR 'h7200
`define RD_REQ_DESC_0_BASE_ADDR 'h3000
`define RD_RESP_DESC_0_BASE_ADDR 'h4000
`define WR_REQ_DESC_0_BASE_ADDR 'h5000
`define WR_RESP_DESC_0_BASE_ADDR 'h6000
`define RD_REQ_DESC_1_BASE_ADDR 'h3100
`define RD_REQ_DESC_2_BASE_ADDR 'h3200
`define RD_REQ_DESC_3_BASE_ADDR 'h3300
`define RD_REQ_DESC_4_BASE_ADDR 'h3400
`define RD_REQ_DESC_5_BASE_ADDR 'h3500
`define RD_REQ_DESC_6_BASE_ADDR 'h3600
`define RD_REQ_DESC_7_BASE_ADDR 'h3700
`define RD_REQ_DESC_8_BASE_ADDR 'h3800
`define RD_REQ_DESC_9_BASE_ADDR 'h3900
`define RD_REQ_DESC_A_BASE_ADDR 'h3A00
`define RD_REQ_DESC_B_BASE_ADDR 'h3B00
`define RD_REQ_DESC_C_BASE_ADDR 'h3C00
`define RD_REQ_DESC_D_BASE_ADDR 'h3D00
`define RD_REQ_DESC_E_BASE_ADDR 'h3E00
`define RD_REQ_DESC_F_BASE_ADDR 'h3F00
`define RD_RESP_DESC_1_BASE_ADDR 'h4100
`define RD_RESP_DESC_2_BASE_ADDR 'h4200
`define RD_RESP_DESC_3_BASE_ADDR 'h4300
`define RD_RESP_DESC_4_BASE_ADDR 'h4400
`define RD_RESP_DESC_5_BASE_ADDR 'h4500
`define RD_RESP_DESC_6_BASE_ADDR 'h4600
`define RD_RESP_DESC_7_BASE_ADDR 'h4700
`define RD_RESP_DESC_8_BASE_ADDR 'h4800
`define RD_RESP_DESC_9_BASE_ADDR 'h4900
`define RD_RESP_DESC_A_BASE_ADDR 'h4A00
`define RD_RESP_DESC_B_BASE_ADDR 'h4B00
`define RD_RESP_DESC_C_BASE_ADDR 'h4C00
`define RD_RESP_DESC_D_BASE_ADDR 'h4D00
`define RD_RESP_DESC_E_BASE_ADDR 'h4E00
`define RD_RESP_DESC_F_BASE_ADDR 'h4F00
`define WR_REQ_DESC_1_BASE_ADDR 'h5100
`define WR_REQ_DESC_2_BASE_ADDR 'h5200
`define WR_REQ_DESC_3_BASE_ADDR 'h5300
`define WR_REQ_DESC_4_BASE_ADDR 'h5400
`define WR_REQ_DESC_5_BASE_ADDR 'h5500
`define WR_REQ_DESC_6_BASE_ADDR 'h5600
`define WR_REQ_DESC_7_BASE_ADDR 'h5700
`define WR_REQ_DESC_8_BASE_ADDR 'h5800
`define WR_REQ_DESC_9_BASE_ADDR 'h5900
`define WR_REQ_DESC_A_BASE_ADDR 'h5A00
`define WR_REQ_DESC_B_BASE_ADDR 'h5B00
`define WR_REQ_DESC_C_BASE_ADDR 'h5C00
`define WR_REQ_DESC_D_BASE_ADDR 'h5D00
`define WR_REQ_DESC_E_BASE_ADDR 'h5E00
`define WR_REQ_DESC_F_BASE_ADDR 'h5F00
`define WR_RESP_DESC_1_BASE_ADDR 'h6100
`define WR_RESP_DESC_2_BASE_ADDR 'h6200
`define WR_RESP_DESC_3_BASE_ADDR 'h6300
`define WR_RESP_DESC_4_BASE_ADDR 'h6400
`define WR_RESP_DESC_5_BASE_ADDR 'h6500
`define WR_RESP_DESC_6_BASE_ADDR 'h6600
`define WR_RESP_DESC_7_BASE_ADDR 'h6700
`define WR_RESP_DESC_8_BASE_ADDR 'h6800
`define WR_RESP_DESC_9_BASE_ADDR 'h6900
`define WR_RESP_DESC_A_BASE_ADDR 'h6A00
`define WR_RESP_DESC_B_BASE_ADDR 'h6B00
`define WR_RESP_DESC_C_BASE_ADDR 'h6C00
`define WR_RESP_DESC_D_BASE_ADDR 'h6D00
`define WR_RESP_DESC_E_BASE_ADDR 'h6E00
`define WR_RESP_DESC_F_BASE_ADDR 'h6F00
`define SN_REQ_DESC_0_BASE_ADDR 'h7000
`define SN_RESP_DESC_0_BASE_ADDR 'h7200
`define SN_REQ_DESC_1_BASE_ADDR 'h7020
`define SN_REQ_DESC_2_BASE_ADDR 'h7040
`define SN_REQ_DESC_3_BASE_ADDR 'h7060
`define SN_REQ_DESC_4_BASE_ADDR 'h7080
`define SN_REQ_DESC_5_BASE_ADDR 'h70A0
`define SN_REQ_DESC_6_BASE_ADDR 'h70C0
`define SN_REQ_DESC_7_BASE_ADDR 'h70E0
`define SN_REQ_DESC_8_BASE_ADDR 'h7100
`define SN_REQ_DESC_9_BASE_ADDR 'h7120
`define SN_REQ_DESC_A_BASE_ADDR 'h7140
`define SN_REQ_DESC_B_BASE_ADDR 'h7160
`define SN_REQ_DESC_C_BASE_ADDR 'h7180
`define SN_REQ_DESC_D_BASE_ADDR 'h71A0
`define SN_REQ_DESC_E_BASE_ADDR 'h71C0
`define SN_REQ_DESC_F_BASE_ADDR 'h71E0
`define SN_RESP_DESC_1_BASE_ADDR 'h7220
`define SN_RESP_DESC_2_BASE_ADDR 'h7240
`define SN_RESP_DESC_3_BASE_ADDR 'h7260
`define SN_RESP_DESC_4_BASE_ADDR 'h7280
`define SN_RESP_DESC_5_BASE_ADDR 'h72A0
`define SN_RESP_DESC_6_BASE_ADDR 'h72C0
`define SN_RESP_DESC_7_BASE_ADDR 'h72E0
`define SN_RESP_DESC_8_BASE_ADDR 'h7300
`define SN_RESP_DESC_9_BASE_ADDR 'h7320
`define SN_RESP_DESC_A_BASE_ADDR 'h7340
`define SN_RESP_DESC_B_BASE_ADDR 'h7360
`define SN_RESP_DESC_C_BASE_ADDR 'h7380
`define SN_RESP_DESC_D_BASE_ADDR 'h73A0
`define SN_RESP_DESC_E_BASE_ADDR 'h73C0
`define SN_RESP_DESC_F_BASE_ADDR 'h73E0
`define XX_DESCSIZE 'h100
`define SN_DESCSIZE 'h20


`define RD_REQ_DESC_N_TXN_TYPE_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h0
`define RD_REQ_DESC_N_SIZE_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h4
`define RD_REQ_DESC_N_AXSIZE_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h8
`define RD_REQ_DESC_N_ATTR_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'hC
`define RD_REQ_DESC_N_AXADDR_0_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h10
`define RD_REQ_DESC_N_AXADDR_1_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h14
`define RD_REQ_DESC_N_AXADDR_2_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h18
`define RD_REQ_DESC_N_AXADDR_3_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h1C
`define RD_REQ_DESC_N_AXID_0_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h20
`define RD_REQ_DESC_N_AXID_1_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h24
`define RD_REQ_DESC_N_AXID_2_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h28
`define RD_REQ_DESC_N_AXID_3_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h2C
`define RD_REQ_DESC_N_AXUSER_0_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h30
`define RD_REQ_DESC_N_AXUSER_1_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h34
`define RD_REQ_DESC_N_AXUSER_2_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h38
`define RD_REQ_DESC_N_AXUSER_3_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h3C
`define RD_REQ_DESC_N_AXUSER_4_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h40
`define RD_REQ_DESC_N_AXUSER_5_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h44
`define RD_REQ_DESC_N_AXUSER_6_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h48
`define RD_REQ_DESC_N_AXUSER_7_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h4C
`define RD_REQ_DESC_N_AXUSER_8_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h50
`define RD_REQ_DESC_N_AXUSER_9_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h54
`define RD_REQ_DESC_N_AXUSER_10_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h58
`define RD_REQ_DESC_N_AXUSER_11_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h5C
`define RD_REQ_DESC_N_AXUSER_12_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h60
`define RD_REQ_DESC_N_AXUSER_13_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h64
`define RD_REQ_DESC_N_AXUSER_14_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h68
`define RD_REQ_DESC_N_AXUSER_15_REG_ADDR `RD_REQ_DESC_N_BASE_ADDR + 'h6C
`define RD_RESP_DESC_N_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h0
`define RD_RESP_DESC_N_DATA_SIZE_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h4
`define RD_RESP_DESC_N_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h8
`define RD_RESP_DESC_N_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'hC
`define RD_RESP_DESC_N_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h10
`define RD_RESP_DESC_N_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h14
`define RD_RESP_DESC_N_RESP_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h18
`define RD_RESP_DESC_N_XID_0_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h1C
`define RD_RESP_DESC_N_XID_1_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h20
`define RD_RESP_DESC_N_XID_2_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h24
`define RD_RESP_DESC_N_XID_3_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h28
`define RD_RESP_DESC_N_XUSER_0_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h2C
`define RD_RESP_DESC_N_XUSER_1_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h30
`define RD_RESP_DESC_N_XUSER_2_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h34
`define RD_RESP_DESC_N_XUSER_3_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h38
`define RD_RESP_DESC_N_XUSER_4_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h3C
`define RD_RESP_DESC_N_XUSER_5_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h40
`define RD_RESP_DESC_N_XUSER_6_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h44
`define RD_RESP_DESC_N_XUSER_7_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h48
`define RD_RESP_DESC_N_XUSER_8_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h4C
`define RD_RESP_DESC_N_XUSER_9_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h50
`define RD_RESP_DESC_N_XUSER_10_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h54
`define RD_RESP_DESC_N_XUSER_11_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h58
`define RD_RESP_DESC_N_XUSER_12_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h5C
`define RD_RESP_DESC_N_XUSER_13_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h60
`define RD_RESP_DESC_N_XUSER_14_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h64
`define RD_RESP_DESC_N_XUSER_15_REG_ADDR `RD_RESP_DESC_N_BASE_ADDR + 'h68
`define WR_REQ_DESC_N_TXN_TYPE_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h0
`define WR_REQ_DESC_N_SIZE_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h4
`define WR_REQ_DESC_N_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h8
`define WR_REQ_DESC_N_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hC
`define WR_REQ_DESC_N_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h10
`define WR_REQ_DESC_N_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h14
`define WR_REQ_DESC_N_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h18
`define WR_REQ_DESC_N_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h1C
`define WR_REQ_DESC_N_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h20
`define WR_REQ_DESC_N_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h24
`define WR_REQ_DESC_N_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h28
`define WR_REQ_DESC_N_AXSIZE_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h2C
`define WR_REQ_DESC_N_ATTR_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h30
`define WR_REQ_DESC_N_AXADDR_0_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h34
`define WR_REQ_DESC_N_AXADDR_1_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h38
`define WR_REQ_DESC_N_AXADDR_2_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h3C
`define WR_REQ_DESC_N_AXADDR_3_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h40
`define WR_REQ_DESC_N_AXID_0_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h44
`define WR_REQ_DESC_N_AXID_1_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h48
`define WR_REQ_DESC_N_AXID_2_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h4C
`define WR_REQ_DESC_N_AXID_3_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h50
`define WR_REQ_DESC_N_AXUSER_0_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h54
`define WR_REQ_DESC_N_AXUSER_1_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h58
`define WR_REQ_DESC_N_AXUSER_2_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h5C
`define WR_REQ_DESC_N_AXUSER_3_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h60
`define WR_REQ_DESC_N_AXUSER_4_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h64
`define WR_REQ_DESC_N_AXUSER_5_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h68
`define WR_REQ_DESC_N_AXUSER_6_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h6C
`define WR_REQ_DESC_N_AXUSER_7_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h70
`define WR_REQ_DESC_N_AXUSER_8_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h74
`define WR_REQ_DESC_N_AXUSER_9_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h78
`define WR_REQ_DESC_N_AXUSER_10_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h7C
`define WR_REQ_DESC_N_AXUSER_11_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h80
`define WR_REQ_DESC_N_AXUSER_12_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h84
`define WR_REQ_DESC_N_AXUSER_13_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h88
`define WR_REQ_DESC_N_AXUSER_14_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h8C
`define WR_REQ_DESC_N_AXUSER_15_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h90
`define WR_REQ_DESC_N_WUSER_0_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h94
`define WR_REQ_DESC_N_WUSER_1_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h98
`define WR_REQ_DESC_N_WUSER_2_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'h9C
`define WR_REQ_DESC_N_WUSER_3_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hA0
`define WR_REQ_DESC_N_WUSER_4_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hA4
`define WR_REQ_DESC_N_WUSER_5_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hA8
`define WR_REQ_DESC_N_WUSER_6_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hAC
`define WR_REQ_DESC_N_WUSER_7_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hB0
`define WR_REQ_DESC_N_WUSER_8_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hB4
`define WR_REQ_DESC_N_WUSER_9_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hB8
`define WR_REQ_DESC_N_WUSER_10_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hBC
`define WR_REQ_DESC_N_WUSER_11_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hC0
`define WR_REQ_DESC_N_WUSER_12_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hC4
`define WR_REQ_DESC_N_WUSER_13_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hC8
`define WR_REQ_DESC_N_WUSER_14_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hCC
`define WR_REQ_DESC_N_WUSER_15_REG_ADDR `WR_REQ_DESC_N_BASE_ADDR + 'hD0
`define WR_RESP_DESC_N_RESP_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h0
`define WR_RESP_DESC_N_XID_0_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h4
`define WR_RESP_DESC_N_XID_1_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h8
`define WR_RESP_DESC_N_XID_2_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'hC
`define WR_RESP_DESC_N_XID_3_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h10
`define WR_RESP_DESC_N_XUSER_0_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h14
`define WR_RESP_DESC_N_XUSER_1_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h18
`define WR_RESP_DESC_N_XUSER_2_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h1C
`define WR_RESP_DESC_N_XUSER_3_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h20
`define WR_RESP_DESC_N_XUSER_4_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h24
`define WR_RESP_DESC_N_XUSER_5_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h28
`define WR_RESP_DESC_N_XUSER_6_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h2C
`define WR_RESP_DESC_N_XUSER_7_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h30
`define WR_RESP_DESC_N_XUSER_8_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h34
`define WR_RESP_DESC_N_XUSER_9_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h38
`define WR_RESP_DESC_N_XUSER_10_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h3C
`define WR_RESP_DESC_N_XUSER_11_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h40
`define WR_RESP_DESC_N_XUSER_12_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h44
`define WR_RESP_DESC_N_XUSER_13_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h48
`define WR_RESP_DESC_N_XUSER_14_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h4C
`define WR_RESP_DESC_N_XUSER_15_REG_ADDR `WR_RESP_DESC_N_BASE_ADDR + 'h50
`define SN_REQ_DESC_N_ATTR_REG_ADDR `SN_REQ_DESC_N_BASE_ADDR + 'h0
`define SN_REQ_DESC_N_ACADDR_0_REG_ADDR `SN_REQ_DESC_N_BASE_ADDR + 'h4
`define SN_REQ_DESC_N_ACADDR_1_REG_ADDR `SN_REQ_DESC_N_BASE_ADDR + 'h8
`define SN_REQ_DESC_N_ACADDR_2_REG_ADDR `SN_REQ_DESC_N_BASE_ADDR + 'hC
`define SN_REQ_DESC_N_ACADDR_3_REG_ADDR `SN_REQ_DESC_N_BASE_ADDR + 'h10
`define SN_RESP_DESC_N_RESP_REG_ADDR `SN_RESP_DESC_N_BASE_ADDR + 'h0


`define RD_REQ_DESC_0_TXN_TYPE_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h0
`define RD_REQ_DESC_0_SIZE_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h4
`define RD_REQ_DESC_0_AXSIZE_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h8
`define RD_REQ_DESC_0_ATTR_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'hC
`define RD_REQ_DESC_0_AXADDR_0_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h10
`define RD_REQ_DESC_0_AXADDR_1_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h14
`define RD_REQ_DESC_0_AXADDR_2_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h18
`define RD_REQ_DESC_0_AXADDR_3_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h1C
`define RD_REQ_DESC_0_AXID_0_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h20
`define RD_REQ_DESC_0_AXID_1_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h24
`define RD_REQ_DESC_0_AXID_2_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h28
`define RD_REQ_DESC_0_AXID_3_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h2C
`define RD_REQ_DESC_0_AXUSER_0_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h30
`define RD_REQ_DESC_0_AXUSER_1_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h34
`define RD_REQ_DESC_0_AXUSER_2_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h38
`define RD_REQ_DESC_0_AXUSER_3_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h3C
`define RD_REQ_DESC_0_AXUSER_4_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h40
`define RD_REQ_DESC_0_AXUSER_5_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h44
`define RD_REQ_DESC_0_AXUSER_6_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h48
`define RD_REQ_DESC_0_AXUSER_7_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h4C
`define RD_REQ_DESC_0_AXUSER_8_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h50
`define RD_REQ_DESC_0_AXUSER_9_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h54
`define RD_REQ_DESC_0_AXUSER_10_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h58
`define RD_REQ_DESC_0_AXUSER_11_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h5C
`define RD_REQ_DESC_0_AXUSER_12_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h60
`define RD_REQ_DESC_0_AXUSER_13_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h64
`define RD_REQ_DESC_0_AXUSER_14_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h68
`define RD_REQ_DESC_0_AXUSER_15_REG_ADDR `RD_REQ_DESC_0_BASE_ADDR + 'h6C
`define RD_RESP_DESC_0_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h0
`define RD_RESP_DESC_0_DATA_SIZE_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h4
`define RD_RESP_DESC_0_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h8
`define RD_RESP_DESC_0_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'hC
`define RD_RESP_DESC_0_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h10
`define RD_RESP_DESC_0_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h14
`define RD_RESP_DESC_0_RESP_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h18
`define RD_RESP_DESC_0_XID_0_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h1C
`define RD_RESP_DESC_0_XID_1_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h20
`define RD_RESP_DESC_0_XID_2_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h24
`define RD_RESP_DESC_0_XID_3_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h28
`define RD_RESP_DESC_0_XUSER_0_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h2C
`define RD_RESP_DESC_0_XUSER_1_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h30
`define RD_RESP_DESC_0_XUSER_2_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h34
`define RD_RESP_DESC_0_XUSER_3_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h38
`define RD_RESP_DESC_0_XUSER_4_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h3C
`define RD_RESP_DESC_0_XUSER_5_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h40
`define RD_RESP_DESC_0_XUSER_6_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h44
`define RD_RESP_DESC_0_XUSER_7_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h48
`define RD_RESP_DESC_0_XUSER_8_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h4C
`define RD_RESP_DESC_0_XUSER_9_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h50
`define RD_RESP_DESC_0_XUSER_10_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h54
`define RD_RESP_DESC_0_XUSER_11_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h58
`define RD_RESP_DESC_0_XUSER_12_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h5C
`define RD_RESP_DESC_0_XUSER_13_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h60
`define RD_RESP_DESC_0_XUSER_14_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h64
`define RD_RESP_DESC_0_XUSER_15_REG_ADDR `RD_RESP_DESC_0_BASE_ADDR + 'h68
`define WR_REQ_DESC_0_TXN_TYPE_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h0
`define WR_REQ_DESC_0_SIZE_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h4
`define WR_REQ_DESC_0_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h8
`define WR_REQ_DESC_0_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hC
`define WR_REQ_DESC_0_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h10
`define WR_REQ_DESC_0_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h14
`define WR_REQ_DESC_0_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h18
`define WR_REQ_DESC_0_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h1C
`define WR_REQ_DESC_0_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h20
`define WR_REQ_DESC_0_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h24
`define WR_REQ_DESC_0_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h28
`define WR_REQ_DESC_0_AXSIZE_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h2C
`define WR_REQ_DESC_0_ATTR_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h30
`define WR_REQ_DESC_0_AXADDR_0_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h34
`define WR_REQ_DESC_0_AXADDR_1_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h38
`define WR_REQ_DESC_0_AXADDR_2_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h3C
`define WR_REQ_DESC_0_AXADDR_3_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h40
`define WR_REQ_DESC_0_AXID_0_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h44
`define WR_REQ_DESC_0_AXID_1_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h48
`define WR_REQ_DESC_0_AXID_2_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h4C
`define WR_REQ_DESC_0_AXID_3_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h50
`define WR_REQ_DESC_0_AXUSER_0_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h54
`define WR_REQ_DESC_0_AXUSER_1_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h58
`define WR_REQ_DESC_0_AXUSER_2_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h5C
`define WR_REQ_DESC_0_AXUSER_3_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h60
`define WR_REQ_DESC_0_AXUSER_4_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h64
`define WR_REQ_DESC_0_AXUSER_5_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h68
`define WR_REQ_DESC_0_AXUSER_6_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h6C
`define WR_REQ_DESC_0_AXUSER_7_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h70
`define WR_REQ_DESC_0_AXUSER_8_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h74
`define WR_REQ_DESC_0_AXUSER_9_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h78
`define WR_REQ_DESC_0_AXUSER_10_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h7C
`define WR_REQ_DESC_0_AXUSER_11_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h80
`define WR_REQ_DESC_0_AXUSER_12_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h84
`define WR_REQ_DESC_0_AXUSER_13_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h88
`define WR_REQ_DESC_0_AXUSER_14_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h8C
`define WR_REQ_DESC_0_AXUSER_15_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h90
`define WR_REQ_DESC_0_WUSER_0_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h94
`define WR_REQ_DESC_0_WUSER_1_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h98
`define WR_REQ_DESC_0_WUSER_2_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'h9C
`define WR_REQ_DESC_0_WUSER_3_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hA0
`define WR_REQ_DESC_0_WUSER_4_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hA4
`define WR_REQ_DESC_0_WUSER_5_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hA8
`define WR_REQ_DESC_0_WUSER_6_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hAC
`define WR_REQ_DESC_0_WUSER_7_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hB0
`define WR_REQ_DESC_0_WUSER_8_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hB4
`define WR_REQ_DESC_0_WUSER_9_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hB8
`define WR_REQ_DESC_0_WUSER_10_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hBC
`define WR_REQ_DESC_0_WUSER_11_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hC0
`define WR_REQ_DESC_0_WUSER_12_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hC4
`define WR_REQ_DESC_0_WUSER_13_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hC8
`define WR_REQ_DESC_0_WUSER_14_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hCC
`define WR_REQ_DESC_0_WUSER_15_REG_ADDR `WR_REQ_DESC_0_BASE_ADDR + 'hD0
`define WR_RESP_DESC_0_RESP_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h0
`define WR_RESP_DESC_0_XID_0_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h4
`define WR_RESP_DESC_0_XID_1_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h8
`define WR_RESP_DESC_0_XID_2_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'hC
`define WR_RESP_DESC_0_XID_3_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h10
`define WR_RESP_DESC_0_XUSER_0_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h14
`define WR_RESP_DESC_0_XUSER_1_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h18
`define WR_RESP_DESC_0_XUSER_2_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h1C
`define WR_RESP_DESC_0_XUSER_3_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h20
`define WR_RESP_DESC_0_XUSER_4_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h24
`define WR_RESP_DESC_0_XUSER_5_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h28
`define WR_RESP_DESC_0_XUSER_6_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h2C
`define WR_RESP_DESC_0_XUSER_7_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h30
`define WR_RESP_DESC_0_XUSER_8_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h34
`define WR_RESP_DESC_0_XUSER_9_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h38
`define WR_RESP_DESC_0_XUSER_10_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h3C
`define WR_RESP_DESC_0_XUSER_11_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h40
`define WR_RESP_DESC_0_XUSER_12_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h44
`define WR_RESP_DESC_0_XUSER_13_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h48
`define WR_RESP_DESC_0_XUSER_14_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h4C
`define WR_RESP_DESC_0_XUSER_15_REG_ADDR `WR_RESP_DESC_0_BASE_ADDR + 'h50
`define SN_REQ_DESC_0_ATTR_REG_ADDR `SN_REQ_DESC_0_BASE_ADDR + 'h0
`define SN_REQ_DESC_0_ACADDR_0_REG_ADDR `SN_REQ_DESC_0_BASE_ADDR + 'h4
`define SN_REQ_DESC_0_ACADDR_1_REG_ADDR `SN_REQ_DESC_0_BASE_ADDR + 'h8
`define SN_REQ_DESC_0_ACADDR_2_REG_ADDR `SN_REQ_DESC_0_BASE_ADDR + 'hC
`define SN_REQ_DESC_0_ACADDR_3_REG_ADDR `SN_REQ_DESC_0_BASE_ADDR + 'h10
`define SN_RESP_DESC_0_RESP_REG_ADDR `SN_RESP_DESC_0_BASE_ADDR + 'h0


`define RD_REQ_DESC_1_TXN_TYPE_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h0
`define RD_REQ_DESC_1_SIZE_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h4
`define RD_REQ_DESC_1_AXSIZE_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h8
`define RD_REQ_DESC_1_ATTR_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'hC
`define RD_REQ_DESC_1_AXADDR_0_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h10
`define RD_REQ_DESC_1_AXADDR_1_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h14
`define RD_REQ_DESC_1_AXADDR_2_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h18
`define RD_REQ_DESC_1_AXADDR_3_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h1C
`define RD_REQ_DESC_1_AXID_0_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h20
`define RD_REQ_DESC_1_AXID_1_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h24
`define RD_REQ_DESC_1_AXID_2_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h28
`define RD_REQ_DESC_1_AXID_3_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h2C
`define RD_REQ_DESC_1_AXUSER_0_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h30
`define RD_REQ_DESC_1_AXUSER_1_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h34
`define RD_REQ_DESC_1_AXUSER_2_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h38
`define RD_REQ_DESC_1_AXUSER_3_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h3C
`define RD_REQ_DESC_1_AXUSER_4_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h40
`define RD_REQ_DESC_1_AXUSER_5_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h44
`define RD_REQ_DESC_1_AXUSER_6_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h48
`define RD_REQ_DESC_1_AXUSER_7_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h4C
`define RD_REQ_DESC_1_AXUSER_8_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h50
`define RD_REQ_DESC_1_AXUSER_9_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h54
`define RD_REQ_DESC_1_AXUSER_10_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h58
`define RD_REQ_DESC_1_AXUSER_11_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h5C
`define RD_REQ_DESC_1_AXUSER_12_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h60
`define RD_REQ_DESC_1_AXUSER_13_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h64
`define RD_REQ_DESC_1_AXUSER_14_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h68
`define RD_REQ_DESC_1_AXUSER_15_REG_ADDR `RD_REQ_DESC_1_BASE_ADDR + 'h6C
`define RD_RESP_DESC_1_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h0
`define RD_RESP_DESC_1_DATA_SIZE_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h4
`define RD_RESP_DESC_1_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h8
`define RD_RESP_DESC_1_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'hC
`define RD_RESP_DESC_1_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h10
`define RD_RESP_DESC_1_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h14
`define RD_RESP_DESC_1_RESP_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h18
`define RD_RESP_DESC_1_XID_0_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h1C
`define RD_RESP_DESC_1_XID_1_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h20
`define RD_RESP_DESC_1_XID_2_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h24
`define RD_RESP_DESC_1_XID_3_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h28
`define RD_RESP_DESC_1_XUSER_0_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h2C
`define RD_RESP_DESC_1_XUSER_1_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h30
`define RD_RESP_DESC_1_XUSER_2_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h34
`define RD_RESP_DESC_1_XUSER_3_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h38
`define RD_RESP_DESC_1_XUSER_4_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h3C
`define RD_RESP_DESC_1_XUSER_5_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h40
`define RD_RESP_DESC_1_XUSER_6_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h44
`define RD_RESP_DESC_1_XUSER_7_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h48
`define RD_RESP_DESC_1_XUSER_8_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h4C
`define RD_RESP_DESC_1_XUSER_9_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h50
`define RD_RESP_DESC_1_XUSER_10_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h54
`define RD_RESP_DESC_1_XUSER_11_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h58
`define RD_RESP_DESC_1_XUSER_12_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h5C
`define RD_RESP_DESC_1_XUSER_13_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h60
`define RD_RESP_DESC_1_XUSER_14_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h64
`define RD_RESP_DESC_1_XUSER_15_REG_ADDR `RD_RESP_DESC_1_BASE_ADDR + 'h68
`define WR_REQ_DESC_1_TXN_TYPE_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h0
`define WR_REQ_DESC_1_SIZE_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h4
`define WR_REQ_DESC_1_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h8
`define WR_REQ_DESC_1_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hC
`define WR_REQ_DESC_1_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h10
`define WR_REQ_DESC_1_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h14
`define WR_REQ_DESC_1_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h18
`define WR_REQ_DESC_1_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h1C
`define WR_REQ_DESC_1_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h20
`define WR_REQ_DESC_1_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h24
`define WR_REQ_DESC_1_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h28
`define WR_REQ_DESC_1_AXSIZE_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h2C
`define WR_REQ_DESC_1_ATTR_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h30
`define WR_REQ_DESC_1_AXADDR_0_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h34
`define WR_REQ_DESC_1_AXADDR_1_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h38
`define WR_REQ_DESC_1_AXADDR_2_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h3C
`define WR_REQ_DESC_1_AXADDR_3_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h40
`define WR_REQ_DESC_1_AXID_0_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h44
`define WR_REQ_DESC_1_AXID_1_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h48
`define WR_REQ_DESC_1_AXID_2_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h4C
`define WR_REQ_DESC_1_AXID_3_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h50
`define WR_REQ_DESC_1_AXUSER_0_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h54
`define WR_REQ_DESC_1_AXUSER_1_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h58
`define WR_REQ_DESC_1_AXUSER_2_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h5C
`define WR_REQ_DESC_1_AXUSER_3_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h60
`define WR_REQ_DESC_1_AXUSER_4_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h64
`define WR_REQ_DESC_1_AXUSER_5_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h68
`define WR_REQ_DESC_1_AXUSER_6_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h6C
`define WR_REQ_DESC_1_AXUSER_7_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h70
`define WR_REQ_DESC_1_AXUSER_8_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h74
`define WR_REQ_DESC_1_AXUSER_9_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h78
`define WR_REQ_DESC_1_AXUSER_10_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h7C
`define WR_REQ_DESC_1_AXUSER_11_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h80
`define WR_REQ_DESC_1_AXUSER_12_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h84
`define WR_REQ_DESC_1_AXUSER_13_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h88
`define WR_REQ_DESC_1_AXUSER_14_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h8C
`define WR_REQ_DESC_1_AXUSER_15_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h90
`define WR_REQ_DESC_1_WUSER_0_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h94
`define WR_REQ_DESC_1_WUSER_1_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h98
`define WR_REQ_DESC_1_WUSER_2_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'h9C
`define WR_REQ_DESC_1_WUSER_3_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hA0
`define WR_REQ_DESC_1_WUSER_4_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hA4
`define WR_REQ_DESC_1_WUSER_5_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hA8
`define WR_REQ_DESC_1_WUSER_6_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hAC
`define WR_REQ_DESC_1_WUSER_7_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hB0
`define WR_REQ_DESC_1_WUSER_8_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hB4
`define WR_REQ_DESC_1_WUSER_9_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hB8
`define WR_REQ_DESC_1_WUSER_10_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hBC
`define WR_REQ_DESC_1_WUSER_11_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hC0
`define WR_REQ_DESC_1_WUSER_12_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hC4
`define WR_REQ_DESC_1_WUSER_13_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hC8
`define WR_REQ_DESC_1_WUSER_14_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hCC
`define WR_REQ_DESC_1_WUSER_15_REG_ADDR `WR_REQ_DESC_1_BASE_ADDR + 'hD0
`define WR_RESP_DESC_1_RESP_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h0
`define WR_RESP_DESC_1_XID_0_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h4
`define WR_RESP_DESC_1_XID_1_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h8
`define WR_RESP_DESC_1_XID_2_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'hC
`define WR_RESP_DESC_1_XID_3_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h10
`define WR_RESP_DESC_1_XUSER_0_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h14
`define WR_RESP_DESC_1_XUSER_1_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h18
`define WR_RESP_DESC_1_XUSER_2_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h1C
`define WR_RESP_DESC_1_XUSER_3_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h20
`define WR_RESP_DESC_1_XUSER_4_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h24
`define WR_RESP_DESC_1_XUSER_5_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h28
`define WR_RESP_DESC_1_XUSER_6_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h2C
`define WR_RESP_DESC_1_XUSER_7_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h30
`define WR_RESP_DESC_1_XUSER_8_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h34
`define WR_RESP_DESC_1_XUSER_9_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h38
`define WR_RESP_DESC_1_XUSER_10_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h3C
`define WR_RESP_DESC_1_XUSER_11_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h40
`define WR_RESP_DESC_1_XUSER_12_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h44
`define WR_RESP_DESC_1_XUSER_13_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h48
`define WR_RESP_DESC_1_XUSER_14_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h4C
`define WR_RESP_DESC_1_XUSER_15_REG_ADDR `WR_RESP_DESC_1_BASE_ADDR + 'h50
`define SN_REQ_DESC_1_ATTR_REG_ADDR `SN_REQ_DESC_1_BASE_ADDR + 'h0
`define SN_REQ_DESC_1_ACADDR_0_REG_ADDR `SN_REQ_DESC_1_BASE_ADDR + 'h4
`define SN_REQ_DESC_1_ACADDR_1_REG_ADDR `SN_REQ_DESC_1_BASE_ADDR + 'h8
`define SN_REQ_DESC_1_ACADDR_2_REG_ADDR `SN_REQ_DESC_1_BASE_ADDR + 'hC
`define SN_REQ_DESC_1_ACADDR_3_REG_ADDR `SN_REQ_DESC_1_BASE_ADDR + 'h10
`define SN_RESP_DESC_1_RESP_REG_ADDR `SN_RESP_DESC_1_BASE_ADDR + 'h0


`define RD_REQ_DESC_2_TXN_TYPE_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h0
`define RD_REQ_DESC_2_SIZE_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h4
`define RD_REQ_DESC_2_AXSIZE_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h8
`define RD_REQ_DESC_2_ATTR_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'hC
`define RD_REQ_DESC_2_AXADDR_0_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h10
`define RD_REQ_DESC_2_AXADDR_1_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h14
`define RD_REQ_DESC_2_AXADDR_2_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h18
`define RD_REQ_DESC_2_AXADDR_3_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h1C
`define RD_REQ_DESC_2_AXID_0_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h20
`define RD_REQ_DESC_2_AXID_1_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h24
`define RD_REQ_DESC_2_AXID_2_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h28
`define RD_REQ_DESC_2_AXID_3_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h2C
`define RD_REQ_DESC_2_AXUSER_0_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h30
`define RD_REQ_DESC_2_AXUSER_1_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h34
`define RD_REQ_DESC_2_AXUSER_2_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h38
`define RD_REQ_DESC_2_AXUSER_3_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h3C
`define RD_REQ_DESC_2_AXUSER_4_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h40
`define RD_REQ_DESC_2_AXUSER_5_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h44
`define RD_REQ_DESC_2_AXUSER_6_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h48
`define RD_REQ_DESC_2_AXUSER_7_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h4C
`define RD_REQ_DESC_2_AXUSER_8_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h50
`define RD_REQ_DESC_2_AXUSER_9_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h54
`define RD_REQ_DESC_2_AXUSER_10_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h58
`define RD_REQ_DESC_2_AXUSER_11_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h5C
`define RD_REQ_DESC_2_AXUSER_12_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h60
`define RD_REQ_DESC_2_AXUSER_13_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h64
`define RD_REQ_DESC_2_AXUSER_14_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h68
`define RD_REQ_DESC_2_AXUSER_15_REG_ADDR `RD_REQ_DESC_2_BASE_ADDR + 'h6C
`define RD_RESP_DESC_2_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h0
`define RD_RESP_DESC_2_DATA_SIZE_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h4
`define RD_RESP_DESC_2_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h8
`define RD_RESP_DESC_2_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'hC
`define RD_RESP_DESC_2_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h10
`define RD_RESP_DESC_2_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h14
`define RD_RESP_DESC_2_RESP_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h18
`define RD_RESP_DESC_2_XID_0_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h1C
`define RD_RESP_DESC_2_XID_1_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h20
`define RD_RESP_DESC_2_XID_2_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h24
`define RD_RESP_DESC_2_XID_3_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h28
`define RD_RESP_DESC_2_XUSER_0_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h2C
`define RD_RESP_DESC_2_XUSER_1_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h30
`define RD_RESP_DESC_2_XUSER_2_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h34
`define RD_RESP_DESC_2_XUSER_3_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h38
`define RD_RESP_DESC_2_XUSER_4_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h3C
`define RD_RESP_DESC_2_XUSER_5_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h40
`define RD_RESP_DESC_2_XUSER_6_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h44
`define RD_RESP_DESC_2_XUSER_7_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h48
`define RD_RESP_DESC_2_XUSER_8_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h4C
`define RD_RESP_DESC_2_XUSER_9_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h50
`define RD_RESP_DESC_2_XUSER_10_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h54
`define RD_RESP_DESC_2_XUSER_11_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h58
`define RD_RESP_DESC_2_XUSER_12_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h5C
`define RD_RESP_DESC_2_XUSER_13_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h60
`define RD_RESP_DESC_2_XUSER_14_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h64
`define RD_RESP_DESC_2_XUSER_15_REG_ADDR `RD_RESP_DESC_2_BASE_ADDR + 'h68
`define WR_REQ_DESC_2_TXN_TYPE_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h0
`define WR_REQ_DESC_2_SIZE_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h4
`define WR_REQ_DESC_2_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h8
`define WR_REQ_DESC_2_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hC
`define WR_REQ_DESC_2_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h10
`define WR_REQ_DESC_2_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h14
`define WR_REQ_DESC_2_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h18
`define WR_REQ_DESC_2_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h1C
`define WR_REQ_DESC_2_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h20
`define WR_REQ_DESC_2_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h24
`define WR_REQ_DESC_2_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h28
`define WR_REQ_DESC_2_AXSIZE_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h2C
`define WR_REQ_DESC_2_ATTR_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h30
`define WR_REQ_DESC_2_AXADDR_0_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h34
`define WR_REQ_DESC_2_AXADDR_1_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h38
`define WR_REQ_DESC_2_AXADDR_2_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h3C
`define WR_REQ_DESC_2_AXADDR_3_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h40
`define WR_REQ_DESC_2_AXID_0_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h44
`define WR_REQ_DESC_2_AXID_1_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h48
`define WR_REQ_DESC_2_AXID_2_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h4C
`define WR_REQ_DESC_2_AXID_3_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h50
`define WR_REQ_DESC_2_AXUSER_0_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h54
`define WR_REQ_DESC_2_AXUSER_1_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h58
`define WR_REQ_DESC_2_AXUSER_2_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h5C
`define WR_REQ_DESC_2_AXUSER_3_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h60
`define WR_REQ_DESC_2_AXUSER_4_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h64
`define WR_REQ_DESC_2_AXUSER_5_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h68
`define WR_REQ_DESC_2_AXUSER_6_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h6C
`define WR_REQ_DESC_2_AXUSER_7_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h70
`define WR_REQ_DESC_2_AXUSER_8_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h74
`define WR_REQ_DESC_2_AXUSER_9_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h78
`define WR_REQ_DESC_2_AXUSER_10_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h7C
`define WR_REQ_DESC_2_AXUSER_11_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h80
`define WR_REQ_DESC_2_AXUSER_12_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h84
`define WR_REQ_DESC_2_AXUSER_13_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h88
`define WR_REQ_DESC_2_AXUSER_14_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h8C
`define WR_REQ_DESC_2_AXUSER_15_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h90
`define WR_REQ_DESC_2_WUSER_0_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h94
`define WR_REQ_DESC_2_WUSER_1_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h98
`define WR_REQ_DESC_2_WUSER_2_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'h9C
`define WR_REQ_DESC_2_WUSER_3_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hA0
`define WR_REQ_DESC_2_WUSER_4_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hA4
`define WR_REQ_DESC_2_WUSER_5_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hA8
`define WR_REQ_DESC_2_WUSER_6_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hAC
`define WR_REQ_DESC_2_WUSER_7_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hB0
`define WR_REQ_DESC_2_WUSER_8_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hB4
`define WR_REQ_DESC_2_WUSER_9_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hB8
`define WR_REQ_DESC_2_WUSER_10_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hBC
`define WR_REQ_DESC_2_WUSER_11_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hC0
`define WR_REQ_DESC_2_WUSER_12_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hC4
`define WR_REQ_DESC_2_WUSER_13_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hC8
`define WR_REQ_DESC_2_WUSER_14_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hCC
`define WR_REQ_DESC_2_WUSER_15_REG_ADDR `WR_REQ_DESC_2_BASE_ADDR + 'hD0
`define WR_RESP_DESC_2_RESP_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h0
`define WR_RESP_DESC_2_XID_0_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h4
`define WR_RESP_DESC_2_XID_1_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h8
`define WR_RESP_DESC_2_XID_2_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'hC
`define WR_RESP_DESC_2_XID_3_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h10
`define WR_RESP_DESC_2_XUSER_0_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h14
`define WR_RESP_DESC_2_XUSER_1_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h18
`define WR_RESP_DESC_2_XUSER_2_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h1C
`define WR_RESP_DESC_2_XUSER_3_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h20
`define WR_RESP_DESC_2_XUSER_4_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h24
`define WR_RESP_DESC_2_XUSER_5_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h28
`define WR_RESP_DESC_2_XUSER_6_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h2C
`define WR_RESP_DESC_2_XUSER_7_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h30
`define WR_RESP_DESC_2_XUSER_8_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h34
`define WR_RESP_DESC_2_XUSER_9_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h38
`define WR_RESP_DESC_2_XUSER_10_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h3C
`define WR_RESP_DESC_2_XUSER_11_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h40
`define WR_RESP_DESC_2_XUSER_12_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h44
`define WR_RESP_DESC_2_XUSER_13_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h48
`define WR_RESP_DESC_2_XUSER_14_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h4C
`define WR_RESP_DESC_2_XUSER_15_REG_ADDR `WR_RESP_DESC_2_BASE_ADDR + 'h50
`define SN_REQ_DESC_2_ATTR_REG_ADDR `SN_REQ_DESC_2_BASE_ADDR + 'h0
`define SN_REQ_DESC_2_ACADDR_0_REG_ADDR `SN_REQ_DESC_2_BASE_ADDR + 'h4
`define SN_REQ_DESC_2_ACADDR_1_REG_ADDR `SN_REQ_DESC_2_BASE_ADDR + 'h8
`define SN_REQ_DESC_2_ACADDR_2_REG_ADDR `SN_REQ_DESC_2_BASE_ADDR + 'hC
`define SN_REQ_DESC_2_ACADDR_3_REG_ADDR `SN_REQ_DESC_2_BASE_ADDR + 'h10
`define SN_RESP_DESC_2_RESP_REG_ADDR `SN_RESP_DESC_2_BASE_ADDR + 'h0


`define RD_REQ_DESC_3_TXN_TYPE_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h0
`define RD_REQ_DESC_3_SIZE_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h4
`define RD_REQ_DESC_3_AXSIZE_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h8
`define RD_REQ_DESC_3_ATTR_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'hC
`define RD_REQ_DESC_3_AXADDR_0_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h10
`define RD_REQ_DESC_3_AXADDR_1_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h14
`define RD_REQ_DESC_3_AXADDR_2_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h18
`define RD_REQ_DESC_3_AXADDR_3_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h1C
`define RD_REQ_DESC_3_AXID_0_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h20
`define RD_REQ_DESC_3_AXID_1_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h24
`define RD_REQ_DESC_3_AXID_2_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h28
`define RD_REQ_DESC_3_AXID_3_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h2C
`define RD_REQ_DESC_3_AXUSER_0_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h30
`define RD_REQ_DESC_3_AXUSER_1_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h34
`define RD_REQ_DESC_3_AXUSER_2_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h38
`define RD_REQ_DESC_3_AXUSER_3_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h3C
`define RD_REQ_DESC_3_AXUSER_4_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h40
`define RD_REQ_DESC_3_AXUSER_5_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h44
`define RD_REQ_DESC_3_AXUSER_6_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h48
`define RD_REQ_DESC_3_AXUSER_7_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h4C
`define RD_REQ_DESC_3_AXUSER_8_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h50
`define RD_REQ_DESC_3_AXUSER_9_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h54
`define RD_REQ_DESC_3_AXUSER_10_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h58
`define RD_REQ_DESC_3_AXUSER_11_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h5C
`define RD_REQ_DESC_3_AXUSER_12_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h60
`define RD_REQ_DESC_3_AXUSER_13_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h64
`define RD_REQ_DESC_3_AXUSER_14_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h68
`define RD_REQ_DESC_3_AXUSER_15_REG_ADDR `RD_REQ_DESC_3_BASE_ADDR + 'h6C
`define RD_RESP_DESC_3_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h0
`define RD_RESP_DESC_3_DATA_SIZE_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h4
`define RD_RESP_DESC_3_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h8
`define RD_RESP_DESC_3_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'hC
`define RD_RESP_DESC_3_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h10
`define RD_RESP_DESC_3_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h14
`define RD_RESP_DESC_3_RESP_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h18
`define RD_RESP_DESC_3_XID_0_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h1C
`define RD_RESP_DESC_3_XID_1_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h20
`define RD_RESP_DESC_3_XID_2_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h24
`define RD_RESP_DESC_3_XID_3_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h28
`define RD_RESP_DESC_3_XUSER_0_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h2C
`define RD_RESP_DESC_3_XUSER_1_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h30
`define RD_RESP_DESC_3_XUSER_2_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h34
`define RD_RESP_DESC_3_XUSER_3_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h38
`define RD_RESP_DESC_3_XUSER_4_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h3C
`define RD_RESP_DESC_3_XUSER_5_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h40
`define RD_RESP_DESC_3_XUSER_6_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h44
`define RD_RESP_DESC_3_XUSER_7_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h48
`define RD_RESP_DESC_3_XUSER_8_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h4C
`define RD_RESP_DESC_3_XUSER_9_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h50
`define RD_RESP_DESC_3_XUSER_10_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h54
`define RD_RESP_DESC_3_XUSER_11_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h58
`define RD_RESP_DESC_3_XUSER_12_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h5C
`define RD_RESP_DESC_3_XUSER_13_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h60
`define RD_RESP_DESC_3_XUSER_14_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h64
`define RD_RESP_DESC_3_XUSER_15_REG_ADDR `RD_RESP_DESC_3_BASE_ADDR + 'h68
`define WR_REQ_DESC_3_TXN_TYPE_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h0
`define WR_REQ_DESC_3_SIZE_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h4
`define WR_REQ_DESC_3_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h8
`define WR_REQ_DESC_3_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hC
`define WR_REQ_DESC_3_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h10
`define WR_REQ_DESC_3_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h14
`define WR_REQ_DESC_3_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h18
`define WR_REQ_DESC_3_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h1C
`define WR_REQ_DESC_3_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h20
`define WR_REQ_DESC_3_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h24
`define WR_REQ_DESC_3_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h28
`define WR_REQ_DESC_3_AXSIZE_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h2C
`define WR_REQ_DESC_3_ATTR_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h30
`define WR_REQ_DESC_3_AXADDR_0_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h34
`define WR_REQ_DESC_3_AXADDR_1_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h38
`define WR_REQ_DESC_3_AXADDR_2_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h3C
`define WR_REQ_DESC_3_AXADDR_3_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h40
`define WR_REQ_DESC_3_AXID_0_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h44
`define WR_REQ_DESC_3_AXID_1_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h48
`define WR_REQ_DESC_3_AXID_2_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h4C
`define WR_REQ_DESC_3_AXID_3_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h50
`define WR_REQ_DESC_3_AXUSER_0_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h54
`define WR_REQ_DESC_3_AXUSER_1_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h58
`define WR_REQ_DESC_3_AXUSER_2_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h5C
`define WR_REQ_DESC_3_AXUSER_3_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h60
`define WR_REQ_DESC_3_AXUSER_4_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h64
`define WR_REQ_DESC_3_AXUSER_5_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h68
`define WR_REQ_DESC_3_AXUSER_6_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h6C
`define WR_REQ_DESC_3_AXUSER_7_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h70
`define WR_REQ_DESC_3_AXUSER_8_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h74
`define WR_REQ_DESC_3_AXUSER_9_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h78
`define WR_REQ_DESC_3_AXUSER_10_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h7C
`define WR_REQ_DESC_3_AXUSER_11_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h80
`define WR_REQ_DESC_3_AXUSER_12_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h84
`define WR_REQ_DESC_3_AXUSER_13_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h88
`define WR_REQ_DESC_3_AXUSER_14_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h8C
`define WR_REQ_DESC_3_AXUSER_15_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h90
`define WR_REQ_DESC_3_WUSER_0_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h94
`define WR_REQ_DESC_3_WUSER_1_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h98
`define WR_REQ_DESC_3_WUSER_2_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'h9C
`define WR_REQ_DESC_3_WUSER_3_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hA0
`define WR_REQ_DESC_3_WUSER_4_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hA4
`define WR_REQ_DESC_3_WUSER_5_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hA8
`define WR_REQ_DESC_3_WUSER_6_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hAC
`define WR_REQ_DESC_3_WUSER_7_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hB0
`define WR_REQ_DESC_3_WUSER_8_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hB4
`define WR_REQ_DESC_3_WUSER_9_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hB8
`define WR_REQ_DESC_3_WUSER_10_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hBC
`define WR_REQ_DESC_3_WUSER_11_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hC0
`define WR_REQ_DESC_3_WUSER_12_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hC4
`define WR_REQ_DESC_3_WUSER_13_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hC8
`define WR_REQ_DESC_3_WUSER_14_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hCC
`define WR_REQ_DESC_3_WUSER_15_REG_ADDR `WR_REQ_DESC_3_BASE_ADDR + 'hD0
`define WR_RESP_DESC_3_RESP_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h0
`define WR_RESP_DESC_3_XID_0_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h4
`define WR_RESP_DESC_3_XID_1_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h8
`define WR_RESP_DESC_3_XID_2_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'hC
`define WR_RESP_DESC_3_XID_3_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h10
`define WR_RESP_DESC_3_XUSER_0_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h14
`define WR_RESP_DESC_3_XUSER_1_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h18
`define WR_RESP_DESC_3_XUSER_2_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h1C
`define WR_RESP_DESC_3_XUSER_3_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h20
`define WR_RESP_DESC_3_XUSER_4_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h24
`define WR_RESP_DESC_3_XUSER_5_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h28
`define WR_RESP_DESC_3_XUSER_6_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h2C
`define WR_RESP_DESC_3_XUSER_7_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h30
`define WR_RESP_DESC_3_XUSER_8_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h34
`define WR_RESP_DESC_3_XUSER_9_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h38
`define WR_RESP_DESC_3_XUSER_10_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h3C
`define WR_RESP_DESC_3_XUSER_11_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h40
`define WR_RESP_DESC_3_XUSER_12_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h44
`define WR_RESP_DESC_3_XUSER_13_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h48
`define WR_RESP_DESC_3_XUSER_14_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h4C
`define WR_RESP_DESC_3_XUSER_15_REG_ADDR `WR_RESP_DESC_3_BASE_ADDR + 'h50
`define SN_REQ_DESC_3_ATTR_REG_ADDR `SN_REQ_DESC_3_BASE_ADDR + 'h0
`define SN_REQ_DESC_3_ACADDR_0_REG_ADDR `SN_REQ_DESC_3_BASE_ADDR + 'h4
`define SN_REQ_DESC_3_ACADDR_1_REG_ADDR `SN_REQ_DESC_3_BASE_ADDR + 'h8
`define SN_REQ_DESC_3_ACADDR_2_REG_ADDR `SN_REQ_DESC_3_BASE_ADDR + 'hC
`define SN_REQ_DESC_3_ACADDR_3_REG_ADDR `SN_REQ_DESC_3_BASE_ADDR + 'h10
`define SN_RESP_DESC_3_RESP_REG_ADDR `SN_RESP_DESC_3_BASE_ADDR + 'h0


`define RD_REQ_DESC_4_TXN_TYPE_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h0
`define RD_REQ_DESC_4_SIZE_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h4
`define RD_REQ_DESC_4_AXSIZE_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h8
`define RD_REQ_DESC_4_ATTR_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'hC
`define RD_REQ_DESC_4_AXADDR_0_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h10
`define RD_REQ_DESC_4_AXADDR_1_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h14
`define RD_REQ_DESC_4_AXADDR_2_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h18
`define RD_REQ_DESC_4_AXADDR_3_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h1C
`define RD_REQ_DESC_4_AXID_0_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h20
`define RD_REQ_DESC_4_AXID_1_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h24
`define RD_REQ_DESC_4_AXID_2_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h28
`define RD_REQ_DESC_4_AXID_3_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h2C
`define RD_REQ_DESC_4_AXUSER_0_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h30
`define RD_REQ_DESC_4_AXUSER_1_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h34
`define RD_REQ_DESC_4_AXUSER_2_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h38
`define RD_REQ_DESC_4_AXUSER_3_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h3C
`define RD_REQ_DESC_4_AXUSER_4_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h40
`define RD_REQ_DESC_4_AXUSER_5_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h44
`define RD_REQ_DESC_4_AXUSER_6_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h48
`define RD_REQ_DESC_4_AXUSER_7_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h4C
`define RD_REQ_DESC_4_AXUSER_8_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h50
`define RD_REQ_DESC_4_AXUSER_9_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h54
`define RD_REQ_DESC_4_AXUSER_10_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h58
`define RD_REQ_DESC_4_AXUSER_11_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h5C
`define RD_REQ_DESC_4_AXUSER_12_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h60
`define RD_REQ_DESC_4_AXUSER_13_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h64
`define RD_REQ_DESC_4_AXUSER_14_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h68
`define RD_REQ_DESC_4_AXUSER_15_REG_ADDR `RD_REQ_DESC_4_BASE_ADDR + 'h6C
`define RD_RESP_DESC_4_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h0
`define RD_RESP_DESC_4_DATA_SIZE_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h4
`define RD_RESP_DESC_4_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h8
`define RD_RESP_DESC_4_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'hC
`define RD_RESP_DESC_4_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h10
`define RD_RESP_DESC_4_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h14
`define RD_RESP_DESC_4_RESP_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h18
`define RD_RESP_DESC_4_XID_0_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h1C
`define RD_RESP_DESC_4_XID_1_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h20
`define RD_RESP_DESC_4_XID_2_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h24
`define RD_RESP_DESC_4_XID_3_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h28
`define RD_RESP_DESC_4_XUSER_0_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h2C
`define RD_RESP_DESC_4_XUSER_1_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h30
`define RD_RESP_DESC_4_XUSER_2_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h34
`define RD_RESP_DESC_4_XUSER_3_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h38
`define RD_RESP_DESC_4_XUSER_4_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h3C
`define RD_RESP_DESC_4_XUSER_5_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h40
`define RD_RESP_DESC_4_XUSER_6_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h44
`define RD_RESP_DESC_4_XUSER_7_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h48
`define RD_RESP_DESC_4_XUSER_8_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h4C
`define RD_RESP_DESC_4_XUSER_9_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h50
`define RD_RESP_DESC_4_XUSER_10_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h54
`define RD_RESP_DESC_4_XUSER_11_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h58
`define RD_RESP_DESC_4_XUSER_12_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h5C
`define RD_RESP_DESC_4_XUSER_13_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h60
`define RD_RESP_DESC_4_XUSER_14_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h64
`define RD_RESP_DESC_4_XUSER_15_REG_ADDR `RD_RESP_DESC_4_BASE_ADDR + 'h68
`define WR_REQ_DESC_4_TXN_TYPE_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h0
`define WR_REQ_DESC_4_SIZE_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h4
`define WR_REQ_DESC_4_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h8
`define WR_REQ_DESC_4_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hC
`define WR_REQ_DESC_4_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h10
`define WR_REQ_DESC_4_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h14
`define WR_REQ_DESC_4_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h18
`define WR_REQ_DESC_4_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h1C
`define WR_REQ_DESC_4_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h20
`define WR_REQ_DESC_4_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h24
`define WR_REQ_DESC_4_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h28
`define WR_REQ_DESC_4_AXSIZE_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h2C
`define WR_REQ_DESC_4_ATTR_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h30
`define WR_REQ_DESC_4_AXADDR_0_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h34
`define WR_REQ_DESC_4_AXADDR_1_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h38
`define WR_REQ_DESC_4_AXADDR_2_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h3C
`define WR_REQ_DESC_4_AXADDR_3_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h40
`define WR_REQ_DESC_4_AXID_0_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h44
`define WR_REQ_DESC_4_AXID_1_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h48
`define WR_REQ_DESC_4_AXID_2_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h4C
`define WR_REQ_DESC_4_AXID_3_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h50
`define WR_REQ_DESC_4_AXUSER_0_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h54
`define WR_REQ_DESC_4_AXUSER_1_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h58
`define WR_REQ_DESC_4_AXUSER_2_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h5C
`define WR_REQ_DESC_4_AXUSER_3_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h60
`define WR_REQ_DESC_4_AXUSER_4_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h64
`define WR_REQ_DESC_4_AXUSER_5_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h68
`define WR_REQ_DESC_4_AXUSER_6_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h6C
`define WR_REQ_DESC_4_AXUSER_7_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h70
`define WR_REQ_DESC_4_AXUSER_8_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h74
`define WR_REQ_DESC_4_AXUSER_9_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h78
`define WR_REQ_DESC_4_AXUSER_10_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h7C
`define WR_REQ_DESC_4_AXUSER_11_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h80
`define WR_REQ_DESC_4_AXUSER_12_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h84
`define WR_REQ_DESC_4_AXUSER_13_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h88
`define WR_REQ_DESC_4_AXUSER_14_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h8C
`define WR_REQ_DESC_4_AXUSER_15_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h90
`define WR_REQ_DESC_4_WUSER_0_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h94
`define WR_REQ_DESC_4_WUSER_1_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h98
`define WR_REQ_DESC_4_WUSER_2_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'h9C
`define WR_REQ_DESC_4_WUSER_3_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hA0
`define WR_REQ_DESC_4_WUSER_4_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hA4
`define WR_REQ_DESC_4_WUSER_5_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hA8
`define WR_REQ_DESC_4_WUSER_6_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hAC
`define WR_REQ_DESC_4_WUSER_7_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hB0
`define WR_REQ_DESC_4_WUSER_8_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hB4
`define WR_REQ_DESC_4_WUSER_9_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hB8
`define WR_REQ_DESC_4_WUSER_10_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hBC
`define WR_REQ_DESC_4_WUSER_11_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hC0
`define WR_REQ_DESC_4_WUSER_12_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hC4
`define WR_REQ_DESC_4_WUSER_13_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hC8
`define WR_REQ_DESC_4_WUSER_14_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hCC
`define WR_REQ_DESC_4_WUSER_15_REG_ADDR `WR_REQ_DESC_4_BASE_ADDR + 'hD0
`define WR_RESP_DESC_4_RESP_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h0
`define WR_RESP_DESC_4_XID_0_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h4
`define WR_RESP_DESC_4_XID_1_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h8
`define WR_RESP_DESC_4_XID_2_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'hC
`define WR_RESP_DESC_4_XID_3_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h10
`define WR_RESP_DESC_4_XUSER_0_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h14
`define WR_RESP_DESC_4_XUSER_1_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h18
`define WR_RESP_DESC_4_XUSER_2_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h1C
`define WR_RESP_DESC_4_XUSER_3_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h20
`define WR_RESP_DESC_4_XUSER_4_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h24
`define WR_RESP_DESC_4_XUSER_5_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h28
`define WR_RESP_DESC_4_XUSER_6_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h2C
`define WR_RESP_DESC_4_XUSER_7_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h30
`define WR_RESP_DESC_4_XUSER_8_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h34
`define WR_RESP_DESC_4_XUSER_9_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h38
`define WR_RESP_DESC_4_XUSER_10_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h3C
`define WR_RESP_DESC_4_XUSER_11_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h40
`define WR_RESP_DESC_4_XUSER_12_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h44
`define WR_RESP_DESC_4_XUSER_13_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h48
`define WR_RESP_DESC_4_XUSER_14_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h4C
`define WR_RESP_DESC_4_XUSER_15_REG_ADDR `WR_RESP_DESC_4_BASE_ADDR + 'h50
`define SN_REQ_DESC_4_ATTR_REG_ADDR `SN_REQ_DESC_4_BASE_ADDR + 'h0
`define SN_REQ_DESC_4_ACADDR_0_REG_ADDR `SN_REQ_DESC_4_BASE_ADDR + 'h4
`define SN_REQ_DESC_4_ACADDR_1_REG_ADDR `SN_REQ_DESC_4_BASE_ADDR + 'h8
`define SN_REQ_DESC_4_ACADDR_2_REG_ADDR `SN_REQ_DESC_4_BASE_ADDR + 'hC
`define SN_REQ_DESC_4_ACADDR_3_REG_ADDR `SN_REQ_DESC_4_BASE_ADDR + 'h10
`define SN_RESP_DESC_4_RESP_REG_ADDR `SN_RESP_DESC_4_BASE_ADDR + 'h0


`define RD_REQ_DESC_5_TXN_TYPE_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h0
`define RD_REQ_DESC_5_SIZE_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h4
`define RD_REQ_DESC_5_AXSIZE_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h8
`define RD_REQ_DESC_5_ATTR_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'hC
`define RD_REQ_DESC_5_AXADDR_0_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h10
`define RD_REQ_DESC_5_AXADDR_1_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h14
`define RD_REQ_DESC_5_AXADDR_2_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h18
`define RD_REQ_DESC_5_AXADDR_3_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h1C
`define RD_REQ_DESC_5_AXID_0_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h20
`define RD_REQ_DESC_5_AXID_1_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h24
`define RD_REQ_DESC_5_AXID_2_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h28
`define RD_REQ_DESC_5_AXID_3_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h2C
`define RD_REQ_DESC_5_AXUSER_0_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h30
`define RD_REQ_DESC_5_AXUSER_1_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h34
`define RD_REQ_DESC_5_AXUSER_2_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h38
`define RD_REQ_DESC_5_AXUSER_3_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h3C
`define RD_REQ_DESC_5_AXUSER_4_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h40
`define RD_REQ_DESC_5_AXUSER_5_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h44
`define RD_REQ_DESC_5_AXUSER_6_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h48
`define RD_REQ_DESC_5_AXUSER_7_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h4C
`define RD_REQ_DESC_5_AXUSER_8_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h50
`define RD_REQ_DESC_5_AXUSER_9_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h54
`define RD_REQ_DESC_5_AXUSER_10_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h58
`define RD_REQ_DESC_5_AXUSER_11_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h5C
`define RD_REQ_DESC_5_AXUSER_12_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h60
`define RD_REQ_DESC_5_AXUSER_13_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h64
`define RD_REQ_DESC_5_AXUSER_14_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h68
`define RD_REQ_DESC_5_AXUSER_15_REG_ADDR `RD_REQ_DESC_5_BASE_ADDR + 'h6C
`define RD_RESP_DESC_5_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h0
`define RD_RESP_DESC_5_DATA_SIZE_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h4
`define RD_RESP_DESC_5_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h8
`define RD_RESP_DESC_5_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'hC
`define RD_RESP_DESC_5_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h10
`define RD_RESP_DESC_5_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h14
`define RD_RESP_DESC_5_RESP_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h18
`define RD_RESP_DESC_5_XID_0_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h1C
`define RD_RESP_DESC_5_XID_1_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h20
`define RD_RESP_DESC_5_XID_2_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h24
`define RD_RESP_DESC_5_XID_3_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h28
`define RD_RESP_DESC_5_XUSER_0_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h2C
`define RD_RESP_DESC_5_XUSER_1_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h30
`define RD_RESP_DESC_5_XUSER_2_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h34
`define RD_RESP_DESC_5_XUSER_3_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h38
`define RD_RESP_DESC_5_XUSER_4_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h3C
`define RD_RESP_DESC_5_XUSER_5_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h40
`define RD_RESP_DESC_5_XUSER_6_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h44
`define RD_RESP_DESC_5_XUSER_7_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h48
`define RD_RESP_DESC_5_XUSER_8_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h4C
`define RD_RESP_DESC_5_XUSER_9_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h50
`define RD_RESP_DESC_5_XUSER_10_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h54
`define RD_RESP_DESC_5_XUSER_11_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h58
`define RD_RESP_DESC_5_XUSER_12_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h5C
`define RD_RESP_DESC_5_XUSER_13_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h60
`define RD_RESP_DESC_5_XUSER_14_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h64
`define RD_RESP_DESC_5_XUSER_15_REG_ADDR `RD_RESP_DESC_5_BASE_ADDR + 'h68
`define WR_REQ_DESC_5_TXN_TYPE_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h0
`define WR_REQ_DESC_5_SIZE_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h4
`define WR_REQ_DESC_5_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h8
`define WR_REQ_DESC_5_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hC
`define WR_REQ_DESC_5_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h10
`define WR_REQ_DESC_5_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h14
`define WR_REQ_DESC_5_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h18
`define WR_REQ_DESC_5_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h1C
`define WR_REQ_DESC_5_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h20
`define WR_REQ_DESC_5_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h24
`define WR_REQ_DESC_5_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h28
`define WR_REQ_DESC_5_AXSIZE_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h2C
`define WR_REQ_DESC_5_ATTR_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h30
`define WR_REQ_DESC_5_AXADDR_0_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h34
`define WR_REQ_DESC_5_AXADDR_1_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h38
`define WR_REQ_DESC_5_AXADDR_2_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h3C
`define WR_REQ_DESC_5_AXADDR_3_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h40
`define WR_REQ_DESC_5_AXID_0_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h44
`define WR_REQ_DESC_5_AXID_1_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h48
`define WR_REQ_DESC_5_AXID_2_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h4C
`define WR_REQ_DESC_5_AXID_3_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h50
`define WR_REQ_DESC_5_AXUSER_0_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h54
`define WR_REQ_DESC_5_AXUSER_1_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h58
`define WR_REQ_DESC_5_AXUSER_2_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h5C
`define WR_REQ_DESC_5_AXUSER_3_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h60
`define WR_REQ_DESC_5_AXUSER_4_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h64
`define WR_REQ_DESC_5_AXUSER_5_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h68
`define WR_REQ_DESC_5_AXUSER_6_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h6C
`define WR_REQ_DESC_5_AXUSER_7_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h70
`define WR_REQ_DESC_5_AXUSER_8_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h74
`define WR_REQ_DESC_5_AXUSER_9_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h78
`define WR_REQ_DESC_5_AXUSER_10_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h7C
`define WR_REQ_DESC_5_AXUSER_11_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h80
`define WR_REQ_DESC_5_AXUSER_12_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h84
`define WR_REQ_DESC_5_AXUSER_13_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h88
`define WR_REQ_DESC_5_AXUSER_14_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h8C
`define WR_REQ_DESC_5_AXUSER_15_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h90
`define WR_REQ_DESC_5_WUSER_0_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h94
`define WR_REQ_DESC_5_WUSER_1_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h98
`define WR_REQ_DESC_5_WUSER_2_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'h9C
`define WR_REQ_DESC_5_WUSER_3_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hA0
`define WR_REQ_DESC_5_WUSER_4_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hA4
`define WR_REQ_DESC_5_WUSER_5_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hA8
`define WR_REQ_DESC_5_WUSER_6_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hAC
`define WR_REQ_DESC_5_WUSER_7_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hB0
`define WR_REQ_DESC_5_WUSER_8_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hB4
`define WR_REQ_DESC_5_WUSER_9_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hB8
`define WR_REQ_DESC_5_WUSER_10_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hBC
`define WR_REQ_DESC_5_WUSER_11_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hC0
`define WR_REQ_DESC_5_WUSER_12_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hC4
`define WR_REQ_DESC_5_WUSER_13_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hC8
`define WR_REQ_DESC_5_WUSER_14_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hCC
`define WR_REQ_DESC_5_WUSER_15_REG_ADDR `WR_REQ_DESC_5_BASE_ADDR + 'hD0
`define WR_RESP_DESC_5_RESP_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h0
`define WR_RESP_DESC_5_XID_0_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h4
`define WR_RESP_DESC_5_XID_1_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h8
`define WR_RESP_DESC_5_XID_2_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'hC
`define WR_RESP_DESC_5_XID_3_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h10
`define WR_RESP_DESC_5_XUSER_0_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h14
`define WR_RESP_DESC_5_XUSER_1_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h18
`define WR_RESP_DESC_5_XUSER_2_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h1C
`define WR_RESP_DESC_5_XUSER_3_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h20
`define WR_RESP_DESC_5_XUSER_4_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h24
`define WR_RESP_DESC_5_XUSER_5_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h28
`define WR_RESP_DESC_5_XUSER_6_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h2C
`define WR_RESP_DESC_5_XUSER_7_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h30
`define WR_RESP_DESC_5_XUSER_8_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h34
`define WR_RESP_DESC_5_XUSER_9_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h38
`define WR_RESP_DESC_5_XUSER_10_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h3C
`define WR_RESP_DESC_5_XUSER_11_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h40
`define WR_RESP_DESC_5_XUSER_12_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h44
`define WR_RESP_DESC_5_XUSER_13_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h48
`define WR_RESP_DESC_5_XUSER_14_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h4C
`define WR_RESP_DESC_5_XUSER_15_REG_ADDR `WR_RESP_DESC_5_BASE_ADDR + 'h50
`define SN_REQ_DESC_5_ATTR_REG_ADDR `SN_REQ_DESC_5_BASE_ADDR + 'h0
`define SN_REQ_DESC_5_ACADDR_0_REG_ADDR `SN_REQ_DESC_5_BASE_ADDR + 'h4
`define SN_REQ_DESC_5_ACADDR_1_REG_ADDR `SN_REQ_DESC_5_BASE_ADDR + 'h8
`define SN_REQ_DESC_5_ACADDR_2_REG_ADDR `SN_REQ_DESC_5_BASE_ADDR + 'hC
`define SN_REQ_DESC_5_ACADDR_3_REG_ADDR `SN_REQ_DESC_5_BASE_ADDR + 'h10
`define SN_RESP_DESC_5_RESP_REG_ADDR `SN_RESP_DESC_5_BASE_ADDR + 'h0


`define RD_REQ_DESC_6_TXN_TYPE_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h0
`define RD_REQ_DESC_6_SIZE_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h4
`define RD_REQ_DESC_6_AXSIZE_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h8
`define RD_REQ_DESC_6_ATTR_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'hC
`define RD_REQ_DESC_6_AXADDR_0_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h10
`define RD_REQ_DESC_6_AXADDR_1_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h14
`define RD_REQ_DESC_6_AXADDR_2_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h18
`define RD_REQ_DESC_6_AXADDR_3_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h1C
`define RD_REQ_DESC_6_AXID_0_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h20
`define RD_REQ_DESC_6_AXID_1_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h24
`define RD_REQ_DESC_6_AXID_2_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h28
`define RD_REQ_DESC_6_AXID_3_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h2C
`define RD_REQ_DESC_6_AXUSER_0_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h30
`define RD_REQ_DESC_6_AXUSER_1_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h34
`define RD_REQ_DESC_6_AXUSER_2_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h38
`define RD_REQ_DESC_6_AXUSER_3_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h3C
`define RD_REQ_DESC_6_AXUSER_4_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h40
`define RD_REQ_DESC_6_AXUSER_5_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h44
`define RD_REQ_DESC_6_AXUSER_6_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h48
`define RD_REQ_DESC_6_AXUSER_7_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h4C
`define RD_REQ_DESC_6_AXUSER_8_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h50
`define RD_REQ_DESC_6_AXUSER_9_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h54
`define RD_REQ_DESC_6_AXUSER_10_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h58
`define RD_REQ_DESC_6_AXUSER_11_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h5C
`define RD_REQ_DESC_6_AXUSER_12_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h60
`define RD_REQ_DESC_6_AXUSER_13_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h64
`define RD_REQ_DESC_6_AXUSER_14_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h68
`define RD_REQ_DESC_6_AXUSER_15_REG_ADDR `RD_REQ_DESC_6_BASE_ADDR + 'h6C
`define RD_RESP_DESC_6_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h0
`define RD_RESP_DESC_6_DATA_SIZE_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h4
`define RD_RESP_DESC_6_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h8
`define RD_RESP_DESC_6_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'hC
`define RD_RESP_DESC_6_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h10
`define RD_RESP_DESC_6_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h14
`define RD_RESP_DESC_6_RESP_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h18
`define RD_RESP_DESC_6_XID_0_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h1C
`define RD_RESP_DESC_6_XID_1_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h20
`define RD_RESP_DESC_6_XID_2_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h24
`define RD_RESP_DESC_6_XID_3_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h28
`define RD_RESP_DESC_6_XUSER_0_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h2C
`define RD_RESP_DESC_6_XUSER_1_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h30
`define RD_RESP_DESC_6_XUSER_2_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h34
`define RD_RESP_DESC_6_XUSER_3_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h38
`define RD_RESP_DESC_6_XUSER_4_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h3C
`define RD_RESP_DESC_6_XUSER_5_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h40
`define RD_RESP_DESC_6_XUSER_6_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h44
`define RD_RESP_DESC_6_XUSER_7_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h48
`define RD_RESP_DESC_6_XUSER_8_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h4C
`define RD_RESP_DESC_6_XUSER_9_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h50
`define RD_RESP_DESC_6_XUSER_10_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h54
`define RD_RESP_DESC_6_XUSER_11_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h58
`define RD_RESP_DESC_6_XUSER_12_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h5C
`define RD_RESP_DESC_6_XUSER_13_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h60
`define RD_RESP_DESC_6_XUSER_14_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h64
`define RD_RESP_DESC_6_XUSER_15_REG_ADDR `RD_RESP_DESC_6_BASE_ADDR + 'h68
`define WR_REQ_DESC_6_TXN_TYPE_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h0
`define WR_REQ_DESC_6_SIZE_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h4
`define WR_REQ_DESC_6_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h8
`define WR_REQ_DESC_6_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hC
`define WR_REQ_DESC_6_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h10
`define WR_REQ_DESC_6_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h14
`define WR_REQ_DESC_6_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h18
`define WR_REQ_DESC_6_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h1C
`define WR_REQ_DESC_6_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h20
`define WR_REQ_DESC_6_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h24
`define WR_REQ_DESC_6_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h28
`define WR_REQ_DESC_6_AXSIZE_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h2C
`define WR_REQ_DESC_6_ATTR_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h30
`define WR_REQ_DESC_6_AXADDR_0_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h34
`define WR_REQ_DESC_6_AXADDR_1_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h38
`define WR_REQ_DESC_6_AXADDR_2_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h3C
`define WR_REQ_DESC_6_AXADDR_3_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h40
`define WR_REQ_DESC_6_AXID_0_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h44
`define WR_REQ_DESC_6_AXID_1_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h48
`define WR_REQ_DESC_6_AXID_2_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h4C
`define WR_REQ_DESC_6_AXID_3_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h50
`define WR_REQ_DESC_6_AXUSER_0_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h54
`define WR_REQ_DESC_6_AXUSER_1_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h58
`define WR_REQ_DESC_6_AXUSER_2_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h5C
`define WR_REQ_DESC_6_AXUSER_3_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h60
`define WR_REQ_DESC_6_AXUSER_4_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h64
`define WR_REQ_DESC_6_AXUSER_5_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h68
`define WR_REQ_DESC_6_AXUSER_6_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h6C
`define WR_REQ_DESC_6_AXUSER_7_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h70
`define WR_REQ_DESC_6_AXUSER_8_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h74
`define WR_REQ_DESC_6_AXUSER_9_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h78
`define WR_REQ_DESC_6_AXUSER_10_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h7C
`define WR_REQ_DESC_6_AXUSER_11_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h80
`define WR_REQ_DESC_6_AXUSER_12_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h84
`define WR_REQ_DESC_6_AXUSER_13_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h88
`define WR_REQ_DESC_6_AXUSER_14_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h8C
`define WR_REQ_DESC_6_AXUSER_15_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h90
`define WR_REQ_DESC_6_WUSER_0_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h94
`define WR_REQ_DESC_6_WUSER_1_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h98
`define WR_REQ_DESC_6_WUSER_2_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'h9C
`define WR_REQ_DESC_6_WUSER_3_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hA0
`define WR_REQ_DESC_6_WUSER_4_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hA4
`define WR_REQ_DESC_6_WUSER_5_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hA8
`define WR_REQ_DESC_6_WUSER_6_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hAC
`define WR_REQ_DESC_6_WUSER_7_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hB0
`define WR_REQ_DESC_6_WUSER_8_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hB4
`define WR_REQ_DESC_6_WUSER_9_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hB8
`define WR_REQ_DESC_6_WUSER_10_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hBC
`define WR_REQ_DESC_6_WUSER_11_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hC0
`define WR_REQ_DESC_6_WUSER_12_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hC4
`define WR_REQ_DESC_6_WUSER_13_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hC8
`define WR_REQ_DESC_6_WUSER_14_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hCC
`define WR_REQ_DESC_6_WUSER_15_REG_ADDR `WR_REQ_DESC_6_BASE_ADDR + 'hD0
`define WR_RESP_DESC_6_RESP_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h0
`define WR_RESP_DESC_6_XID_0_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h4
`define WR_RESP_DESC_6_XID_1_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h8
`define WR_RESP_DESC_6_XID_2_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'hC
`define WR_RESP_DESC_6_XID_3_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h10
`define WR_RESP_DESC_6_XUSER_0_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h14
`define WR_RESP_DESC_6_XUSER_1_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h18
`define WR_RESP_DESC_6_XUSER_2_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h1C
`define WR_RESP_DESC_6_XUSER_3_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h20
`define WR_RESP_DESC_6_XUSER_4_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h24
`define WR_RESP_DESC_6_XUSER_5_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h28
`define WR_RESP_DESC_6_XUSER_6_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h2C
`define WR_RESP_DESC_6_XUSER_7_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h30
`define WR_RESP_DESC_6_XUSER_8_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h34
`define WR_RESP_DESC_6_XUSER_9_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h38
`define WR_RESP_DESC_6_XUSER_10_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h3C
`define WR_RESP_DESC_6_XUSER_11_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h40
`define WR_RESP_DESC_6_XUSER_12_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h44
`define WR_RESP_DESC_6_XUSER_13_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h48
`define WR_RESP_DESC_6_XUSER_14_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h4C
`define WR_RESP_DESC_6_XUSER_15_REG_ADDR `WR_RESP_DESC_6_BASE_ADDR + 'h50
`define SN_REQ_DESC_6_ATTR_REG_ADDR `SN_REQ_DESC_6_BASE_ADDR + 'h0
`define SN_REQ_DESC_6_ACADDR_0_REG_ADDR `SN_REQ_DESC_6_BASE_ADDR + 'h4
`define SN_REQ_DESC_6_ACADDR_1_REG_ADDR `SN_REQ_DESC_6_BASE_ADDR + 'h8
`define SN_REQ_DESC_6_ACADDR_2_REG_ADDR `SN_REQ_DESC_6_BASE_ADDR + 'hC
`define SN_REQ_DESC_6_ACADDR_3_REG_ADDR `SN_REQ_DESC_6_BASE_ADDR + 'h10
`define SN_RESP_DESC_6_RESP_REG_ADDR `SN_RESP_DESC_6_BASE_ADDR + 'h0


`define RD_REQ_DESC_7_TXN_TYPE_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h0
`define RD_REQ_DESC_7_SIZE_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h4
`define RD_REQ_DESC_7_AXSIZE_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h8
`define RD_REQ_DESC_7_ATTR_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'hC
`define RD_REQ_DESC_7_AXADDR_0_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h10
`define RD_REQ_DESC_7_AXADDR_1_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h14
`define RD_REQ_DESC_7_AXADDR_2_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h18
`define RD_REQ_DESC_7_AXADDR_3_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h1C
`define RD_REQ_DESC_7_AXID_0_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h20
`define RD_REQ_DESC_7_AXID_1_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h24
`define RD_REQ_DESC_7_AXID_2_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h28
`define RD_REQ_DESC_7_AXID_3_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h2C
`define RD_REQ_DESC_7_AXUSER_0_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h30
`define RD_REQ_DESC_7_AXUSER_1_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h34
`define RD_REQ_DESC_7_AXUSER_2_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h38
`define RD_REQ_DESC_7_AXUSER_3_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h3C
`define RD_REQ_DESC_7_AXUSER_4_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h40
`define RD_REQ_DESC_7_AXUSER_5_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h44
`define RD_REQ_DESC_7_AXUSER_6_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h48
`define RD_REQ_DESC_7_AXUSER_7_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h4C
`define RD_REQ_DESC_7_AXUSER_8_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h50
`define RD_REQ_DESC_7_AXUSER_9_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h54
`define RD_REQ_DESC_7_AXUSER_10_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h58
`define RD_REQ_DESC_7_AXUSER_11_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h5C
`define RD_REQ_DESC_7_AXUSER_12_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h60
`define RD_REQ_DESC_7_AXUSER_13_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h64
`define RD_REQ_DESC_7_AXUSER_14_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h68
`define RD_REQ_DESC_7_AXUSER_15_REG_ADDR `RD_REQ_DESC_7_BASE_ADDR + 'h6C
`define RD_RESP_DESC_7_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h0
`define RD_RESP_DESC_7_DATA_SIZE_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h4
`define RD_RESP_DESC_7_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h8
`define RD_RESP_DESC_7_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'hC
`define RD_RESP_DESC_7_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h10
`define RD_RESP_DESC_7_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h14
`define RD_RESP_DESC_7_RESP_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h18
`define RD_RESP_DESC_7_XID_0_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h1C
`define RD_RESP_DESC_7_XID_1_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h20
`define RD_RESP_DESC_7_XID_2_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h24
`define RD_RESP_DESC_7_XID_3_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h28
`define RD_RESP_DESC_7_XUSER_0_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h2C
`define RD_RESP_DESC_7_XUSER_1_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h30
`define RD_RESP_DESC_7_XUSER_2_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h34
`define RD_RESP_DESC_7_XUSER_3_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h38
`define RD_RESP_DESC_7_XUSER_4_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h3C
`define RD_RESP_DESC_7_XUSER_5_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h40
`define RD_RESP_DESC_7_XUSER_6_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h44
`define RD_RESP_DESC_7_XUSER_7_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h48
`define RD_RESP_DESC_7_XUSER_8_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h4C
`define RD_RESP_DESC_7_XUSER_9_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h50
`define RD_RESP_DESC_7_XUSER_10_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h54
`define RD_RESP_DESC_7_XUSER_11_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h58
`define RD_RESP_DESC_7_XUSER_12_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h5C
`define RD_RESP_DESC_7_XUSER_13_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h60
`define RD_RESP_DESC_7_XUSER_14_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h64
`define RD_RESP_DESC_7_XUSER_15_REG_ADDR `RD_RESP_DESC_7_BASE_ADDR + 'h68
`define WR_REQ_DESC_7_TXN_TYPE_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h0
`define WR_REQ_DESC_7_SIZE_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h4
`define WR_REQ_DESC_7_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h8
`define WR_REQ_DESC_7_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hC
`define WR_REQ_DESC_7_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h10
`define WR_REQ_DESC_7_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h14
`define WR_REQ_DESC_7_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h18
`define WR_REQ_DESC_7_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h1C
`define WR_REQ_DESC_7_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h20
`define WR_REQ_DESC_7_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h24
`define WR_REQ_DESC_7_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h28
`define WR_REQ_DESC_7_AXSIZE_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h2C
`define WR_REQ_DESC_7_ATTR_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h30
`define WR_REQ_DESC_7_AXADDR_0_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h34
`define WR_REQ_DESC_7_AXADDR_1_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h38
`define WR_REQ_DESC_7_AXADDR_2_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h3C
`define WR_REQ_DESC_7_AXADDR_3_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h40
`define WR_REQ_DESC_7_AXID_0_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h44
`define WR_REQ_DESC_7_AXID_1_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h48
`define WR_REQ_DESC_7_AXID_2_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h4C
`define WR_REQ_DESC_7_AXID_3_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h50
`define WR_REQ_DESC_7_AXUSER_0_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h54
`define WR_REQ_DESC_7_AXUSER_1_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h58
`define WR_REQ_DESC_7_AXUSER_2_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h5C
`define WR_REQ_DESC_7_AXUSER_3_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h60
`define WR_REQ_DESC_7_AXUSER_4_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h64
`define WR_REQ_DESC_7_AXUSER_5_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h68
`define WR_REQ_DESC_7_AXUSER_6_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h6C
`define WR_REQ_DESC_7_AXUSER_7_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h70
`define WR_REQ_DESC_7_AXUSER_8_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h74
`define WR_REQ_DESC_7_AXUSER_9_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h78
`define WR_REQ_DESC_7_AXUSER_10_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h7C
`define WR_REQ_DESC_7_AXUSER_11_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h80
`define WR_REQ_DESC_7_AXUSER_12_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h84
`define WR_REQ_DESC_7_AXUSER_13_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h88
`define WR_REQ_DESC_7_AXUSER_14_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h8C
`define WR_REQ_DESC_7_AXUSER_15_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h90
`define WR_REQ_DESC_7_WUSER_0_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h94
`define WR_REQ_DESC_7_WUSER_1_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h98
`define WR_REQ_DESC_7_WUSER_2_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'h9C
`define WR_REQ_DESC_7_WUSER_3_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hA0
`define WR_REQ_DESC_7_WUSER_4_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hA4
`define WR_REQ_DESC_7_WUSER_5_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hA8
`define WR_REQ_DESC_7_WUSER_6_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hAC
`define WR_REQ_DESC_7_WUSER_7_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hB0
`define WR_REQ_DESC_7_WUSER_8_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hB4
`define WR_REQ_DESC_7_WUSER_9_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hB8
`define WR_REQ_DESC_7_WUSER_10_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hBC
`define WR_REQ_DESC_7_WUSER_11_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hC0
`define WR_REQ_DESC_7_WUSER_12_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hC4
`define WR_REQ_DESC_7_WUSER_13_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hC8
`define WR_REQ_DESC_7_WUSER_14_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hCC
`define WR_REQ_DESC_7_WUSER_15_REG_ADDR `WR_REQ_DESC_7_BASE_ADDR + 'hD0
`define WR_RESP_DESC_7_RESP_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h0
`define WR_RESP_DESC_7_XID_0_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h4
`define WR_RESP_DESC_7_XID_1_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h8
`define WR_RESP_DESC_7_XID_2_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'hC
`define WR_RESP_DESC_7_XID_3_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h10
`define WR_RESP_DESC_7_XUSER_0_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h14
`define WR_RESP_DESC_7_XUSER_1_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h18
`define WR_RESP_DESC_7_XUSER_2_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h1C
`define WR_RESP_DESC_7_XUSER_3_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h20
`define WR_RESP_DESC_7_XUSER_4_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h24
`define WR_RESP_DESC_7_XUSER_5_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h28
`define WR_RESP_DESC_7_XUSER_6_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h2C
`define WR_RESP_DESC_7_XUSER_7_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h30
`define WR_RESP_DESC_7_XUSER_8_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h34
`define WR_RESP_DESC_7_XUSER_9_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h38
`define WR_RESP_DESC_7_XUSER_10_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h3C
`define WR_RESP_DESC_7_XUSER_11_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h40
`define WR_RESP_DESC_7_XUSER_12_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h44
`define WR_RESP_DESC_7_XUSER_13_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h48
`define WR_RESP_DESC_7_XUSER_14_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h4C
`define WR_RESP_DESC_7_XUSER_15_REG_ADDR `WR_RESP_DESC_7_BASE_ADDR + 'h50
`define SN_REQ_DESC_7_ATTR_REG_ADDR `SN_REQ_DESC_7_BASE_ADDR + 'h0
`define SN_REQ_DESC_7_ACADDR_0_REG_ADDR `SN_REQ_DESC_7_BASE_ADDR + 'h4
`define SN_REQ_DESC_7_ACADDR_1_REG_ADDR `SN_REQ_DESC_7_BASE_ADDR + 'h8
`define SN_REQ_DESC_7_ACADDR_2_REG_ADDR `SN_REQ_DESC_7_BASE_ADDR + 'hC
`define SN_REQ_DESC_7_ACADDR_3_REG_ADDR `SN_REQ_DESC_7_BASE_ADDR + 'h10
`define SN_RESP_DESC_7_RESP_REG_ADDR `SN_RESP_DESC_7_BASE_ADDR + 'h0


`define RD_REQ_DESC_8_TXN_TYPE_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h0
`define RD_REQ_DESC_8_SIZE_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h4
`define RD_REQ_DESC_8_AXSIZE_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h8
`define RD_REQ_DESC_8_ATTR_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'hC
`define RD_REQ_DESC_8_AXADDR_0_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h10
`define RD_REQ_DESC_8_AXADDR_1_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h14
`define RD_REQ_DESC_8_AXADDR_2_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h18
`define RD_REQ_DESC_8_AXADDR_3_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h1C
`define RD_REQ_DESC_8_AXID_0_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h20
`define RD_REQ_DESC_8_AXID_1_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h24
`define RD_REQ_DESC_8_AXID_2_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h28
`define RD_REQ_DESC_8_AXID_3_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h2C
`define RD_REQ_DESC_8_AXUSER_0_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h30
`define RD_REQ_DESC_8_AXUSER_1_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h34
`define RD_REQ_DESC_8_AXUSER_2_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h38
`define RD_REQ_DESC_8_AXUSER_3_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h3C
`define RD_REQ_DESC_8_AXUSER_4_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h40
`define RD_REQ_DESC_8_AXUSER_5_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h44
`define RD_REQ_DESC_8_AXUSER_6_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h48
`define RD_REQ_DESC_8_AXUSER_7_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h4C
`define RD_REQ_DESC_8_AXUSER_8_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h50
`define RD_REQ_DESC_8_AXUSER_9_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h54
`define RD_REQ_DESC_8_AXUSER_10_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h58
`define RD_REQ_DESC_8_AXUSER_11_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h5C
`define RD_REQ_DESC_8_AXUSER_12_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h60
`define RD_REQ_DESC_8_AXUSER_13_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h64
`define RD_REQ_DESC_8_AXUSER_14_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h68
`define RD_REQ_DESC_8_AXUSER_15_REG_ADDR `RD_REQ_DESC_8_BASE_ADDR + 'h6C
`define RD_RESP_DESC_8_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h0
`define RD_RESP_DESC_8_DATA_SIZE_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h4
`define RD_RESP_DESC_8_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h8
`define RD_RESP_DESC_8_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'hC
`define RD_RESP_DESC_8_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h10
`define RD_RESP_DESC_8_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h14
`define RD_RESP_DESC_8_RESP_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h18
`define RD_RESP_DESC_8_XID_0_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h1C
`define RD_RESP_DESC_8_XID_1_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h20
`define RD_RESP_DESC_8_XID_2_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h24
`define RD_RESP_DESC_8_XID_3_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h28
`define RD_RESP_DESC_8_XUSER_0_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h2C
`define RD_RESP_DESC_8_XUSER_1_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h30
`define RD_RESP_DESC_8_XUSER_2_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h34
`define RD_RESP_DESC_8_XUSER_3_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h38
`define RD_RESP_DESC_8_XUSER_4_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h3C
`define RD_RESP_DESC_8_XUSER_5_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h40
`define RD_RESP_DESC_8_XUSER_6_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h44
`define RD_RESP_DESC_8_XUSER_7_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h48
`define RD_RESP_DESC_8_XUSER_8_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h4C
`define RD_RESP_DESC_8_XUSER_9_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h50
`define RD_RESP_DESC_8_XUSER_10_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h54
`define RD_RESP_DESC_8_XUSER_11_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h58
`define RD_RESP_DESC_8_XUSER_12_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h5C
`define RD_RESP_DESC_8_XUSER_13_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h60
`define RD_RESP_DESC_8_XUSER_14_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h64
`define RD_RESP_DESC_8_XUSER_15_REG_ADDR `RD_RESP_DESC_8_BASE_ADDR + 'h68
`define WR_REQ_DESC_8_TXN_TYPE_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h0
`define WR_REQ_DESC_8_SIZE_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h4
`define WR_REQ_DESC_8_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h8
`define WR_REQ_DESC_8_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hC
`define WR_REQ_DESC_8_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h10
`define WR_REQ_DESC_8_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h14
`define WR_REQ_DESC_8_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h18
`define WR_REQ_DESC_8_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h1C
`define WR_REQ_DESC_8_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h20
`define WR_REQ_DESC_8_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h24
`define WR_REQ_DESC_8_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h28
`define WR_REQ_DESC_8_AXSIZE_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h2C
`define WR_REQ_DESC_8_ATTR_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h30
`define WR_REQ_DESC_8_AXADDR_0_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h34
`define WR_REQ_DESC_8_AXADDR_1_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h38
`define WR_REQ_DESC_8_AXADDR_2_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h3C
`define WR_REQ_DESC_8_AXADDR_3_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h40
`define WR_REQ_DESC_8_AXID_0_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h44
`define WR_REQ_DESC_8_AXID_1_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h48
`define WR_REQ_DESC_8_AXID_2_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h4C
`define WR_REQ_DESC_8_AXID_3_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h50
`define WR_REQ_DESC_8_AXUSER_0_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h54
`define WR_REQ_DESC_8_AXUSER_1_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h58
`define WR_REQ_DESC_8_AXUSER_2_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h5C
`define WR_REQ_DESC_8_AXUSER_3_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h60
`define WR_REQ_DESC_8_AXUSER_4_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h64
`define WR_REQ_DESC_8_AXUSER_5_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h68
`define WR_REQ_DESC_8_AXUSER_6_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h6C
`define WR_REQ_DESC_8_AXUSER_7_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h70
`define WR_REQ_DESC_8_AXUSER_8_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h74
`define WR_REQ_DESC_8_AXUSER_9_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h78
`define WR_REQ_DESC_8_AXUSER_10_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h7C
`define WR_REQ_DESC_8_AXUSER_11_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h80
`define WR_REQ_DESC_8_AXUSER_12_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h84
`define WR_REQ_DESC_8_AXUSER_13_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h88
`define WR_REQ_DESC_8_AXUSER_14_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h8C
`define WR_REQ_DESC_8_AXUSER_15_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h90
`define WR_REQ_DESC_8_WUSER_0_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h94
`define WR_REQ_DESC_8_WUSER_1_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h98
`define WR_REQ_DESC_8_WUSER_2_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'h9C
`define WR_REQ_DESC_8_WUSER_3_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hA0
`define WR_REQ_DESC_8_WUSER_4_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hA4
`define WR_REQ_DESC_8_WUSER_5_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hA8
`define WR_REQ_DESC_8_WUSER_6_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hAC
`define WR_REQ_DESC_8_WUSER_7_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hB0
`define WR_REQ_DESC_8_WUSER_8_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hB4
`define WR_REQ_DESC_8_WUSER_9_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hB8
`define WR_REQ_DESC_8_WUSER_10_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hBC
`define WR_REQ_DESC_8_WUSER_11_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hC0
`define WR_REQ_DESC_8_WUSER_12_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hC4
`define WR_REQ_DESC_8_WUSER_13_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hC8
`define WR_REQ_DESC_8_WUSER_14_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hCC
`define WR_REQ_DESC_8_WUSER_15_REG_ADDR `WR_REQ_DESC_8_BASE_ADDR + 'hD0
`define WR_RESP_DESC_8_RESP_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h0
`define WR_RESP_DESC_8_XID_0_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h4
`define WR_RESP_DESC_8_XID_1_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h8
`define WR_RESP_DESC_8_XID_2_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'hC
`define WR_RESP_DESC_8_XID_3_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h10
`define WR_RESP_DESC_8_XUSER_0_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h14
`define WR_RESP_DESC_8_XUSER_1_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h18
`define WR_RESP_DESC_8_XUSER_2_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h1C
`define WR_RESP_DESC_8_XUSER_3_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h20
`define WR_RESP_DESC_8_XUSER_4_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h24
`define WR_RESP_DESC_8_XUSER_5_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h28
`define WR_RESP_DESC_8_XUSER_6_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h2C
`define WR_RESP_DESC_8_XUSER_7_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h30
`define WR_RESP_DESC_8_XUSER_8_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h34
`define WR_RESP_DESC_8_XUSER_9_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h38
`define WR_RESP_DESC_8_XUSER_10_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h3C
`define WR_RESP_DESC_8_XUSER_11_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h40
`define WR_RESP_DESC_8_XUSER_12_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h44
`define WR_RESP_DESC_8_XUSER_13_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h48
`define WR_RESP_DESC_8_XUSER_14_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h4C
`define WR_RESP_DESC_8_XUSER_15_REG_ADDR `WR_RESP_DESC_8_BASE_ADDR + 'h50
`define SN_REQ_DESC_8_ATTR_REG_ADDR `SN_REQ_DESC_8_BASE_ADDR + 'h0
`define SN_REQ_DESC_8_ACADDR_0_REG_ADDR `SN_REQ_DESC_8_BASE_ADDR + 'h4
`define SN_REQ_DESC_8_ACADDR_1_REG_ADDR `SN_REQ_DESC_8_BASE_ADDR + 'h8
`define SN_REQ_DESC_8_ACADDR_2_REG_ADDR `SN_REQ_DESC_8_BASE_ADDR + 'hC
`define SN_REQ_DESC_8_ACADDR_3_REG_ADDR `SN_REQ_DESC_8_BASE_ADDR + 'h10
`define SN_RESP_DESC_8_RESP_REG_ADDR `SN_RESP_DESC_8_BASE_ADDR + 'h0


`define RD_REQ_DESC_9_TXN_TYPE_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h0
`define RD_REQ_DESC_9_SIZE_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h4
`define RD_REQ_DESC_9_AXSIZE_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h8
`define RD_REQ_DESC_9_ATTR_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'hC
`define RD_REQ_DESC_9_AXADDR_0_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h10
`define RD_REQ_DESC_9_AXADDR_1_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h14
`define RD_REQ_DESC_9_AXADDR_2_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h18
`define RD_REQ_DESC_9_AXADDR_3_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h1C
`define RD_REQ_DESC_9_AXID_0_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h20
`define RD_REQ_DESC_9_AXID_1_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h24
`define RD_REQ_DESC_9_AXID_2_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h28
`define RD_REQ_DESC_9_AXID_3_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h2C
`define RD_REQ_DESC_9_AXUSER_0_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h30
`define RD_REQ_DESC_9_AXUSER_1_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h34
`define RD_REQ_DESC_9_AXUSER_2_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h38
`define RD_REQ_DESC_9_AXUSER_3_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h3C
`define RD_REQ_DESC_9_AXUSER_4_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h40
`define RD_REQ_DESC_9_AXUSER_5_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h44
`define RD_REQ_DESC_9_AXUSER_6_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h48
`define RD_REQ_DESC_9_AXUSER_7_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h4C
`define RD_REQ_DESC_9_AXUSER_8_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h50
`define RD_REQ_DESC_9_AXUSER_9_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h54
`define RD_REQ_DESC_9_AXUSER_10_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h58
`define RD_REQ_DESC_9_AXUSER_11_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h5C
`define RD_REQ_DESC_9_AXUSER_12_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h60
`define RD_REQ_DESC_9_AXUSER_13_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h64
`define RD_REQ_DESC_9_AXUSER_14_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h68
`define RD_REQ_DESC_9_AXUSER_15_REG_ADDR `RD_REQ_DESC_9_BASE_ADDR + 'h6C
`define RD_RESP_DESC_9_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h0
`define RD_RESP_DESC_9_DATA_SIZE_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h4
`define RD_RESP_DESC_9_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h8
`define RD_RESP_DESC_9_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'hC
`define RD_RESP_DESC_9_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h10
`define RD_RESP_DESC_9_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h14
`define RD_RESP_DESC_9_RESP_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h18
`define RD_RESP_DESC_9_XID_0_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h1C
`define RD_RESP_DESC_9_XID_1_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h20
`define RD_RESP_DESC_9_XID_2_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h24
`define RD_RESP_DESC_9_XID_3_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h28
`define RD_RESP_DESC_9_XUSER_0_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h2C
`define RD_RESP_DESC_9_XUSER_1_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h30
`define RD_RESP_DESC_9_XUSER_2_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h34
`define RD_RESP_DESC_9_XUSER_3_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h38
`define RD_RESP_DESC_9_XUSER_4_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h3C
`define RD_RESP_DESC_9_XUSER_5_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h40
`define RD_RESP_DESC_9_XUSER_6_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h44
`define RD_RESP_DESC_9_XUSER_7_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h48
`define RD_RESP_DESC_9_XUSER_8_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h4C
`define RD_RESP_DESC_9_XUSER_9_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h50
`define RD_RESP_DESC_9_XUSER_10_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h54
`define RD_RESP_DESC_9_XUSER_11_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h58
`define RD_RESP_DESC_9_XUSER_12_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h5C
`define RD_RESP_DESC_9_XUSER_13_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h60
`define RD_RESP_DESC_9_XUSER_14_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h64
`define RD_RESP_DESC_9_XUSER_15_REG_ADDR `RD_RESP_DESC_9_BASE_ADDR + 'h68
`define WR_REQ_DESC_9_TXN_TYPE_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h0
`define WR_REQ_DESC_9_SIZE_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h4
`define WR_REQ_DESC_9_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h8
`define WR_REQ_DESC_9_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hC
`define WR_REQ_DESC_9_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h10
`define WR_REQ_DESC_9_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h14
`define WR_REQ_DESC_9_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h18
`define WR_REQ_DESC_9_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h1C
`define WR_REQ_DESC_9_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h20
`define WR_REQ_DESC_9_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h24
`define WR_REQ_DESC_9_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h28
`define WR_REQ_DESC_9_AXSIZE_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h2C
`define WR_REQ_DESC_9_ATTR_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h30
`define WR_REQ_DESC_9_AXADDR_0_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h34
`define WR_REQ_DESC_9_AXADDR_1_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h38
`define WR_REQ_DESC_9_AXADDR_2_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h3C
`define WR_REQ_DESC_9_AXADDR_3_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h40
`define WR_REQ_DESC_9_AXID_0_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h44
`define WR_REQ_DESC_9_AXID_1_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h48
`define WR_REQ_DESC_9_AXID_2_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h4C
`define WR_REQ_DESC_9_AXID_3_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h50
`define WR_REQ_DESC_9_AXUSER_0_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h54
`define WR_REQ_DESC_9_AXUSER_1_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h58
`define WR_REQ_DESC_9_AXUSER_2_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h5C
`define WR_REQ_DESC_9_AXUSER_3_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h60
`define WR_REQ_DESC_9_AXUSER_4_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h64
`define WR_REQ_DESC_9_AXUSER_5_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h68
`define WR_REQ_DESC_9_AXUSER_6_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h6C
`define WR_REQ_DESC_9_AXUSER_7_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h70
`define WR_REQ_DESC_9_AXUSER_8_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h74
`define WR_REQ_DESC_9_AXUSER_9_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h78
`define WR_REQ_DESC_9_AXUSER_10_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h7C
`define WR_REQ_DESC_9_AXUSER_11_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h80
`define WR_REQ_DESC_9_AXUSER_12_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h84
`define WR_REQ_DESC_9_AXUSER_13_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h88
`define WR_REQ_DESC_9_AXUSER_14_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h8C
`define WR_REQ_DESC_9_AXUSER_15_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h90
`define WR_REQ_DESC_9_WUSER_0_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h94
`define WR_REQ_DESC_9_WUSER_1_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h98
`define WR_REQ_DESC_9_WUSER_2_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'h9C
`define WR_REQ_DESC_9_WUSER_3_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hA0
`define WR_REQ_DESC_9_WUSER_4_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hA4
`define WR_REQ_DESC_9_WUSER_5_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hA8
`define WR_REQ_DESC_9_WUSER_6_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hAC
`define WR_REQ_DESC_9_WUSER_7_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hB0
`define WR_REQ_DESC_9_WUSER_8_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hB4
`define WR_REQ_DESC_9_WUSER_9_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hB8
`define WR_REQ_DESC_9_WUSER_10_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hBC
`define WR_REQ_DESC_9_WUSER_11_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hC0
`define WR_REQ_DESC_9_WUSER_12_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hC4
`define WR_REQ_DESC_9_WUSER_13_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hC8
`define WR_REQ_DESC_9_WUSER_14_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hCC
`define WR_REQ_DESC_9_WUSER_15_REG_ADDR `WR_REQ_DESC_9_BASE_ADDR + 'hD0
`define WR_RESP_DESC_9_RESP_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h0
`define WR_RESP_DESC_9_XID_0_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h4
`define WR_RESP_DESC_9_XID_1_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h8
`define WR_RESP_DESC_9_XID_2_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'hC
`define WR_RESP_DESC_9_XID_3_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h10
`define WR_RESP_DESC_9_XUSER_0_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h14
`define WR_RESP_DESC_9_XUSER_1_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h18
`define WR_RESP_DESC_9_XUSER_2_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h1C
`define WR_RESP_DESC_9_XUSER_3_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h20
`define WR_RESP_DESC_9_XUSER_4_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h24
`define WR_RESP_DESC_9_XUSER_5_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h28
`define WR_RESP_DESC_9_XUSER_6_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h2C
`define WR_RESP_DESC_9_XUSER_7_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h30
`define WR_RESP_DESC_9_XUSER_8_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h34
`define WR_RESP_DESC_9_XUSER_9_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h38
`define WR_RESP_DESC_9_XUSER_10_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h3C
`define WR_RESP_DESC_9_XUSER_11_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h40
`define WR_RESP_DESC_9_XUSER_12_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h44
`define WR_RESP_DESC_9_XUSER_13_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h48
`define WR_RESP_DESC_9_XUSER_14_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h4C
`define WR_RESP_DESC_9_XUSER_15_REG_ADDR `WR_RESP_DESC_9_BASE_ADDR + 'h50
`define SN_REQ_DESC_9_ATTR_REG_ADDR `SN_REQ_DESC_9_BASE_ADDR + 'h0
`define SN_REQ_DESC_9_ACADDR_0_REG_ADDR `SN_REQ_DESC_9_BASE_ADDR + 'h4
`define SN_REQ_DESC_9_ACADDR_1_REG_ADDR `SN_REQ_DESC_9_BASE_ADDR + 'h8
`define SN_REQ_DESC_9_ACADDR_2_REG_ADDR `SN_REQ_DESC_9_BASE_ADDR + 'hC
`define SN_REQ_DESC_9_ACADDR_3_REG_ADDR `SN_REQ_DESC_9_BASE_ADDR + 'h10
`define SN_RESP_DESC_9_RESP_REG_ADDR `SN_RESP_DESC_9_BASE_ADDR + 'h0


`define RD_REQ_DESC_A_TXN_TYPE_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h0
`define RD_REQ_DESC_A_SIZE_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h4
`define RD_REQ_DESC_A_AXSIZE_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h8
`define RD_REQ_DESC_A_ATTR_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'hC
`define RD_REQ_DESC_A_AXADDR_0_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h10
`define RD_REQ_DESC_A_AXADDR_1_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h14
`define RD_REQ_DESC_A_AXADDR_2_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h18
`define RD_REQ_DESC_A_AXADDR_3_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h1C
`define RD_REQ_DESC_A_AXID_0_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h20
`define RD_REQ_DESC_A_AXID_1_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h24
`define RD_REQ_DESC_A_AXID_2_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h28
`define RD_REQ_DESC_A_AXID_3_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h2C
`define RD_REQ_DESC_A_AXUSER_0_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h30
`define RD_REQ_DESC_A_AXUSER_1_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h34
`define RD_REQ_DESC_A_AXUSER_2_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h38
`define RD_REQ_DESC_A_AXUSER_3_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h3C
`define RD_REQ_DESC_A_AXUSER_4_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h40
`define RD_REQ_DESC_A_AXUSER_5_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h44
`define RD_REQ_DESC_A_AXUSER_6_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h48
`define RD_REQ_DESC_A_AXUSER_7_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h4C
`define RD_REQ_DESC_A_AXUSER_8_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h50
`define RD_REQ_DESC_A_AXUSER_9_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h54
`define RD_REQ_DESC_A_AXUSER_10_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h58
`define RD_REQ_DESC_A_AXUSER_11_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h5C
`define RD_REQ_DESC_A_AXUSER_12_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h60
`define RD_REQ_DESC_A_AXUSER_13_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h64
`define RD_REQ_DESC_A_AXUSER_14_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h68
`define RD_REQ_DESC_A_AXUSER_15_REG_ADDR `RD_REQ_DESC_A_BASE_ADDR + 'h6C
`define RD_RESP_DESC_A_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h0
`define RD_RESP_DESC_A_DATA_SIZE_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h4
`define RD_RESP_DESC_A_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h8
`define RD_RESP_DESC_A_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'hC
`define RD_RESP_DESC_A_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h10
`define RD_RESP_DESC_A_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h14
`define RD_RESP_DESC_A_RESP_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h18
`define RD_RESP_DESC_A_XID_0_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h1C
`define RD_RESP_DESC_A_XID_1_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h20
`define RD_RESP_DESC_A_XID_2_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h24
`define RD_RESP_DESC_A_XID_3_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h28
`define RD_RESP_DESC_A_XUSER_0_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h2C
`define RD_RESP_DESC_A_XUSER_1_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h30
`define RD_RESP_DESC_A_XUSER_2_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h34
`define RD_RESP_DESC_A_XUSER_3_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h38
`define RD_RESP_DESC_A_XUSER_4_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h3C
`define RD_RESP_DESC_A_XUSER_5_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h40
`define RD_RESP_DESC_A_XUSER_6_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h44
`define RD_RESP_DESC_A_XUSER_7_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h48
`define RD_RESP_DESC_A_XUSER_8_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h4C
`define RD_RESP_DESC_A_XUSER_9_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h50
`define RD_RESP_DESC_A_XUSER_10_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h54
`define RD_RESP_DESC_A_XUSER_11_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h58
`define RD_RESP_DESC_A_XUSER_12_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h5C
`define RD_RESP_DESC_A_XUSER_13_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h60
`define RD_RESP_DESC_A_XUSER_14_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h64
`define RD_RESP_DESC_A_XUSER_15_REG_ADDR `RD_RESP_DESC_A_BASE_ADDR + 'h68
`define WR_REQ_DESC_A_TXN_TYPE_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h0
`define WR_REQ_DESC_A_SIZE_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h4
`define WR_REQ_DESC_A_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h8
`define WR_REQ_DESC_A_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hC
`define WR_REQ_DESC_A_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h10
`define WR_REQ_DESC_A_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h14
`define WR_REQ_DESC_A_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h18
`define WR_REQ_DESC_A_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h1C
`define WR_REQ_DESC_A_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h20
`define WR_REQ_DESC_A_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h24
`define WR_REQ_DESC_A_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h28
`define WR_REQ_DESC_A_AXSIZE_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h2C
`define WR_REQ_DESC_A_ATTR_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h30
`define WR_REQ_DESC_A_AXADDR_0_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h34
`define WR_REQ_DESC_A_AXADDR_1_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h38
`define WR_REQ_DESC_A_AXADDR_2_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h3C
`define WR_REQ_DESC_A_AXADDR_3_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h40
`define WR_REQ_DESC_A_AXID_0_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h44
`define WR_REQ_DESC_A_AXID_1_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h48
`define WR_REQ_DESC_A_AXID_2_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h4C
`define WR_REQ_DESC_A_AXID_3_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h50
`define WR_REQ_DESC_A_AXUSER_0_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h54
`define WR_REQ_DESC_A_AXUSER_1_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h58
`define WR_REQ_DESC_A_AXUSER_2_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h5C
`define WR_REQ_DESC_A_AXUSER_3_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h60
`define WR_REQ_DESC_A_AXUSER_4_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h64
`define WR_REQ_DESC_A_AXUSER_5_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h68
`define WR_REQ_DESC_A_AXUSER_6_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h6C
`define WR_REQ_DESC_A_AXUSER_7_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h70
`define WR_REQ_DESC_A_AXUSER_8_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h74
`define WR_REQ_DESC_A_AXUSER_9_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h78
`define WR_REQ_DESC_A_AXUSER_10_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h7C
`define WR_REQ_DESC_A_AXUSER_11_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h80
`define WR_REQ_DESC_A_AXUSER_12_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h84
`define WR_REQ_DESC_A_AXUSER_13_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h88
`define WR_REQ_DESC_A_AXUSER_14_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h8C
`define WR_REQ_DESC_A_AXUSER_15_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h90
`define WR_REQ_DESC_A_WUSER_0_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h94
`define WR_REQ_DESC_A_WUSER_1_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h98
`define WR_REQ_DESC_A_WUSER_2_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'h9C
`define WR_REQ_DESC_A_WUSER_3_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hA0
`define WR_REQ_DESC_A_WUSER_4_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hA4
`define WR_REQ_DESC_A_WUSER_5_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hA8
`define WR_REQ_DESC_A_WUSER_6_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hAC
`define WR_REQ_DESC_A_WUSER_7_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hB0
`define WR_REQ_DESC_A_WUSER_8_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hB4
`define WR_REQ_DESC_A_WUSER_9_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hB8
`define WR_REQ_DESC_A_WUSER_10_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hBC
`define WR_REQ_DESC_A_WUSER_11_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hC0
`define WR_REQ_DESC_A_WUSER_12_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hC4
`define WR_REQ_DESC_A_WUSER_13_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hC8
`define WR_REQ_DESC_A_WUSER_14_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hCC
`define WR_REQ_DESC_A_WUSER_15_REG_ADDR `WR_REQ_DESC_A_BASE_ADDR + 'hD0
`define WR_RESP_DESC_A_RESP_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h0
`define WR_RESP_DESC_A_XID_0_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h4
`define WR_RESP_DESC_A_XID_1_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h8
`define WR_RESP_DESC_A_XID_2_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'hC
`define WR_RESP_DESC_A_XID_3_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h10
`define WR_RESP_DESC_A_XUSER_0_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h14
`define WR_RESP_DESC_A_XUSER_1_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h18
`define WR_RESP_DESC_A_XUSER_2_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h1C
`define WR_RESP_DESC_A_XUSER_3_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h20
`define WR_RESP_DESC_A_XUSER_4_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h24
`define WR_RESP_DESC_A_XUSER_5_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h28
`define WR_RESP_DESC_A_XUSER_6_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h2C
`define WR_RESP_DESC_A_XUSER_7_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h30
`define WR_RESP_DESC_A_XUSER_8_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h34
`define WR_RESP_DESC_A_XUSER_9_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h38
`define WR_RESP_DESC_A_XUSER_10_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h3C
`define WR_RESP_DESC_A_XUSER_11_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h40
`define WR_RESP_DESC_A_XUSER_12_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h44
`define WR_RESP_DESC_A_XUSER_13_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h48
`define WR_RESP_DESC_A_XUSER_14_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h4C
`define WR_RESP_DESC_A_XUSER_15_REG_ADDR `WR_RESP_DESC_A_BASE_ADDR + 'h50
`define SN_REQ_DESC_A_ATTR_REG_ADDR `SN_REQ_DESC_A_BASE_ADDR + 'h0
`define SN_REQ_DESC_A_ACADDR_0_REG_ADDR `SN_REQ_DESC_A_BASE_ADDR + 'h4
`define SN_REQ_DESC_A_ACADDR_1_REG_ADDR `SN_REQ_DESC_A_BASE_ADDR + 'h8
`define SN_REQ_DESC_A_ACADDR_2_REG_ADDR `SN_REQ_DESC_A_BASE_ADDR + 'hC
`define SN_REQ_DESC_A_ACADDR_3_REG_ADDR `SN_REQ_DESC_A_BASE_ADDR + 'h10
`define SN_RESP_DESC_A_RESP_REG_ADDR `SN_RESP_DESC_A_BASE_ADDR + 'h0


`define RD_REQ_DESC_B_TXN_TYPE_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h0
`define RD_REQ_DESC_B_SIZE_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h4
`define RD_REQ_DESC_B_AXSIZE_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h8
`define RD_REQ_DESC_B_ATTR_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'hC
`define RD_REQ_DESC_B_AXADDR_0_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h10
`define RD_REQ_DESC_B_AXADDR_1_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h14
`define RD_REQ_DESC_B_AXADDR_2_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h18
`define RD_REQ_DESC_B_AXADDR_3_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h1C
`define RD_REQ_DESC_B_AXID_0_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h20
`define RD_REQ_DESC_B_AXID_1_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h24
`define RD_REQ_DESC_B_AXID_2_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h28
`define RD_REQ_DESC_B_AXID_3_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h2C
`define RD_REQ_DESC_B_AXUSER_0_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h30
`define RD_REQ_DESC_B_AXUSER_1_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h34
`define RD_REQ_DESC_B_AXUSER_2_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h38
`define RD_REQ_DESC_B_AXUSER_3_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h3C
`define RD_REQ_DESC_B_AXUSER_4_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h40
`define RD_REQ_DESC_B_AXUSER_5_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h44
`define RD_REQ_DESC_B_AXUSER_6_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h48
`define RD_REQ_DESC_B_AXUSER_7_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h4C
`define RD_REQ_DESC_B_AXUSER_8_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h50
`define RD_REQ_DESC_B_AXUSER_9_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h54
`define RD_REQ_DESC_B_AXUSER_10_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h58
`define RD_REQ_DESC_B_AXUSER_11_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h5C
`define RD_REQ_DESC_B_AXUSER_12_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h60
`define RD_REQ_DESC_B_AXUSER_13_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h64
`define RD_REQ_DESC_B_AXUSER_14_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h68
`define RD_REQ_DESC_B_AXUSER_15_REG_ADDR `RD_REQ_DESC_B_BASE_ADDR + 'h6C
`define RD_RESP_DESC_B_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h0
`define RD_RESP_DESC_B_DATA_SIZE_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h4
`define RD_RESP_DESC_B_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h8
`define RD_RESP_DESC_B_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'hC
`define RD_RESP_DESC_B_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h10
`define RD_RESP_DESC_B_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h14
`define RD_RESP_DESC_B_RESP_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h18
`define RD_RESP_DESC_B_XID_0_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h1C
`define RD_RESP_DESC_B_XID_1_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h20
`define RD_RESP_DESC_B_XID_2_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h24
`define RD_RESP_DESC_B_XID_3_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h28
`define RD_RESP_DESC_B_XUSER_0_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h2C
`define RD_RESP_DESC_B_XUSER_1_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h30
`define RD_RESP_DESC_B_XUSER_2_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h34
`define RD_RESP_DESC_B_XUSER_3_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h38
`define RD_RESP_DESC_B_XUSER_4_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h3C
`define RD_RESP_DESC_B_XUSER_5_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h40
`define RD_RESP_DESC_B_XUSER_6_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h44
`define RD_RESP_DESC_B_XUSER_7_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h48
`define RD_RESP_DESC_B_XUSER_8_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h4C
`define RD_RESP_DESC_B_XUSER_9_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h50
`define RD_RESP_DESC_B_XUSER_10_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h54
`define RD_RESP_DESC_B_XUSER_11_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h58
`define RD_RESP_DESC_B_XUSER_12_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h5C
`define RD_RESP_DESC_B_XUSER_13_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h60
`define RD_RESP_DESC_B_XUSER_14_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h64
`define RD_RESP_DESC_B_XUSER_15_REG_ADDR `RD_RESP_DESC_B_BASE_ADDR + 'h68
`define WR_REQ_DESC_B_TXN_TYPE_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h0
`define WR_REQ_DESC_B_SIZE_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h4
`define WR_REQ_DESC_B_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h8
`define WR_REQ_DESC_B_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hC
`define WR_REQ_DESC_B_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h10
`define WR_REQ_DESC_B_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h14
`define WR_REQ_DESC_B_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h18
`define WR_REQ_DESC_B_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h1C
`define WR_REQ_DESC_B_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h20
`define WR_REQ_DESC_B_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h24
`define WR_REQ_DESC_B_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h28
`define WR_REQ_DESC_B_AXSIZE_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h2C
`define WR_REQ_DESC_B_ATTR_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h30
`define WR_REQ_DESC_B_AXADDR_0_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h34
`define WR_REQ_DESC_B_AXADDR_1_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h38
`define WR_REQ_DESC_B_AXADDR_2_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h3C
`define WR_REQ_DESC_B_AXADDR_3_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h40
`define WR_REQ_DESC_B_AXID_0_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h44
`define WR_REQ_DESC_B_AXID_1_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h48
`define WR_REQ_DESC_B_AXID_2_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h4C
`define WR_REQ_DESC_B_AXID_3_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h50
`define WR_REQ_DESC_B_AXUSER_0_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h54
`define WR_REQ_DESC_B_AXUSER_1_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h58
`define WR_REQ_DESC_B_AXUSER_2_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h5C
`define WR_REQ_DESC_B_AXUSER_3_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h60
`define WR_REQ_DESC_B_AXUSER_4_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h64
`define WR_REQ_DESC_B_AXUSER_5_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h68
`define WR_REQ_DESC_B_AXUSER_6_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h6C
`define WR_REQ_DESC_B_AXUSER_7_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h70
`define WR_REQ_DESC_B_AXUSER_8_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h74
`define WR_REQ_DESC_B_AXUSER_9_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h78
`define WR_REQ_DESC_B_AXUSER_10_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h7C
`define WR_REQ_DESC_B_AXUSER_11_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h80
`define WR_REQ_DESC_B_AXUSER_12_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h84
`define WR_REQ_DESC_B_AXUSER_13_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h88
`define WR_REQ_DESC_B_AXUSER_14_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h8C
`define WR_REQ_DESC_B_AXUSER_15_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h90
`define WR_REQ_DESC_B_WUSER_0_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h94
`define WR_REQ_DESC_B_WUSER_1_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h98
`define WR_REQ_DESC_B_WUSER_2_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'h9C
`define WR_REQ_DESC_B_WUSER_3_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hA0
`define WR_REQ_DESC_B_WUSER_4_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hA4
`define WR_REQ_DESC_B_WUSER_5_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hA8
`define WR_REQ_DESC_B_WUSER_6_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hAC
`define WR_REQ_DESC_B_WUSER_7_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hB0
`define WR_REQ_DESC_B_WUSER_8_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hB4
`define WR_REQ_DESC_B_WUSER_9_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hB8
`define WR_REQ_DESC_B_WUSER_10_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hBC
`define WR_REQ_DESC_B_WUSER_11_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hC0
`define WR_REQ_DESC_B_WUSER_12_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hC4
`define WR_REQ_DESC_B_WUSER_13_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hC8
`define WR_REQ_DESC_B_WUSER_14_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hCC
`define WR_REQ_DESC_B_WUSER_15_REG_ADDR `WR_REQ_DESC_B_BASE_ADDR + 'hD0
`define WR_RESP_DESC_B_RESP_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h0
`define WR_RESP_DESC_B_XID_0_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h4
`define WR_RESP_DESC_B_XID_1_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h8
`define WR_RESP_DESC_B_XID_2_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'hC
`define WR_RESP_DESC_B_XID_3_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h10
`define WR_RESP_DESC_B_XUSER_0_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h14
`define WR_RESP_DESC_B_XUSER_1_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h18
`define WR_RESP_DESC_B_XUSER_2_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h1C
`define WR_RESP_DESC_B_XUSER_3_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h20
`define WR_RESP_DESC_B_XUSER_4_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h24
`define WR_RESP_DESC_B_XUSER_5_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h28
`define WR_RESP_DESC_B_XUSER_6_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h2C
`define WR_RESP_DESC_B_XUSER_7_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h30
`define WR_RESP_DESC_B_XUSER_8_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h34
`define WR_RESP_DESC_B_XUSER_9_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h38
`define WR_RESP_DESC_B_XUSER_10_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h3C
`define WR_RESP_DESC_B_XUSER_11_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h40
`define WR_RESP_DESC_B_XUSER_12_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h44
`define WR_RESP_DESC_B_XUSER_13_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h48
`define WR_RESP_DESC_B_XUSER_14_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h4C
`define WR_RESP_DESC_B_XUSER_15_REG_ADDR `WR_RESP_DESC_B_BASE_ADDR + 'h50
`define SN_REQ_DESC_B_ATTR_REG_ADDR `SN_REQ_DESC_B_BASE_ADDR + 'h0
`define SN_REQ_DESC_B_ACADDR_0_REG_ADDR `SN_REQ_DESC_B_BASE_ADDR + 'h4
`define SN_REQ_DESC_B_ACADDR_1_REG_ADDR `SN_REQ_DESC_B_BASE_ADDR + 'h8
`define SN_REQ_DESC_B_ACADDR_2_REG_ADDR `SN_REQ_DESC_B_BASE_ADDR + 'hC
`define SN_REQ_DESC_B_ACADDR_3_REG_ADDR `SN_REQ_DESC_B_BASE_ADDR + 'h10
`define SN_RESP_DESC_B_RESP_REG_ADDR `SN_RESP_DESC_B_BASE_ADDR + 'h0


`define RD_REQ_DESC_C_TXN_TYPE_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h0
`define RD_REQ_DESC_C_SIZE_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h4
`define RD_REQ_DESC_C_AXSIZE_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h8
`define RD_REQ_DESC_C_ATTR_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'hC
`define RD_REQ_DESC_C_AXADDR_0_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h10
`define RD_REQ_DESC_C_AXADDR_1_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h14
`define RD_REQ_DESC_C_AXADDR_2_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h18
`define RD_REQ_DESC_C_AXADDR_3_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h1C
`define RD_REQ_DESC_C_AXID_0_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h20
`define RD_REQ_DESC_C_AXID_1_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h24
`define RD_REQ_DESC_C_AXID_2_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h28
`define RD_REQ_DESC_C_AXID_3_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h2C
`define RD_REQ_DESC_C_AXUSER_0_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h30
`define RD_REQ_DESC_C_AXUSER_1_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h34
`define RD_REQ_DESC_C_AXUSER_2_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h38
`define RD_REQ_DESC_C_AXUSER_3_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h3C
`define RD_REQ_DESC_C_AXUSER_4_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h40
`define RD_REQ_DESC_C_AXUSER_5_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h44
`define RD_REQ_DESC_C_AXUSER_6_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h48
`define RD_REQ_DESC_C_AXUSER_7_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h4C
`define RD_REQ_DESC_C_AXUSER_8_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h50
`define RD_REQ_DESC_C_AXUSER_9_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h54
`define RD_REQ_DESC_C_AXUSER_10_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h58
`define RD_REQ_DESC_C_AXUSER_11_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h5C
`define RD_REQ_DESC_C_AXUSER_12_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h60
`define RD_REQ_DESC_C_AXUSER_13_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h64
`define RD_REQ_DESC_C_AXUSER_14_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h68
`define RD_REQ_DESC_C_AXUSER_15_REG_ADDR `RD_REQ_DESC_C_BASE_ADDR + 'h6C
`define RD_RESP_DESC_C_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h0
`define RD_RESP_DESC_C_DATA_SIZE_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h4
`define RD_RESP_DESC_C_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h8
`define RD_RESP_DESC_C_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'hC
`define RD_RESP_DESC_C_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h10
`define RD_RESP_DESC_C_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h14
`define RD_RESP_DESC_C_RESP_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h18
`define RD_RESP_DESC_C_XID_0_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h1C
`define RD_RESP_DESC_C_XID_1_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h20
`define RD_RESP_DESC_C_XID_2_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h24
`define RD_RESP_DESC_C_XID_3_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h28
`define RD_RESP_DESC_C_XUSER_0_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h2C
`define RD_RESP_DESC_C_XUSER_1_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h30
`define RD_RESP_DESC_C_XUSER_2_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h34
`define RD_RESP_DESC_C_XUSER_3_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h38
`define RD_RESP_DESC_C_XUSER_4_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h3C
`define RD_RESP_DESC_C_XUSER_5_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h40
`define RD_RESP_DESC_C_XUSER_6_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h44
`define RD_RESP_DESC_C_XUSER_7_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h48
`define RD_RESP_DESC_C_XUSER_8_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h4C
`define RD_RESP_DESC_C_XUSER_9_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h50
`define RD_RESP_DESC_C_XUSER_10_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h54
`define RD_RESP_DESC_C_XUSER_11_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h58
`define RD_RESP_DESC_C_XUSER_12_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h5C
`define RD_RESP_DESC_C_XUSER_13_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h60
`define RD_RESP_DESC_C_XUSER_14_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h64
`define RD_RESP_DESC_C_XUSER_15_REG_ADDR `RD_RESP_DESC_C_BASE_ADDR + 'h68
`define WR_REQ_DESC_C_TXN_TYPE_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h0
`define WR_REQ_DESC_C_SIZE_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h4
`define WR_REQ_DESC_C_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h8
`define WR_REQ_DESC_C_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hC
`define WR_REQ_DESC_C_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h10
`define WR_REQ_DESC_C_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h14
`define WR_REQ_DESC_C_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h18
`define WR_REQ_DESC_C_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h1C
`define WR_REQ_DESC_C_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h20
`define WR_REQ_DESC_C_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h24
`define WR_REQ_DESC_C_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h28
`define WR_REQ_DESC_C_AXSIZE_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h2C
`define WR_REQ_DESC_C_ATTR_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h30
`define WR_REQ_DESC_C_AXADDR_0_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h34
`define WR_REQ_DESC_C_AXADDR_1_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h38
`define WR_REQ_DESC_C_AXADDR_2_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h3C
`define WR_REQ_DESC_C_AXADDR_3_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h40
`define WR_REQ_DESC_C_AXID_0_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h44
`define WR_REQ_DESC_C_AXID_1_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h48
`define WR_REQ_DESC_C_AXID_2_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h4C
`define WR_REQ_DESC_C_AXID_3_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h50
`define WR_REQ_DESC_C_AXUSER_0_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h54
`define WR_REQ_DESC_C_AXUSER_1_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h58
`define WR_REQ_DESC_C_AXUSER_2_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h5C
`define WR_REQ_DESC_C_AXUSER_3_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h60
`define WR_REQ_DESC_C_AXUSER_4_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h64
`define WR_REQ_DESC_C_AXUSER_5_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h68
`define WR_REQ_DESC_C_AXUSER_6_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h6C
`define WR_REQ_DESC_C_AXUSER_7_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h70
`define WR_REQ_DESC_C_AXUSER_8_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h74
`define WR_REQ_DESC_C_AXUSER_9_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h78
`define WR_REQ_DESC_C_AXUSER_10_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h7C
`define WR_REQ_DESC_C_AXUSER_11_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h80
`define WR_REQ_DESC_C_AXUSER_12_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h84
`define WR_REQ_DESC_C_AXUSER_13_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h88
`define WR_REQ_DESC_C_AXUSER_14_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h8C
`define WR_REQ_DESC_C_AXUSER_15_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h90
`define WR_REQ_DESC_C_WUSER_0_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h94
`define WR_REQ_DESC_C_WUSER_1_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h98
`define WR_REQ_DESC_C_WUSER_2_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'h9C
`define WR_REQ_DESC_C_WUSER_3_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hA0
`define WR_REQ_DESC_C_WUSER_4_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hA4
`define WR_REQ_DESC_C_WUSER_5_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hA8
`define WR_REQ_DESC_C_WUSER_6_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hAC
`define WR_REQ_DESC_C_WUSER_7_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hB0
`define WR_REQ_DESC_C_WUSER_8_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hB4
`define WR_REQ_DESC_C_WUSER_9_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hB8
`define WR_REQ_DESC_C_WUSER_10_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hBC
`define WR_REQ_DESC_C_WUSER_11_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hC0
`define WR_REQ_DESC_C_WUSER_12_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hC4
`define WR_REQ_DESC_C_WUSER_13_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hC8
`define WR_REQ_DESC_C_WUSER_14_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hCC
`define WR_REQ_DESC_C_WUSER_15_REG_ADDR `WR_REQ_DESC_C_BASE_ADDR + 'hD0
`define WR_RESP_DESC_C_RESP_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h0
`define WR_RESP_DESC_C_XID_0_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h4
`define WR_RESP_DESC_C_XID_1_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h8
`define WR_RESP_DESC_C_XID_2_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'hC
`define WR_RESP_DESC_C_XID_3_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h10
`define WR_RESP_DESC_C_XUSER_0_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h14
`define WR_RESP_DESC_C_XUSER_1_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h18
`define WR_RESP_DESC_C_XUSER_2_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h1C
`define WR_RESP_DESC_C_XUSER_3_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h20
`define WR_RESP_DESC_C_XUSER_4_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h24
`define WR_RESP_DESC_C_XUSER_5_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h28
`define WR_RESP_DESC_C_XUSER_6_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h2C
`define WR_RESP_DESC_C_XUSER_7_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h30
`define WR_RESP_DESC_C_XUSER_8_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h34
`define WR_RESP_DESC_C_XUSER_9_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h38
`define WR_RESP_DESC_C_XUSER_10_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h3C
`define WR_RESP_DESC_C_XUSER_11_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h40
`define WR_RESP_DESC_C_XUSER_12_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h44
`define WR_RESP_DESC_C_XUSER_13_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h48
`define WR_RESP_DESC_C_XUSER_14_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h4C
`define WR_RESP_DESC_C_XUSER_15_REG_ADDR `WR_RESP_DESC_C_BASE_ADDR + 'h50
`define SN_REQ_DESC_C_ATTR_REG_ADDR `SN_REQ_DESC_C_BASE_ADDR + 'h0
`define SN_REQ_DESC_C_ACADDR_0_REG_ADDR `SN_REQ_DESC_C_BASE_ADDR + 'h4
`define SN_REQ_DESC_C_ACADDR_1_REG_ADDR `SN_REQ_DESC_C_BASE_ADDR + 'h8
`define SN_REQ_DESC_C_ACADDR_2_REG_ADDR `SN_REQ_DESC_C_BASE_ADDR + 'hC
`define SN_REQ_DESC_C_ACADDR_3_REG_ADDR `SN_REQ_DESC_C_BASE_ADDR + 'h10
`define SN_RESP_DESC_C_RESP_REG_ADDR `SN_RESP_DESC_C_BASE_ADDR + 'h0


`define RD_REQ_DESC_D_TXN_TYPE_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h0
`define RD_REQ_DESC_D_SIZE_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h4
`define RD_REQ_DESC_D_AXSIZE_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h8
`define RD_REQ_DESC_D_ATTR_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'hC
`define RD_REQ_DESC_D_AXADDR_0_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h10
`define RD_REQ_DESC_D_AXADDR_1_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h14
`define RD_REQ_DESC_D_AXADDR_2_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h18
`define RD_REQ_DESC_D_AXADDR_3_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h1C
`define RD_REQ_DESC_D_AXID_0_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h20
`define RD_REQ_DESC_D_AXID_1_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h24
`define RD_REQ_DESC_D_AXID_2_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h28
`define RD_REQ_DESC_D_AXID_3_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h2C
`define RD_REQ_DESC_D_AXUSER_0_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h30
`define RD_REQ_DESC_D_AXUSER_1_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h34
`define RD_REQ_DESC_D_AXUSER_2_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h38
`define RD_REQ_DESC_D_AXUSER_3_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h3C
`define RD_REQ_DESC_D_AXUSER_4_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h40
`define RD_REQ_DESC_D_AXUSER_5_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h44
`define RD_REQ_DESC_D_AXUSER_6_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h48
`define RD_REQ_DESC_D_AXUSER_7_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h4C
`define RD_REQ_DESC_D_AXUSER_8_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h50
`define RD_REQ_DESC_D_AXUSER_9_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h54
`define RD_REQ_DESC_D_AXUSER_10_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h58
`define RD_REQ_DESC_D_AXUSER_11_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h5C
`define RD_REQ_DESC_D_AXUSER_12_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h60
`define RD_REQ_DESC_D_AXUSER_13_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h64
`define RD_REQ_DESC_D_AXUSER_14_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h68
`define RD_REQ_DESC_D_AXUSER_15_REG_ADDR `RD_REQ_DESC_D_BASE_ADDR + 'h6C
`define RD_RESP_DESC_D_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h0
`define RD_RESP_DESC_D_DATA_SIZE_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h4
`define RD_RESP_DESC_D_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h8
`define RD_RESP_DESC_D_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'hC
`define RD_RESP_DESC_D_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h10
`define RD_RESP_DESC_D_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h14
`define RD_RESP_DESC_D_RESP_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h18
`define RD_RESP_DESC_D_XID_0_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h1C
`define RD_RESP_DESC_D_XID_1_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h20
`define RD_RESP_DESC_D_XID_2_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h24
`define RD_RESP_DESC_D_XID_3_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h28
`define RD_RESP_DESC_D_XUSER_0_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h2C
`define RD_RESP_DESC_D_XUSER_1_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h30
`define RD_RESP_DESC_D_XUSER_2_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h34
`define RD_RESP_DESC_D_XUSER_3_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h38
`define RD_RESP_DESC_D_XUSER_4_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h3C
`define RD_RESP_DESC_D_XUSER_5_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h40
`define RD_RESP_DESC_D_XUSER_6_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h44
`define RD_RESP_DESC_D_XUSER_7_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h48
`define RD_RESP_DESC_D_XUSER_8_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h4C
`define RD_RESP_DESC_D_XUSER_9_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h50
`define RD_RESP_DESC_D_XUSER_10_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h54
`define RD_RESP_DESC_D_XUSER_11_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h58
`define RD_RESP_DESC_D_XUSER_12_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h5C
`define RD_RESP_DESC_D_XUSER_13_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h60
`define RD_RESP_DESC_D_XUSER_14_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h64
`define RD_RESP_DESC_D_XUSER_15_REG_ADDR `RD_RESP_DESC_D_BASE_ADDR + 'h68
`define WR_REQ_DESC_D_TXN_TYPE_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h0
`define WR_REQ_DESC_D_SIZE_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h4
`define WR_REQ_DESC_D_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h8
`define WR_REQ_DESC_D_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hC
`define WR_REQ_DESC_D_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h10
`define WR_REQ_DESC_D_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h14
`define WR_REQ_DESC_D_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h18
`define WR_REQ_DESC_D_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h1C
`define WR_REQ_DESC_D_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h20
`define WR_REQ_DESC_D_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h24
`define WR_REQ_DESC_D_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h28
`define WR_REQ_DESC_D_AXSIZE_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h2C
`define WR_REQ_DESC_D_ATTR_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h30
`define WR_REQ_DESC_D_AXADDR_0_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h34
`define WR_REQ_DESC_D_AXADDR_1_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h38
`define WR_REQ_DESC_D_AXADDR_2_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h3C
`define WR_REQ_DESC_D_AXADDR_3_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h40
`define WR_REQ_DESC_D_AXID_0_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h44
`define WR_REQ_DESC_D_AXID_1_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h48
`define WR_REQ_DESC_D_AXID_2_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h4C
`define WR_REQ_DESC_D_AXID_3_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h50
`define WR_REQ_DESC_D_AXUSER_0_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h54
`define WR_REQ_DESC_D_AXUSER_1_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h58
`define WR_REQ_DESC_D_AXUSER_2_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h5C
`define WR_REQ_DESC_D_AXUSER_3_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h60
`define WR_REQ_DESC_D_AXUSER_4_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h64
`define WR_REQ_DESC_D_AXUSER_5_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h68
`define WR_REQ_DESC_D_AXUSER_6_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h6C
`define WR_REQ_DESC_D_AXUSER_7_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h70
`define WR_REQ_DESC_D_AXUSER_8_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h74
`define WR_REQ_DESC_D_AXUSER_9_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h78
`define WR_REQ_DESC_D_AXUSER_10_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h7C
`define WR_REQ_DESC_D_AXUSER_11_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h80
`define WR_REQ_DESC_D_AXUSER_12_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h84
`define WR_REQ_DESC_D_AXUSER_13_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h88
`define WR_REQ_DESC_D_AXUSER_14_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h8C
`define WR_REQ_DESC_D_AXUSER_15_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h90
`define WR_REQ_DESC_D_WUSER_0_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h94
`define WR_REQ_DESC_D_WUSER_1_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h98
`define WR_REQ_DESC_D_WUSER_2_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'h9C
`define WR_REQ_DESC_D_WUSER_3_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hA0
`define WR_REQ_DESC_D_WUSER_4_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hA4
`define WR_REQ_DESC_D_WUSER_5_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hA8
`define WR_REQ_DESC_D_WUSER_6_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hAC
`define WR_REQ_DESC_D_WUSER_7_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hB0
`define WR_REQ_DESC_D_WUSER_8_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hB4
`define WR_REQ_DESC_D_WUSER_9_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hB8
`define WR_REQ_DESC_D_WUSER_10_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hBC
`define WR_REQ_DESC_D_WUSER_11_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hC0
`define WR_REQ_DESC_D_WUSER_12_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hC4
`define WR_REQ_DESC_D_WUSER_13_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hC8
`define WR_REQ_DESC_D_WUSER_14_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hCC
`define WR_REQ_DESC_D_WUSER_15_REG_ADDR `WR_REQ_DESC_D_BASE_ADDR + 'hD0
`define WR_RESP_DESC_D_RESP_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h0
`define WR_RESP_DESC_D_XID_0_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h4
`define WR_RESP_DESC_D_XID_1_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h8
`define WR_RESP_DESC_D_XID_2_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'hC
`define WR_RESP_DESC_D_XID_3_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h10
`define WR_RESP_DESC_D_XUSER_0_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h14
`define WR_RESP_DESC_D_XUSER_1_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h18
`define WR_RESP_DESC_D_XUSER_2_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h1C
`define WR_RESP_DESC_D_XUSER_3_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h20
`define WR_RESP_DESC_D_XUSER_4_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h24
`define WR_RESP_DESC_D_XUSER_5_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h28
`define WR_RESP_DESC_D_XUSER_6_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h2C
`define WR_RESP_DESC_D_XUSER_7_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h30
`define WR_RESP_DESC_D_XUSER_8_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h34
`define WR_RESP_DESC_D_XUSER_9_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h38
`define WR_RESP_DESC_D_XUSER_10_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h3C
`define WR_RESP_DESC_D_XUSER_11_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h40
`define WR_RESP_DESC_D_XUSER_12_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h44
`define WR_RESP_DESC_D_XUSER_13_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h48
`define WR_RESP_DESC_D_XUSER_14_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h4C
`define WR_RESP_DESC_D_XUSER_15_REG_ADDR `WR_RESP_DESC_D_BASE_ADDR + 'h50
`define SN_REQ_DESC_D_ATTR_REG_ADDR `SN_REQ_DESC_D_BASE_ADDR + 'h0
`define SN_REQ_DESC_D_ACADDR_0_REG_ADDR `SN_REQ_DESC_D_BASE_ADDR + 'h4
`define SN_REQ_DESC_D_ACADDR_1_REG_ADDR `SN_REQ_DESC_D_BASE_ADDR + 'h8
`define SN_REQ_DESC_D_ACADDR_2_REG_ADDR `SN_REQ_DESC_D_BASE_ADDR + 'hC
`define SN_REQ_DESC_D_ACADDR_3_REG_ADDR `SN_REQ_DESC_D_BASE_ADDR + 'h10
`define SN_RESP_DESC_D_RESP_REG_ADDR `SN_RESP_DESC_D_BASE_ADDR + 'h0


`define RD_REQ_DESC_E_TXN_TYPE_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h0
`define RD_REQ_DESC_E_SIZE_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h4
`define RD_REQ_DESC_E_AXSIZE_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h8
`define RD_REQ_DESC_E_ATTR_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'hC
`define RD_REQ_DESC_E_AXADDR_0_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h10
`define RD_REQ_DESC_E_AXADDR_1_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h14
`define RD_REQ_DESC_E_AXADDR_2_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h18
`define RD_REQ_DESC_E_AXADDR_3_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h1C
`define RD_REQ_DESC_E_AXID_0_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h20
`define RD_REQ_DESC_E_AXID_1_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h24
`define RD_REQ_DESC_E_AXID_2_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h28
`define RD_REQ_DESC_E_AXID_3_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h2C
`define RD_REQ_DESC_E_AXUSER_0_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h30
`define RD_REQ_DESC_E_AXUSER_1_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h34
`define RD_REQ_DESC_E_AXUSER_2_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h38
`define RD_REQ_DESC_E_AXUSER_3_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h3C
`define RD_REQ_DESC_E_AXUSER_4_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h40
`define RD_REQ_DESC_E_AXUSER_5_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h44
`define RD_REQ_DESC_E_AXUSER_6_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h48
`define RD_REQ_DESC_E_AXUSER_7_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h4C
`define RD_REQ_DESC_E_AXUSER_8_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h50
`define RD_REQ_DESC_E_AXUSER_9_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h54
`define RD_REQ_DESC_E_AXUSER_10_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h58
`define RD_REQ_DESC_E_AXUSER_11_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h5C
`define RD_REQ_DESC_E_AXUSER_12_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h60
`define RD_REQ_DESC_E_AXUSER_13_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h64
`define RD_REQ_DESC_E_AXUSER_14_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h68
`define RD_REQ_DESC_E_AXUSER_15_REG_ADDR `RD_REQ_DESC_E_BASE_ADDR + 'h6C
`define RD_RESP_DESC_E_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h0
`define RD_RESP_DESC_E_DATA_SIZE_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h4
`define RD_RESP_DESC_E_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h8
`define RD_RESP_DESC_E_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'hC
`define RD_RESP_DESC_E_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h10
`define RD_RESP_DESC_E_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h14
`define RD_RESP_DESC_E_RESP_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h18
`define RD_RESP_DESC_E_XID_0_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h1C
`define RD_RESP_DESC_E_XID_1_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h20
`define RD_RESP_DESC_E_XID_2_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h24
`define RD_RESP_DESC_E_XID_3_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h28
`define RD_RESP_DESC_E_XUSER_0_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h2C
`define RD_RESP_DESC_E_XUSER_1_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h30
`define RD_RESP_DESC_E_XUSER_2_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h34
`define RD_RESP_DESC_E_XUSER_3_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h38
`define RD_RESP_DESC_E_XUSER_4_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h3C
`define RD_RESP_DESC_E_XUSER_5_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h40
`define RD_RESP_DESC_E_XUSER_6_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h44
`define RD_RESP_DESC_E_XUSER_7_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h48
`define RD_RESP_DESC_E_XUSER_8_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h4C
`define RD_RESP_DESC_E_XUSER_9_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h50
`define RD_RESP_DESC_E_XUSER_10_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h54
`define RD_RESP_DESC_E_XUSER_11_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h58
`define RD_RESP_DESC_E_XUSER_12_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h5C
`define RD_RESP_DESC_E_XUSER_13_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h60
`define RD_RESP_DESC_E_XUSER_14_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h64
`define RD_RESP_DESC_E_XUSER_15_REG_ADDR `RD_RESP_DESC_E_BASE_ADDR + 'h68
`define WR_REQ_DESC_E_TXN_TYPE_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h0
`define WR_REQ_DESC_E_SIZE_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h4
`define WR_REQ_DESC_E_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h8
`define WR_REQ_DESC_E_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hC
`define WR_REQ_DESC_E_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h10
`define WR_REQ_DESC_E_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h14
`define WR_REQ_DESC_E_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h18
`define WR_REQ_DESC_E_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h1C
`define WR_REQ_DESC_E_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h20
`define WR_REQ_DESC_E_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h24
`define WR_REQ_DESC_E_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h28
`define WR_REQ_DESC_E_AXSIZE_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h2C
`define WR_REQ_DESC_E_ATTR_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h30
`define WR_REQ_DESC_E_AXADDR_0_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h34
`define WR_REQ_DESC_E_AXADDR_1_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h38
`define WR_REQ_DESC_E_AXADDR_2_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h3C
`define WR_REQ_DESC_E_AXADDR_3_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h40
`define WR_REQ_DESC_E_AXID_0_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h44
`define WR_REQ_DESC_E_AXID_1_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h48
`define WR_REQ_DESC_E_AXID_2_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h4C
`define WR_REQ_DESC_E_AXID_3_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h50
`define WR_REQ_DESC_E_AXUSER_0_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h54
`define WR_REQ_DESC_E_AXUSER_1_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h58
`define WR_REQ_DESC_E_AXUSER_2_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h5C
`define WR_REQ_DESC_E_AXUSER_3_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h60
`define WR_REQ_DESC_E_AXUSER_4_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h64
`define WR_REQ_DESC_E_AXUSER_5_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h68
`define WR_REQ_DESC_E_AXUSER_6_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h6C
`define WR_REQ_DESC_E_AXUSER_7_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h70
`define WR_REQ_DESC_E_AXUSER_8_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h74
`define WR_REQ_DESC_E_AXUSER_9_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h78
`define WR_REQ_DESC_E_AXUSER_10_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h7C
`define WR_REQ_DESC_E_AXUSER_11_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h80
`define WR_REQ_DESC_E_AXUSER_12_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h84
`define WR_REQ_DESC_E_AXUSER_13_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h88
`define WR_REQ_DESC_E_AXUSER_14_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h8C
`define WR_REQ_DESC_E_AXUSER_15_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h90
`define WR_REQ_DESC_E_WUSER_0_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h94
`define WR_REQ_DESC_E_WUSER_1_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h98
`define WR_REQ_DESC_E_WUSER_2_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'h9C
`define WR_REQ_DESC_E_WUSER_3_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hA0
`define WR_REQ_DESC_E_WUSER_4_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hA4
`define WR_REQ_DESC_E_WUSER_5_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hA8
`define WR_REQ_DESC_E_WUSER_6_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hAC
`define WR_REQ_DESC_E_WUSER_7_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hB0
`define WR_REQ_DESC_E_WUSER_8_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hB4
`define WR_REQ_DESC_E_WUSER_9_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hB8
`define WR_REQ_DESC_E_WUSER_10_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hBC
`define WR_REQ_DESC_E_WUSER_11_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hC0
`define WR_REQ_DESC_E_WUSER_12_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hC4
`define WR_REQ_DESC_E_WUSER_13_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hC8
`define WR_REQ_DESC_E_WUSER_14_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hCC
`define WR_REQ_DESC_E_WUSER_15_REG_ADDR `WR_REQ_DESC_E_BASE_ADDR + 'hD0
`define WR_RESP_DESC_E_RESP_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h0
`define WR_RESP_DESC_E_XID_0_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h4
`define WR_RESP_DESC_E_XID_1_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h8
`define WR_RESP_DESC_E_XID_2_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'hC
`define WR_RESP_DESC_E_XID_3_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h10
`define WR_RESP_DESC_E_XUSER_0_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h14
`define WR_RESP_DESC_E_XUSER_1_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h18
`define WR_RESP_DESC_E_XUSER_2_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h1C
`define WR_RESP_DESC_E_XUSER_3_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h20
`define WR_RESP_DESC_E_XUSER_4_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h24
`define WR_RESP_DESC_E_XUSER_5_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h28
`define WR_RESP_DESC_E_XUSER_6_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h2C
`define WR_RESP_DESC_E_XUSER_7_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h30
`define WR_RESP_DESC_E_XUSER_8_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h34
`define WR_RESP_DESC_E_XUSER_9_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h38
`define WR_RESP_DESC_E_XUSER_10_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h3C
`define WR_RESP_DESC_E_XUSER_11_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h40
`define WR_RESP_DESC_E_XUSER_12_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h44
`define WR_RESP_DESC_E_XUSER_13_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h48
`define WR_RESP_DESC_E_XUSER_14_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h4C
`define WR_RESP_DESC_E_XUSER_15_REG_ADDR `WR_RESP_DESC_E_BASE_ADDR + 'h50
`define SN_REQ_DESC_E_ATTR_REG_ADDR `SN_REQ_DESC_E_BASE_ADDR + 'h0
`define SN_REQ_DESC_E_ACADDR_0_REG_ADDR `SN_REQ_DESC_E_BASE_ADDR + 'h4
`define SN_REQ_DESC_E_ACADDR_1_REG_ADDR `SN_REQ_DESC_E_BASE_ADDR + 'h8
`define SN_REQ_DESC_E_ACADDR_2_REG_ADDR `SN_REQ_DESC_E_BASE_ADDR + 'hC
`define SN_REQ_DESC_E_ACADDR_3_REG_ADDR `SN_REQ_DESC_E_BASE_ADDR + 'h10
`define SN_RESP_DESC_E_RESP_REG_ADDR `SN_RESP_DESC_E_BASE_ADDR + 'h0


`define RD_REQ_DESC_F_TXN_TYPE_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h0
`define RD_REQ_DESC_F_SIZE_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h4
`define RD_REQ_DESC_F_AXSIZE_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h8
`define RD_REQ_DESC_F_ATTR_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'hC
`define RD_REQ_DESC_F_AXADDR_0_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h10
`define RD_REQ_DESC_F_AXADDR_1_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h14
`define RD_REQ_DESC_F_AXADDR_2_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h18
`define RD_REQ_DESC_F_AXADDR_3_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h1C
`define RD_REQ_DESC_F_AXID_0_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h20
`define RD_REQ_DESC_F_AXID_1_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h24
`define RD_REQ_DESC_F_AXID_2_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h28
`define RD_REQ_DESC_F_AXID_3_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h2C
`define RD_REQ_DESC_F_AXUSER_0_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h30
`define RD_REQ_DESC_F_AXUSER_1_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h34
`define RD_REQ_DESC_F_AXUSER_2_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h38
`define RD_REQ_DESC_F_AXUSER_3_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h3C
`define RD_REQ_DESC_F_AXUSER_4_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h40
`define RD_REQ_DESC_F_AXUSER_5_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h44
`define RD_REQ_DESC_F_AXUSER_6_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h48
`define RD_REQ_DESC_F_AXUSER_7_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h4C
`define RD_REQ_DESC_F_AXUSER_8_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h50
`define RD_REQ_DESC_F_AXUSER_9_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h54
`define RD_REQ_DESC_F_AXUSER_10_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h58
`define RD_REQ_DESC_F_AXUSER_11_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h5C
`define RD_REQ_DESC_F_AXUSER_12_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h60
`define RD_REQ_DESC_F_AXUSER_13_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h64
`define RD_REQ_DESC_F_AXUSER_14_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h68
`define RD_REQ_DESC_F_AXUSER_15_REG_ADDR `RD_REQ_DESC_F_BASE_ADDR + 'h6C
`define RD_RESP_DESC_F_DATA_OFFSET_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h0
`define RD_RESP_DESC_F_DATA_SIZE_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h4
`define RD_RESP_DESC_F_DATA_HOST_ADDR_0_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h8
`define RD_RESP_DESC_F_DATA_HOST_ADDR_1_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'hC
`define RD_RESP_DESC_F_DATA_HOST_ADDR_2_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h10
`define RD_RESP_DESC_F_DATA_HOST_ADDR_3_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h14
`define RD_RESP_DESC_F_RESP_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h18
`define RD_RESP_DESC_F_XID_0_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h1C
`define RD_RESP_DESC_F_XID_1_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h20
`define RD_RESP_DESC_F_XID_2_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h24
`define RD_RESP_DESC_F_XID_3_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h28
`define RD_RESP_DESC_F_XUSER_0_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h2C
`define RD_RESP_DESC_F_XUSER_1_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h30
`define RD_RESP_DESC_F_XUSER_2_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h34
`define RD_RESP_DESC_F_XUSER_3_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h38
`define RD_RESP_DESC_F_XUSER_4_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h3C
`define RD_RESP_DESC_F_XUSER_5_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h40
`define RD_RESP_DESC_F_XUSER_6_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h44
`define RD_RESP_DESC_F_XUSER_7_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h48
`define RD_RESP_DESC_F_XUSER_8_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h4C
`define RD_RESP_DESC_F_XUSER_9_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h50
`define RD_RESP_DESC_F_XUSER_10_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h54
`define RD_RESP_DESC_F_XUSER_11_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h58
`define RD_RESP_DESC_F_XUSER_12_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h5C
`define RD_RESP_DESC_F_XUSER_13_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h60
`define RD_RESP_DESC_F_XUSER_14_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h64
`define RD_RESP_DESC_F_XUSER_15_REG_ADDR `RD_RESP_DESC_F_BASE_ADDR + 'h68
`define WR_REQ_DESC_F_TXN_TYPE_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h0
`define WR_REQ_DESC_F_SIZE_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h4
`define WR_REQ_DESC_F_DATA_OFFSET_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h8
`define WR_REQ_DESC_F_DATA_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hC
`define WR_REQ_DESC_F_DATA_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h10
`define WR_REQ_DESC_F_DATA_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h14
`define WR_REQ_DESC_F_DATA_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h18
`define WR_REQ_DESC_F_WSTRB_HOST_ADDR_0_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h1C
`define WR_REQ_DESC_F_WSTRB_HOST_ADDR_1_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h20
`define WR_REQ_DESC_F_WSTRB_HOST_ADDR_2_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h24
`define WR_REQ_DESC_F_WSTRB_HOST_ADDR_3_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h28
`define WR_REQ_DESC_F_AXSIZE_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h2C
`define WR_REQ_DESC_F_ATTR_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h30
`define WR_REQ_DESC_F_AXADDR_0_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h34
`define WR_REQ_DESC_F_AXADDR_1_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h38
`define WR_REQ_DESC_F_AXADDR_2_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h3C
`define WR_REQ_DESC_F_AXADDR_3_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h40
`define WR_REQ_DESC_F_AXID_0_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h44
`define WR_REQ_DESC_F_AXID_1_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h48
`define WR_REQ_DESC_F_AXID_2_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h4C
`define WR_REQ_DESC_F_AXID_3_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h50
`define WR_REQ_DESC_F_AXUSER_0_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h54
`define WR_REQ_DESC_F_AXUSER_1_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h58
`define WR_REQ_DESC_F_AXUSER_2_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h5C
`define WR_REQ_DESC_F_AXUSER_3_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h60
`define WR_REQ_DESC_F_AXUSER_4_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h64
`define WR_REQ_DESC_F_AXUSER_5_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h68
`define WR_REQ_DESC_F_AXUSER_6_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h6C
`define WR_REQ_DESC_F_AXUSER_7_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h70
`define WR_REQ_DESC_F_AXUSER_8_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h74
`define WR_REQ_DESC_F_AXUSER_9_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h78
`define WR_REQ_DESC_F_AXUSER_10_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h7C
`define WR_REQ_DESC_F_AXUSER_11_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h80
`define WR_REQ_DESC_F_AXUSER_12_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h84
`define WR_REQ_DESC_F_AXUSER_13_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h88
`define WR_REQ_DESC_F_AXUSER_14_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h8C
`define WR_REQ_DESC_F_AXUSER_15_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h90
`define WR_REQ_DESC_F_WUSER_0_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h94
`define WR_REQ_DESC_F_WUSER_1_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h98
`define WR_REQ_DESC_F_WUSER_2_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'h9C
`define WR_REQ_DESC_F_WUSER_3_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hA0
`define WR_REQ_DESC_F_WUSER_4_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hA4
`define WR_REQ_DESC_F_WUSER_5_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hA8
`define WR_REQ_DESC_F_WUSER_6_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hAC
`define WR_REQ_DESC_F_WUSER_7_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hB0
`define WR_REQ_DESC_F_WUSER_8_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hB4
`define WR_REQ_DESC_F_WUSER_9_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hB8
`define WR_REQ_DESC_F_WUSER_10_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hBC
`define WR_REQ_DESC_F_WUSER_11_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hC0
`define WR_REQ_DESC_F_WUSER_12_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hC4
`define WR_REQ_DESC_F_WUSER_13_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hC8
`define WR_REQ_DESC_F_WUSER_14_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hCC
`define WR_REQ_DESC_F_WUSER_15_REG_ADDR `WR_REQ_DESC_F_BASE_ADDR + 'hD0
`define WR_RESP_DESC_F_RESP_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h0
`define WR_RESP_DESC_F_XID_0_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h4
`define WR_RESP_DESC_F_XID_1_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h8
`define WR_RESP_DESC_F_XID_2_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'hC
`define WR_RESP_DESC_F_XID_3_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h10
`define WR_RESP_DESC_F_XUSER_0_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h14
`define WR_RESP_DESC_F_XUSER_1_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h18
`define WR_RESP_DESC_F_XUSER_2_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h1C
`define WR_RESP_DESC_F_XUSER_3_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h20
`define WR_RESP_DESC_F_XUSER_4_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h24
`define WR_RESP_DESC_F_XUSER_5_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h28
`define WR_RESP_DESC_F_XUSER_6_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h2C
`define WR_RESP_DESC_F_XUSER_7_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h30
`define WR_RESP_DESC_F_XUSER_8_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h34
`define WR_RESP_DESC_F_XUSER_9_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h38
`define WR_RESP_DESC_F_XUSER_10_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h3C
`define WR_RESP_DESC_F_XUSER_11_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h40
`define WR_RESP_DESC_F_XUSER_12_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h44
`define WR_RESP_DESC_F_XUSER_13_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h48
`define WR_RESP_DESC_F_XUSER_14_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h4C
`define WR_RESP_DESC_F_XUSER_15_REG_ADDR `WR_RESP_DESC_F_BASE_ADDR + 'h50
`define SN_REQ_DESC_F_ATTR_REG_ADDR `SN_REQ_DESC_F_BASE_ADDR + 'h0
`define SN_REQ_DESC_F_ACADDR_0_REG_ADDR `SN_REQ_DESC_F_BASE_ADDR + 'h4
`define SN_REQ_DESC_F_ACADDR_1_REG_ADDR `SN_REQ_DESC_F_BASE_ADDR + 'h8
`define SN_REQ_DESC_F_ACADDR_2_REG_ADDR `SN_REQ_DESC_F_BASE_ADDR + 'hC
`define SN_REQ_DESC_F_ACADDR_3_REG_ADDR `SN_REQ_DESC_F_BASE_ADDR + 'h10
`define SN_RESP_DESC_F_RESP_REG_ADDR `SN_RESP_DESC_F_BASE_ADDR + 'h0


`define RDATA_RAM_REG_ADDR 'h8000
`define WDATA_RAM_REG_ADDR 'hC000
`define WSTRB_RAM_REG_ADDR 'h10000
`define CDDATA_RAM_REG_ADDR 'h14000

