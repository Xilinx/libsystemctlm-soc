/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Alok Mistry.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 *
 * Description: 
 * Converting all regsters in to 2D.
 *
 *
 */

reg [0:0] int_reg_desc_n_txn_type_wr_strb [MAX_DESC-1:0] ;
reg [0:0] int_reg_desc_n_txn_type_wr_rd [MAX_DESC-1:0] ;
reg [3:0] int_reg_desc_n_attr_axregion [MAX_DESC-1:0] ;
reg [3:0] int_reg_desc_n_attr_axqos [MAX_DESC-1:0] ;
reg [2:0] int_reg_desc_n_attr_axprot [MAX_DESC-1:0] ;
reg [3:0] int_reg_desc_n_attr_axcache [MAX_DESC-1:0] ;
reg [1:0] int_reg_desc_n_attr_axlock [MAX_DESC-1:0] ;
reg [1:0] int_reg_desc_n_attr_axburst [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axid_0_axid [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axid_1_axid [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axid_2_axid [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axid_3_axid [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_0_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_1_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_2_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_3_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_4_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_5_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_6_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_7_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_8_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_9_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_10_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_11_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_12_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_13_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_14_axuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axuser_15_axuser [MAX_DESC-1:0] ;
reg [15:0] int_reg_desc_n_size_txn_size [MAX_DESC-1:0] ;
reg [2:0] int_reg_desc_n_axsize_axsize [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axaddr_0_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axaddr_1_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axaddr_2_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_axaddr_3_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_data_offset_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_0_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_1_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_2_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_3_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_4_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_5_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_6_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_7_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_8_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_9_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_10_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_11_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_12_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_13_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_14_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wuser_15_wuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_data_host_addr_0_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_data_host_addr_1_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_data_host_addr_2_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_data_host_addr_3_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wstrb_host_addr_0_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wstrb_host_addr_1_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wstrb_host_addr_2_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_wstrb_host_addr_3_addr [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_0_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_1_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_2_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_3_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_4_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_5_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_6_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_7_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_8_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_9_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_10_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_11_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_12_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_13_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_14_xuser [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_15_xuser [MAX_DESC-1:0] ;

//we

reg [31:0] int_reg_desc_n_xuser_0_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_1_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_2_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_3_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_4_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_5_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_6_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_7_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_8_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_9_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_10_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_11_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_12_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_13_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_14_xuser_we [MAX_DESC-1:0] ;
reg [31:0] int_reg_desc_n_xuser_15_xuser_we [MAX_DESC-1:0] ;




wire [0:0] int_wire_desc_n_txn_type_wr_strb [MAX_DESC-1:0] ;
wire [MAX_DESC-1:0] int_wire_desc_n_txn_type_wr_rd ;
wire [3:0] int_wire_desc_n_attr_axregion [MAX_DESC-1:0] ;
wire [3:0] int_wire_desc_n_attr_axqos [MAX_DESC-1:0] ;
wire [2:0] int_wire_desc_n_attr_axprot [MAX_DESC-1:0] ;
wire [3:0] int_wire_desc_n_attr_axcache [MAX_DESC-1:0] ;
wire [1:0] int_wire_desc_n_attr_axlock [MAX_DESC-1:0] ;
wire [1:0] int_wire_desc_n_attr_axburst [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axid_0_axid [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axid_1_axid [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axid_2_axid [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axid_3_axid [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_0_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_1_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_2_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_3_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_4_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_5_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_6_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_7_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_8_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_9_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_10_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_11_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_12_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_13_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_14_axuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axuser_15_axuser [MAX_DESC-1:0] ;
wire [15:0] int_wire_desc_n_size_txn_size [MAX_DESC-1:0] ;
wire [2:0] int_wire_desc_n_axsize_axsize [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axaddr_0_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axaddr_1_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axaddr_2_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_axaddr_3_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_data_offset_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_0_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_1_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_2_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_3_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_4_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_5_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_6_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_7_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_8_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_9_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_10_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_11_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_12_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_13_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_14_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wuser_15_wuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_data_host_addr_0_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_data_host_addr_1_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_data_host_addr_2_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_data_host_addr_3_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wstrb_host_addr_0_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wstrb_host_addr_1_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wstrb_host_addr_2_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_wstrb_host_addr_3_addr [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_0_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_1_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_2_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_3_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_4_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_5_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_6_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_7_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_8_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_9_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_10_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_11_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_12_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_13_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_14_xuser [MAX_DESC-1:0] ;
wire [31:0] int_wire_desc_n_xuser_15_xuser [MAX_DESC-1:0] ;




genvar i; 


//Concatinating 128 bits of ID/Address.
wire [127:0] int_desc_n_axid_reg[MAX_DESC-1:0];
wire [127:0] int_desc_n_axaddr_reg[MAX_DESC-1:0];

wire [511:0] int_wire_desc_n_axuser[MAX_DESC-1:0];
wire [511:0] int_wire_desc_n_wuser[MAX_DESC-1:0];

// Combining axi ID & Address of 4 registers 
generate
 for (i=0;i<(MAX_DESC);i=i+1) 
 begin: gen_axid
 //Concate AXID of all Registers
 assign int_desc_n_axid_reg[i] = { int_wire_desc_n_axid_3_axid[i] ,int_wire_desc_n_axid_2_axid[i] 
 ,int_wire_desc_n_axid_1_axid[i] ,int_wire_desc_n_axid_0_axid[i]};
 assign int_desc_n_axaddr_reg[i] = { int_wire_desc_n_axaddr_3_addr[i] ,int_wire_desc_n_axaddr_2_addr[i] 
 ,int_wire_desc_n_axaddr_1_addr[i] ,int_wire_desc_n_axaddr_0_addr[i]};
 end
endgenerate

generate 
 for(i=0;i<MAX_DESC;i=i+1) begin:desc_axuser

 assign int_wire_desc_n_axuser[i]= {
 int_wire_desc_n_axuser_15_axuser[i],
 int_wire_desc_n_axuser_14_axuser[i],
 int_wire_desc_n_axuser_13_axuser[i],
 int_wire_desc_n_axuser_12_axuser[i],
 int_wire_desc_n_axuser_11_axuser[i],
 int_wire_desc_n_axuser_10_axuser[i],
 int_wire_desc_n_axuser_9_axuser [i],
 int_wire_desc_n_axuser_8_axuser [i],
 int_wire_desc_n_axuser_7_axuser [i],
 int_wire_desc_n_axuser_6_axuser [i],
 int_wire_desc_n_axuser_5_axuser [i],
 int_wire_desc_n_axuser_4_axuser [i],
 int_wire_desc_n_axuser_3_axuser [i],
 int_wire_desc_n_axuser_2_axuser [i],
 int_wire_desc_n_axuser_1_axuser [i],
 int_wire_desc_n_axuser_0_axuser [i]
 };


 assign int_wire_desc_n_wuser[i]= {
 int_wire_desc_n_wuser_15_wuser[i],
 int_wire_desc_n_wuser_14_wuser[i],
 int_wire_desc_n_wuser_13_wuser[i],
 int_wire_desc_n_wuser_12_wuser[i],
 int_wire_desc_n_wuser_11_wuser[i],
 int_wire_desc_n_wuser_10_wuser[i],
 int_wire_desc_n_wuser_9_wuser [i],
 int_wire_desc_n_wuser_8_wuser [i],
 int_wire_desc_n_wuser_7_wuser [i],
 int_wire_desc_n_wuser_6_wuser [i],
 int_wire_desc_n_wuser_5_wuser [i],
 int_wire_desc_n_wuser_4_wuser [i],
 int_wire_desc_n_wuser_3_wuser [i],
 int_wire_desc_n_wuser_2_wuser [i],
 int_wire_desc_n_wuser_1_wuser [i],
 int_wire_desc_n_wuser_0_wuser [i]
 };
 end
endgenerate





always@( posedge axi_aclk) 
 begin

 //for(i=0;i==0;i=i+1) begin:f1 
 int_reg_desc_n_txn_type_wr_strb [0] <= desc_0_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [0] <= desc_0_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [0] <= desc_0_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [0] <= desc_0_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [0] <= desc_0_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [0] <= desc_0_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [0] <= desc_0_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [0] <= desc_0_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [0] <= desc_0_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [0] <= desc_0_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [0] <= desc_0_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [0] <= desc_0_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [0] <= desc_0_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [0] <= desc_0_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [0] <= desc_0_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [0] <= desc_0_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [0] <= desc_0_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [0] <= desc_0_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [0] <= desc_0_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [0] <= desc_0_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [0] <= desc_0_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [0] <= desc_0_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [0] <= desc_0_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [0] <= desc_0_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [0] <= desc_0_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [0] <= desc_0_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [0] <= desc_0_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [0] <= desc_0_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [0] <= desc_0_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [0] <= desc_0_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [0] <= desc_0_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [0] <= desc_0_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [0] <= desc_0_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [0] <= desc_0_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [0] <= desc_0_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [0] <= desc_0_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [0] <= desc_0_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [0] <= desc_0_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [0] <= desc_0_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [0] <= desc_0_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [0] <= desc_0_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [0] <= desc_0_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [0] <= desc_0_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [0] <= desc_0_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [0] <= desc_0_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [0] <= desc_0_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [0] <= desc_0_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [0] <= desc_0_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [0] <= desc_0_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [0] <= desc_0_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [0] <= desc_0_wuser_15_reg ;
 //end

 int_reg_desc_n_txn_type_wr_strb [1] <= desc_1_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [1] <= desc_1_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [1] <= desc_1_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [1] <= desc_1_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [1] <= desc_1_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [1] <= desc_1_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [1] <= desc_1_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [1] <= desc_1_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [1] <= desc_1_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [1] <= desc_1_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [1] <= desc_1_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [1] <= desc_1_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [1] <= desc_1_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [1] <= desc_1_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [1] <= desc_1_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [1] <= desc_1_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [1] <= desc_1_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [1] <= desc_1_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [1] <= desc_1_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [1] <= desc_1_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [1] <= desc_1_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [1] <= desc_1_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [1] <= desc_1_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [1] <= desc_1_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [1] <= desc_1_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [1] <= desc_1_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [1] <= desc_1_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [1] <= desc_1_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [1] <= desc_1_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [1] <= desc_1_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [1] <= desc_1_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [1] <= desc_1_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [1] <= desc_1_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [1] <= desc_1_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [1] <= desc_1_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [1] <= desc_1_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [1] <= desc_1_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [1] <= desc_1_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [1] <= desc_1_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [1] <= desc_1_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [1] <= desc_1_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [1] <= desc_1_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [1] <= desc_1_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [1] <= desc_1_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [1] <= desc_1_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [1] <= desc_1_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [1] <= desc_1_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [1] <= desc_1_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [1] <= desc_1_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [1] <= desc_1_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [1] <= desc_1_wuser_15_reg ;




 int_reg_desc_n_txn_type_wr_strb [2] <= desc_2_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [2] <= desc_2_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [2] <= desc_2_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [2] <= desc_2_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [2] <= desc_2_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [2] <= desc_2_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [2] <= desc_2_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [2] <= desc_2_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [2] <= desc_2_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [2] <= desc_2_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [2] <= desc_2_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [2] <= desc_2_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [2] <= desc_2_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [2] <= desc_2_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [2] <= desc_2_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [2] <= desc_2_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [2] <= desc_2_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [2] <= desc_2_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [2] <= desc_2_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [2] <= desc_2_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [2] <= desc_2_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [2] <= desc_2_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [2] <= desc_2_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [2] <= desc_2_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [2] <= desc_2_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [2] <= desc_2_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [2] <= desc_2_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [2] <= desc_2_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [2] <= desc_2_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [2] <= desc_2_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [2] <= desc_2_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [2] <= desc_2_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [2] <= desc_2_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [2] <= desc_2_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [2] <= desc_2_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [2] <= desc_2_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [2] <= desc_2_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [2] <= desc_2_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [2] <= desc_2_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [2] <= desc_2_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [2] <= desc_2_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [2] <= desc_2_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [2] <= desc_2_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [2] <= desc_2_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [2] <= desc_2_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [2] <= desc_2_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [2] <= desc_2_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [2] <= desc_2_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [2] <= desc_2_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [2] <= desc_2_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [2] <= desc_2_wuser_15_reg ;









 int_reg_desc_n_txn_type_wr_strb [3] <= desc_3_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [3] <= desc_3_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [3] <= desc_3_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [3] <= desc_3_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [3] <= desc_3_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [3] <= desc_3_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [3] <= desc_3_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [3] <= desc_3_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [3] <= desc_3_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [3] <= desc_3_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [3] <= desc_3_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [3] <= desc_3_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [3] <= desc_3_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [3] <= desc_3_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [3] <= desc_3_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [3] <= desc_3_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [3] <= desc_3_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [3] <= desc_3_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [3] <= desc_3_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [3] <= desc_3_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [3] <= desc_3_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [3] <= desc_3_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [3] <= desc_3_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [3] <= desc_3_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [3] <= desc_3_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [3] <= desc_3_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [3] <= desc_3_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [3] <= desc_3_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [3] <= desc_3_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [3] <= desc_3_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [3] <= desc_3_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [3] <= desc_3_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [3] <= desc_3_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [3] <= desc_3_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [3] <= desc_3_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [3] <= desc_3_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [3] <= desc_3_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [3] <= desc_3_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [3] <= desc_3_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [3] <= desc_3_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [3] <= desc_3_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [3] <= desc_3_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [3] <= desc_3_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [3] <= desc_3_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [3] <= desc_3_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [3] <= desc_3_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [3] <= desc_3_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [3] <= desc_3_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [3] <= desc_3_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [3] <= desc_3_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [3] <= desc_3_wuser_15_reg ;




 int_reg_desc_n_txn_type_wr_strb [4] <= desc_4_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [4] <= desc_4_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [4] <= desc_4_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [4] <= desc_4_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [4] <= desc_4_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [4] <= desc_4_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [4] <= desc_4_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [4] <= desc_4_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [4] <= desc_4_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [4] <= desc_4_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [4] <= desc_4_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [4] <= desc_4_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [4] <= desc_4_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [4] <= desc_4_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [4] <= desc_4_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [4] <= desc_4_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [4] <= desc_4_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [4] <= desc_4_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [4] <= desc_4_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [4] <= desc_4_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [4] <= desc_4_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [4] <= desc_4_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [4] <= desc_4_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [4] <= desc_4_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [4] <= desc_4_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [4] <= desc_4_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [4] <= desc_4_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [4] <= desc_4_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [4] <= desc_4_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [4] <= desc_4_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [4] <= desc_4_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [4] <= desc_4_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [4] <= desc_4_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [4] <= desc_4_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [4] <= desc_4_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [4] <= desc_4_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [4] <= desc_4_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [4] <= desc_4_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [4] <= desc_4_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [4] <= desc_4_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [4] <= desc_4_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [4] <= desc_4_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [4] <= desc_4_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [4] <= desc_4_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [4] <= desc_4_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [4] <= desc_4_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [4] <= desc_4_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [4] <= desc_4_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [4] <= desc_4_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [4] <= desc_4_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [4] <= desc_4_wuser_15_reg ;





 int_reg_desc_n_txn_type_wr_strb [5] <= desc_5_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [5] <= desc_5_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [5] <= desc_5_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [5] <= desc_5_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [5] <= desc_5_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [5] <= desc_5_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [5] <= desc_5_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [5] <= desc_5_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [5] <= desc_5_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [5] <= desc_5_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [5] <= desc_5_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [5] <= desc_5_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [5] <= desc_5_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [5] <= desc_5_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [5] <= desc_5_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [5] <= desc_5_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [5] <= desc_5_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [5] <= desc_5_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [5] <= desc_5_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [5] <= desc_5_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [5] <= desc_5_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [5] <= desc_5_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [5] <= desc_5_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [5] <= desc_5_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [5] <= desc_5_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [5] <= desc_5_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [5] <= desc_5_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [5] <= desc_5_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [5] <= desc_5_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [5] <= desc_5_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [5] <= desc_5_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [5] <= desc_5_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [5] <= desc_5_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [5] <= desc_5_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [5] <= desc_5_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [5] <= desc_5_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [5] <= desc_5_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [5] <= desc_5_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [5] <= desc_5_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [5] <= desc_5_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [5] <= desc_5_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [5] <= desc_5_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [5] <= desc_5_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [5] <= desc_5_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [5] <= desc_5_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [5] <= desc_5_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [5] <= desc_5_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [5] <= desc_5_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [5] <= desc_5_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [5] <= desc_5_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [5] <= desc_5_wuser_15_reg ;






 int_reg_desc_n_txn_type_wr_strb [6] <= desc_6_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [6] <= desc_6_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [6] <= desc_6_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [6] <= desc_6_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [6] <= desc_6_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [6] <= desc_6_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [6] <= desc_6_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [6] <= desc_6_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [6] <= desc_6_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [6] <= desc_6_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [6] <= desc_6_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [6] <= desc_6_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [6] <= desc_6_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [6] <= desc_6_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [6] <= desc_6_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [6] <= desc_6_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [6] <= desc_6_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [6] <= desc_6_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [6] <= desc_6_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [6] <= desc_6_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [6] <= desc_6_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [6] <= desc_6_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [6] <= desc_6_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [6] <= desc_6_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [6] <= desc_6_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [6] <= desc_6_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [6] <= desc_6_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [6] <= desc_6_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [6] <= desc_6_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [6] <= desc_6_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [6] <= desc_6_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [6] <= desc_6_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [6] <= desc_6_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [6] <= desc_6_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [6] <= desc_6_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [6] <= desc_6_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [6] <= desc_6_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [6] <= desc_6_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [6] <= desc_6_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [6] <= desc_6_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [6] <= desc_6_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [6] <= desc_6_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [6] <= desc_6_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [6] <= desc_6_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [6] <= desc_6_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [6] <= desc_6_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [6] <= desc_6_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [6] <= desc_6_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [6] <= desc_6_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [6] <= desc_6_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [6] <= desc_6_wuser_15_reg ;




 int_reg_desc_n_txn_type_wr_strb [7] <= desc_7_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [7] <= desc_7_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [7] <= desc_7_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [7] <= desc_7_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [7] <= desc_7_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [7] <= desc_7_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [7] <= desc_7_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [7] <= desc_7_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [7] <= desc_7_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [7] <= desc_7_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [7] <= desc_7_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [7] <= desc_7_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [7] <= desc_7_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [7] <= desc_7_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [7] <= desc_7_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [7] <= desc_7_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [7] <= desc_7_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [7] <= desc_7_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [7] <= desc_7_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [7] <= desc_7_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [7] <= desc_7_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [7] <= desc_7_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [7] <= desc_7_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [7] <= desc_7_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [7] <= desc_7_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [7] <= desc_7_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [7] <= desc_7_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [7] <= desc_7_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [7] <= desc_7_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [7] <= desc_7_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [7] <= desc_7_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [7] <= desc_7_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [7] <= desc_7_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [7] <= desc_7_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [7] <= desc_7_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [7] <= desc_7_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [7] <= desc_7_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [7] <= desc_7_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [7] <= desc_7_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [7] <= desc_7_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [7] <= desc_7_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [7] <= desc_7_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [7] <= desc_7_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [7] <= desc_7_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [7] <= desc_7_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [7] <= desc_7_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [7] <= desc_7_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [7] <= desc_7_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [7] <= desc_7_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [7] <= desc_7_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [7] <= desc_7_wuser_15_reg ;




 int_reg_desc_n_txn_type_wr_strb [8] <= desc_8_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [8] <= desc_8_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [8] <= desc_8_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [8] <= desc_8_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [8] <= desc_8_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [8] <= desc_8_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [8] <= desc_8_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [8] <= desc_8_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [8] <= desc_8_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [8] <= desc_8_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [8] <= desc_8_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [8] <= desc_8_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [8] <= desc_8_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [8] <= desc_8_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [8] <= desc_8_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [8] <= desc_8_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [8] <= desc_8_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [8] <= desc_8_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [8] <= desc_8_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [8] <= desc_8_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [8] <= desc_8_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [8] <= desc_8_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [8] <= desc_8_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [8] <= desc_8_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [8] <= desc_8_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [8] <= desc_8_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [8] <= desc_8_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [8] <= desc_8_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [8] <= desc_8_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [8] <= desc_8_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [8] <= desc_8_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [8] <= desc_8_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [8] <= desc_8_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [8] <= desc_8_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [8] <= desc_8_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [8] <= desc_8_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [8] <= desc_8_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [8] <= desc_8_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [8] <= desc_8_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [8] <= desc_8_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [8] <= desc_8_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [8] <= desc_8_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [8] <= desc_8_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [8] <= desc_8_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [8] <= desc_8_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [8] <= desc_8_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [8] <= desc_8_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [8] <= desc_8_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [8] <= desc_8_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [8] <= desc_8_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [8] <= desc_8_wuser_15_reg ;



 int_reg_desc_n_txn_type_wr_strb [9] <= desc_9_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [9] <= desc_9_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [9] <= desc_9_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [9] <= desc_9_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [9] <= desc_9_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [9] <= desc_9_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [9] <= desc_9_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [9] <= desc_9_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [9] <= desc_9_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [9] <= desc_9_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [9] <= desc_9_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [9] <= desc_9_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [9] <= desc_9_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [9] <= desc_9_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [9] <= desc_9_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [9] <= desc_9_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [9] <= desc_9_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [9] <= desc_9_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [9] <= desc_9_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [9] <= desc_9_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [9] <= desc_9_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [9] <= desc_9_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [9] <= desc_9_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [9] <= desc_9_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [9] <= desc_9_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [9] <= desc_9_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [9] <= desc_9_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [9] <= desc_9_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [9] <= desc_9_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [9] <= desc_9_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [9] <= desc_9_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [9] <= desc_9_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [9] <= desc_9_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [9] <= desc_9_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [9] <= desc_9_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [9] <= desc_9_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [9] <= desc_9_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [9] <= desc_9_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [9] <= desc_9_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [9] <= desc_9_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [9] <= desc_9_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [9] <= desc_9_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [9] <= desc_9_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [9] <= desc_9_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [9] <= desc_9_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [9] <= desc_9_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [9] <= desc_9_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [9] <= desc_9_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [9] <= desc_9_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [9] <= desc_9_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [9] <= desc_9_wuser_15_reg ;


 
 int_reg_desc_n_txn_type_wr_strb [10] <= desc_10_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [10] <= desc_10_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [10] <= desc_10_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [10] <= desc_10_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [10] <= desc_10_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [10] <= desc_10_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [10] <= desc_10_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [10] <= desc_10_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [10] <= desc_10_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [10] <= desc_10_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [10] <= desc_10_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [10] <= desc_10_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [10] <= desc_10_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [10] <= desc_10_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [10] <= desc_10_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [10] <= desc_10_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [10] <= desc_10_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [10] <= desc_10_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [10] <= desc_10_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [10] <= desc_10_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [10] <= desc_10_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [10] <= desc_10_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [10] <= desc_10_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [10] <= desc_10_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [10] <= desc_10_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [10] <= desc_10_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [10] <= desc_10_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [10] <= desc_10_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [10] <= desc_10_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [10] <= desc_10_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [10] <= desc_10_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [10] <= desc_10_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [10] <= desc_10_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [10] <= desc_10_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [10] <= desc_10_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [10] <= desc_10_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [10] <= desc_10_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [10] <= desc_10_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [10] <= desc_10_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [10] <= desc_10_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [10] <= desc_10_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [10] <= desc_10_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [10] <= desc_10_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [10] <= desc_10_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [10] <= desc_10_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [10] <= desc_10_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [10] <= desc_10_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [10] <= desc_10_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [10] <= desc_10_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [10] <= desc_10_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [10] <= desc_10_wuser_15_reg ;
 

 int_reg_desc_n_txn_type_wr_strb [11] <= desc_11_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [11] <= desc_11_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [11] <= desc_11_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [11] <= desc_11_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [11] <= desc_11_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [11] <= desc_11_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [11] <= desc_11_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [11] <= desc_11_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [11] <= desc_11_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [11] <= desc_11_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [11] <= desc_11_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [11] <= desc_11_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [11] <= desc_11_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [11] <= desc_11_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [11] <= desc_11_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [11] <= desc_11_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [11] <= desc_11_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [11] <= desc_11_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [11] <= desc_11_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [11] <= desc_11_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [11] <= desc_11_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [11] <= desc_11_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [11] <= desc_11_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [11] <= desc_11_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [11] <= desc_11_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [11] <= desc_11_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [11] <= desc_11_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [11] <= desc_11_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [11] <= desc_11_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [11] <= desc_11_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [11] <= desc_11_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [11] <= desc_11_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [11] <= desc_11_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [11] <= desc_11_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [11] <= desc_11_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [11] <= desc_11_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [11] <= desc_11_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [11] <= desc_11_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [11] <= desc_11_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [11] <= desc_11_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [11] <= desc_11_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [11] <= desc_11_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [11] <= desc_11_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [11] <= desc_11_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [11] <= desc_11_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [11] <= desc_11_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [11] <= desc_11_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [11] <= desc_11_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [11] <= desc_11_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [11] <= desc_11_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [11] <= desc_11_wuser_15_reg ;



 int_reg_desc_n_txn_type_wr_strb [12] <= desc_12_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [12] <= desc_12_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [12] <= desc_12_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [12] <= desc_12_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [12] <= desc_12_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [12] <= desc_12_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [12] <= desc_12_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [12] <= desc_12_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [12] <= desc_12_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [12] <= desc_12_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [12] <= desc_12_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [12] <= desc_12_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [12] <= desc_12_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [12] <= desc_12_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [12] <= desc_12_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [12] <= desc_12_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [12] <= desc_12_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [12] <= desc_12_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [12] <= desc_12_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [12] <= desc_12_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [12] <= desc_12_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [12] <= desc_12_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [12] <= desc_12_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [12] <= desc_12_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [12] <= desc_12_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [12] <= desc_12_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [12] <= desc_12_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [12] <= desc_12_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [12] <= desc_12_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [12] <= desc_12_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [12] <= desc_12_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [12] <= desc_12_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [12] <= desc_12_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [12] <= desc_12_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [12] <= desc_12_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [12] <= desc_12_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [12] <= desc_12_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [12] <= desc_12_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [12] <= desc_12_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [12] <= desc_12_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [12] <= desc_12_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [12] <= desc_12_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [12] <= desc_12_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [12] <= desc_12_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [12] <= desc_12_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [12] <= desc_12_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [12] <= desc_12_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [12] <= desc_12_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [12] <= desc_12_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [12] <= desc_12_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [12] <= desc_12_wuser_15_reg ;


 int_reg_desc_n_txn_type_wr_strb [13] <= desc_13_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [13] <= desc_13_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [13] <= desc_13_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [13] <= desc_13_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [13] <= desc_13_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [13] <= desc_13_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [13] <= desc_13_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [13] <= desc_13_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [13] <= desc_13_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [13] <= desc_13_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [13] <= desc_13_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [13] <= desc_13_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [13] <= desc_13_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [13] <= desc_13_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [13] <= desc_13_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [13] <= desc_13_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [13] <= desc_13_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [13] <= desc_13_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [13] <= desc_13_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [13] <= desc_13_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [13] <= desc_13_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [13] <= desc_13_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [13] <= desc_13_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [13] <= desc_13_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [13] <= desc_13_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [13] <= desc_13_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [13] <= desc_13_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [13] <= desc_13_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [13] <= desc_13_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [13] <= desc_13_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [13] <= desc_13_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [13] <= desc_13_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [13] <= desc_13_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [13] <= desc_13_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [13] <= desc_13_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [13] <= desc_13_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [13] <= desc_13_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [13] <= desc_13_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [13] <= desc_13_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [13] <= desc_13_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [13] <= desc_13_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [13] <= desc_13_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [13] <= desc_13_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [13] <= desc_13_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [13] <= desc_13_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [13] <= desc_13_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [13] <= desc_13_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [13] <= desc_13_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [13] <= desc_13_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [13] <= desc_13_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [13] <= desc_13_wuser_15_reg ;




 int_reg_desc_n_txn_type_wr_strb [14] <= desc_14_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [14] <= desc_14_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [14] <= desc_14_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [14] <= desc_14_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [14] <= desc_14_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [14] <= desc_14_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [14] <= desc_14_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [14] <= desc_14_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [14] <= desc_14_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [14] <= desc_14_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [14] <= desc_14_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [14] <= desc_14_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [14] <= desc_14_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [14] <= desc_14_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [14] <= desc_14_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [14] <= desc_14_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [14] <= desc_14_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [14] <= desc_14_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [14] <= desc_14_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [14] <= desc_14_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [14] <= desc_14_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [14] <= desc_14_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [14] <= desc_14_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [14] <= desc_14_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [14] <= desc_14_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [14] <= desc_14_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [14] <= desc_14_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [14] <= desc_14_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [14] <= desc_14_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [14] <= desc_14_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [14] <= desc_14_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [14] <= desc_14_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [14] <= desc_14_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [14] <= desc_14_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [14] <= desc_14_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [14] <= desc_14_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [14] <= desc_14_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [14] <= desc_14_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [14] <= desc_14_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [14] <= desc_14_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [14] <= desc_14_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [14] <= desc_14_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [14] <= desc_14_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [14] <= desc_14_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [14] <= desc_14_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [14] <= desc_14_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [14] <= desc_14_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [14] <= desc_14_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [14] <= desc_14_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [14] <= desc_14_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [14] <= desc_14_wuser_15_reg ;




 int_reg_desc_n_txn_type_wr_strb [15] <= desc_15_txn_type_reg[1] ;
 int_reg_desc_n_txn_type_wr_rd [15] <= desc_15_txn_type_reg[0] ;
 int_reg_desc_n_attr_axregion [15] <= desc_15_attr_reg[18:15] ;
 int_reg_desc_n_attr_axqos [15] <= desc_15_attr_reg[14:11] ;
 int_reg_desc_n_attr_axprot [15] <= desc_15_attr_reg[10:8] ;
 int_reg_desc_n_attr_axcache [15] <= desc_15_attr_reg[7:4] ;
 int_reg_desc_n_attr_axlock [15] <= desc_15_attr_reg[3:2] ;
 int_reg_desc_n_attr_axburst [15] <= desc_15_attr_reg[1:0] ;
 int_reg_desc_n_axid_0_axid [15] <= desc_15_axid_0_reg ;
 int_reg_desc_n_axid_1_axid [15] <= desc_15_axid_1_reg ;
 int_reg_desc_n_axid_2_axid [15] <= desc_15_axid_2_reg ;
 int_reg_desc_n_axid_3_axid [15] <= desc_15_axid_3_reg ;
 int_reg_desc_n_axuser_0_axuser [15] <= desc_15_axuser_0_reg ;
 int_reg_desc_n_axuser_1_axuser [15] <= desc_15_axuser_1_reg ;
 int_reg_desc_n_axuser_2_axuser [15] <= desc_15_axuser_2_reg ;
 int_reg_desc_n_axuser_3_axuser [15] <= desc_15_axuser_3_reg ;
 int_reg_desc_n_axuser_4_axuser [15] <= desc_15_axuser_4_reg ;
 int_reg_desc_n_axuser_5_axuser [15] <= desc_15_axuser_5_reg ;
 int_reg_desc_n_axuser_6_axuser [15] <= desc_15_axuser_6_reg ;
 int_reg_desc_n_axuser_7_axuser [15] <= desc_15_axuser_7_reg ;
 int_reg_desc_n_axuser_8_axuser [15] <= desc_15_axuser_8_reg ;
 int_reg_desc_n_axuser_9_axuser [15] <= desc_15_axuser_9_reg ;
 int_reg_desc_n_axuser_10_axuser [15] <= desc_15_axuser_10_reg ;
 int_reg_desc_n_axuser_11_axuser [15] <= desc_15_axuser_11_reg ;
 int_reg_desc_n_axuser_12_axuser [15] <= desc_15_axuser_12_reg ;
 int_reg_desc_n_axuser_13_axuser [15] <= desc_15_axuser_13_reg ;
 int_reg_desc_n_axuser_14_axuser [15] <= desc_15_axuser_14_reg ;
 int_reg_desc_n_axuser_15_axuser [15] <= desc_15_axuser_15_reg ;
 int_reg_desc_n_size_txn_size [15] <= desc_15_size_reg[15:0] ;
 int_reg_desc_n_axsize_axsize [15] <= desc_15_axsize_reg[2:0] ;
 int_reg_desc_n_axaddr_0_addr [15] <= desc_15_axaddr_0_reg ;
 int_reg_desc_n_axaddr_1_addr [15] <= desc_15_axaddr_1_reg ;
 int_reg_desc_n_axaddr_2_addr [15] <= desc_15_axaddr_2_reg ;
 int_reg_desc_n_axaddr_3_addr [15] <= desc_15_axaddr_3_reg ;
 int_reg_desc_n_data_offset_addr [15] <= desc_15_data_offset_reg ;
 int_reg_desc_n_wuser_0_wuser [15] <= desc_15_wuser_0_reg ;
 int_reg_desc_n_wuser_1_wuser [15] <= desc_15_wuser_1_reg ;
 int_reg_desc_n_wuser_2_wuser [15] <= desc_15_wuser_2_reg ;
 int_reg_desc_n_wuser_3_wuser [15] <= desc_15_wuser_3_reg ;
 int_reg_desc_n_wuser_4_wuser [15] <= desc_15_wuser_4_reg ;
 int_reg_desc_n_wuser_5_wuser [15] <= desc_15_wuser_5_reg ;
 int_reg_desc_n_wuser_6_wuser [15] <= desc_15_wuser_6_reg ;
 int_reg_desc_n_wuser_7_wuser [15] <= desc_15_wuser_7_reg ;
 int_reg_desc_n_wuser_8_wuser [15] <= desc_15_wuser_8_reg ;
 int_reg_desc_n_wuser_9_wuser [15] <= desc_15_wuser_9_reg ;
 int_reg_desc_n_wuser_10_wuser [15] <= desc_15_wuser_10_reg ;
 int_reg_desc_n_wuser_11_wuser [15] <= desc_15_wuser_11_reg ;
 int_reg_desc_n_wuser_12_wuser [15] <= desc_15_wuser_12_reg ;
 int_reg_desc_n_wuser_13_wuser [15] <= desc_15_wuser_13_reg ;
 int_reg_desc_n_wuser_14_wuser [15] <= desc_15_wuser_14_reg ;
 int_reg_desc_n_wuser_15_wuser [15] <= desc_15_wuser_15_reg ;





 int_reg_desc_n_data_host_addr_0_addr [0] <= desc_0_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr [0] <= desc_0_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr [0] <= desc_0_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr [0] <= desc_0_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[0] <= desc_0_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[0] <= desc_0_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[0] <= desc_0_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[0] <= desc_0_wstrb_host_addr_3_reg ;


 int_reg_desc_n_data_host_addr_0_addr[1] <= desc_1_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[1] <= desc_1_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[1] <= desc_1_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[1] <= desc_1_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[1] <= desc_1_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[1] <= desc_1_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[1] <= desc_1_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[1] <= desc_1_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[2] <= desc_2_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[2] <= desc_2_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[2] <= desc_2_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[2] <= desc_2_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[2] <= desc_2_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[2] <= desc_2_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[2] <= desc_2_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[2] <= desc_2_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[3] <= desc_3_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[3] <= desc_3_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[3] <= desc_3_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[3] <= desc_3_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[3] <= desc_3_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[3] <= desc_3_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[3] <= desc_3_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[3] <= desc_3_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[4] <= desc_4_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[4] <= desc_4_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[4] <= desc_4_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[4] <= desc_4_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[4] <= desc_4_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[4] <= desc_4_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[4] <= desc_4_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[4] <= desc_4_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[5] <= desc_5_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[5] <= desc_5_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[5] <= desc_5_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[5] <= desc_5_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[5] <= desc_5_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[5] <= desc_5_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[5] <= desc_5_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[5] <= desc_5_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[6] <= desc_6_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[6] <= desc_6_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[6] <= desc_6_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[6] <= desc_6_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[6] <= desc_6_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[6] <= desc_6_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[6] <= desc_6_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[6] <= desc_6_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[7] <= desc_7_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[7] <= desc_7_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[7] <= desc_7_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[7] <= desc_7_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[7] <= desc_7_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[7] <= desc_7_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[7] <= desc_7_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[7] <= desc_7_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[8] <= desc_8_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[8] <= desc_8_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[8] <= desc_8_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[8] <= desc_8_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[8] <= desc_8_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[8] <= desc_8_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[8] <= desc_8_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[8] <= desc_8_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[9] <= desc_9_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[9] <= desc_9_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[9] <= desc_9_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[9] <= desc_9_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[9] <= desc_9_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[9] <= desc_9_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[9] <= desc_9_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[9] <= desc_9_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[10] <= desc_10_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[10] <= desc_10_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[10] <= desc_10_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[10] <= desc_10_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[10] <= desc_10_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[10] <= desc_10_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[10] <= desc_10_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[10] <= desc_10_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[11] <= desc_11_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[11] <= desc_11_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[11] <= desc_11_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[11] <= desc_11_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[11] <= desc_11_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[11] <= desc_11_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[11] <= desc_11_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[11] <= desc_11_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[12] <= desc_12_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[12] <= desc_12_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[12] <= desc_12_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[12] <= desc_12_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[12] <= desc_12_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[12] <= desc_12_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[12] <= desc_12_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[12] <= desc_12_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[13] <= desc_13_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[13] <= desc_13_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[13] <= desc_13_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[13] <= desc_13_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[13] <= desc_13_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[13] <= desc_13_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[13] <= desc_13_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[13] <= desc_13_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[14] <= desc_14_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[14] <= desc_14_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[14] <= desc_14_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[14] <= desc_14_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[14] <= desc_14_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[14] <= desc_14_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[14] <= desc_14_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[14] <= desc_14_wstrb_host_addr_3_reg ;
 int_reg_desc_n_data_host_addr_0_addr[15] <= desc_15_data_host_addr_0_reg ;
 int_reg_desc_n_data_host_addr_1_addr[15] <= desc_15_data_host_addr_1_reg ;
 int_reg_desc_n_data_host_addr_2_addr[15] <= desc_15_data_host_addr_2_reg ;
 int_reg_desc_n_data_host_addr_3_addr[15] <= desc_15_data_host_addr_3_reg ;
 int_reg_desc_n_wstrb_host_addr_0_addr[15] <= desc_15_wstrb_host_addr_0_reg ;
 int_reg_desc_n_wstrb_host_addr_1_addr[15] <= desc_15_wstrb_host_addr_1_reg ;
 int_reg_desc_n_wstrb_host_addr_2_addr[15] <= desc_15_wstrb_host_addr_2_reg ;
 int_reg_desc_n_wstrb_host_addr_3_addr[15] <= desc_15_wstrb_host_addr_3_reg ;

 end

//end//always
//xuser to be updated by user master
always@(posedge axi_aclk) begin
 uc2rb_desc_0_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[0] ; 
 uc2rb_desc_0_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[0] ;
 uc2rb_desc_0_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[0] ;
 uc2rb_desc_0_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[0] ;
 uc2rb_desc_0_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[0] ;
 uc2rb_desc_0_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[0] ;
 uc2rb_desc_0_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[0] ;
 uc2rb_desc_0_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[0] ;
 uc2rb_desc_0_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[0] ;
 uc2rb_desc_0_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[0] ;
 uc2rb_desc_0_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[0] ;
 uc2rb_desc_0_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[0] ;
 uc2rb_desc_0_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[0] ;
 uc2rb_desc_0_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[0] ;
 uc2rb_desc_0_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[0] ;
 uc2rb_desc_0_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[0] ;
 uc2rb_desc_1_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[1] ;
 uc2rb_desc_1_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[1] ;
 uc2rb_desc_1_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[1] ;
 uc2rb_desc_1_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[1] ;
 uc2rb_desc_1_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[1] ;
 uc2rb_desc_1_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[1] ;
 uc2rb_desc_1_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[1] ;
 uc2rb_desc_1_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[1] ;
 uc2rb_desc_1_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[1] ;
 uc2rb_desc_1_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[1] ;
 uc2rb_desc_1_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[1] ;
 uc2rb_desc_1_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[1] ;
 uc2rb_desc_1_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[1] ;
 uc2rb_desc_1_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[1] ;
 uc2rb_desc_1_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[1] ;
 uc2rb_desc_1_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[1] ;
 uc2rb_desc_2_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[2] ;
 uc2rb_desc_2_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[2] ;
 uc2rb_desc_2_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[2] ;
 uc2rb_desc_2_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[2] ;
 uc2rb_desc_2_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[2] ;
 uc2rb_desc_2_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[2] ;
 uc2rb_desc_2_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[2] ;
 uc2rb_desc_2_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[2] ;
 uc2rb_desc_2_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[2] ;
 uc2rb_desc_2_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[2] ;
 uc2rb_desc_2_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[2] ;
 uc2rb_desc_2_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[2] ;
 uc2rb_desc_2_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[2] ;
 uc2rb_desc_2_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[2] ;
 uc2rb_desc_2_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[2] ;
 uc2rb_desc_2_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[2] ;
 uc2rb_desc_3_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[3] ;
 uc2rb_desc_3_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[3] ;
 uc2rb_desc_3_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[3] ;
 uc2rb_desc_3_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[3] ;
 uc2rb_desc_3_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[3] ;
 uc2rb_desc_3_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[3] ;
 uc2rb_desc_3_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[3] ;
 uc2rb_desc_3_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[3] ;
 uc2rb_desc_3_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[3] ;
 uc2rb_desc_3_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[3] ;
 uc2rb_desc_3_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[3] ;
 uc2rb_desc_3_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[3] ;
 uc2rb_desc_3_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[3] ;
 uc2rb_desc_3_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[3] ;
 uc2rb_desc_3_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[3] ;
 uc2rb_desc_3_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[3] ;
 uc2rb_desc_4_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[4] ;
 uc2rb_desc_4_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[4] ;
 uc2rb_desc_4_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[4] ;
 uc2rb_desc_4_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[4] ;
 uc2rb_desc_4_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[4] ;
 uc2rb_desc_4_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[4] ;
 uc2rb_desc_4_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[4] ;
 uc2rb_desc_4_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[4] ;
 uc2rb_desc_4_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[4] ;
 uc2rb_desc_4_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[4] ;
 uc2rb_desc_4_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[4] ;
 uc2rb_desc_4_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[4] ;
 uc2rb_desc_4_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[4] ;
 uc2rb_desc_4_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[4] ;
 uc2rb_desc_4_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[4] ;
 uc2rb_desc_4_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[4] ;
 uc2rb_desc_5_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[5] ;
 uc2rb_desc_5_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[5] ;
 uc2rb_desc_5_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[5] ;
 uc2rb_desc_5_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[5] ;
 uc2rb_desc_5_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[5] ;
 uc2rb_desc_5_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[5] ;
 uc2rb_desc_5_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[5] ;
 uc2rb_desc_5_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[5] ;
 uc2rb_desc_5_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[5] ;
 uc2rb_desc_5_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[5] ;
 uc2rb_desc_5_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[5] ;
 uc2rb_desc_5_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[5] ;
 uc2rb_desc_5_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[5] ;
 uc2rb_desc_5_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[5] ;
 uc2rb_desc_5_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[5] ;
 uc2rb_desc_5_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[5] ;
 uc2rb_desc_6_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[6] ;
 uc2rb_desc_6_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[6] ;
 uc2rb_desc_6_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[6] ;
 uc2rb_desc_6_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[6] ;
 uc2rb_desc_6_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[6] ;
 uc2rb_desc_6_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[6] ;
 uc2rb_desc_6_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[6] ;
 uc2rb_desc_6_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[6] ;
 uc2rb_desc_6_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[6] ;
 uc2rb_desc_6_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[6] ;
 uc2rb_desc_6_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[6] ;
 uc2rb_desc_6_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[6] ;
 uc2rb_desc_6_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[6] ;
 uc2rb_desc_6_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[6] ;
 uc2rb_desc_6_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[6] ;
 uc2rb_desc_6_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[6] ;
 uc2rb_desc_7_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[7] ;
 uc2rb_desc_7_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[7] ;
 uc2rb_desc_7_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[7] ;
 uc2rb_desc_7_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[7] ;
 uc2rb_desc_7_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[7] ;
 uc2rb_desc_7_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[7] ;
 uc2rb_desc_7_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[7] ;
 uc2rb_desc_7_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[7] ;
 uc2rb_desc_7_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[7] ;
 uc2rb_desc_7_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[7] ;
 uc2rb_desc_7_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[7] ;
 uc2rb_desc_7_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[7] ;
 uc2rb_desc_7_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[7] ;
 uc2rb_desc_7_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[7] ;
 uc2rb_desc_7_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[7] ;
 uc2rb_desc_7_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[7] ;
 uc2rb_desc_8_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[8] ;
 uc2rb_desc_8_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[8] ;
 uc2rb_desc_8_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[8] ;
 uc2rb_desc_8_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[8] ;
 uc2rb_desc_8_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[8] ;
 uc2rb_desc_8_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[8] ;
 uc2rb_desc_8_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[8] ;
 uc2rb_desc_8_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[8] ;
 uc2rb_desc_8_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[8] ;
 uc2rb_desc_8_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[8] ;
 uc2rb_desc_8_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[8] ;
 uc2rb_desc_8_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[8] ;
 uc2rb_desc_8_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[8] ;
 uc2rb_desc_8_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[8] ;
 uc2rb_desc_8_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[8] ;
 uc2rb_desc_8_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[8] ;
 uc2rb_desc_9_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[9] ;
 uc2rb_desc_9_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[9] ;
 uc2rb_desc_9_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[9] ;
 uc2rb_desc_9_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[9] ;
 uc2rb_desc_9_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[9] ;
 uc2rb_desc_9_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[9] ;
 uc2rb_desc_9_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[9] ;
 uc2rb_desc_9_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[9] ;
 uc2rb_desc_9_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[9] ;
 uc2rb_desc_9_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[9] ;
 uc2rb_desc_9_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[9] ;
 uc2rb_desc_9_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[9] ;
 uc2rb_desc_9_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[9] ;
 uc2rb_desc_9_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[9] ;
 uc2rb_desc_9_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[9] ;
 uc2rb_desc_9_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[9] ;
 uc2rb_desc_10_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[10] ;
 uc2rb_desc_10_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[10] ;
 uc2rb_desc_10_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[10] ;
 uc2rb_desc_10_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[10] ;
 uc2rb_desc_10_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[10] ;
 uc2rb_desc_10_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[10] ;
 uc2rb_desc_10_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[10] ;
 uc2rb_desc_10_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[10] ;
 uc2rb_desc_10_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[10] ;
 uc2rb_desc_10_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[10] ;
 uc2rb_desc_10_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[10] ;
 uc2rb_desc_10_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[10] ;
 uc2rb_desc_10_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[10] ;
 uc2rb_desc_10_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[10] ;
 uc2rb_desc_10_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[10] ;
 uc2rb_desc_10_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[10] ;
 uc2rb_desc_11_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[11] ;
 uc2rb_desc_11_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[11] ;
 uc2rb_desc_11_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[11] ;
 uc2rb_desc_11_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[11] ;
 uc2rb_desc_11_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[11] ;
 uc2rb_desc_11_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[11] ;
 uc2rb_desc_11_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[11] ;
 uc2rb_desc_11_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[11] ;
 uc2rb_desc_11_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[11] ;
 uc2rb_desc_11_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[11] ;
 uc2rb_desc_11_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[11] ;
 uc2rb_desc_11_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[11] ;
 uc2rb_desc_11_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[11] ;
 uc2rb_desc_11_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[11] ;
 uc2rb_desc_11_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[11] ;
 uc2rb_desc_11_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[11] ;
 uc2rb_desc_12_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[12] ;
 uc2rb_desc_12_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[12] ;
 uc2rb_desc_12_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[12] ;
 uc2rb_desc_12_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[12] ;
 uc2rb_desc_12_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[12] ;
 uc2rb_desc_12_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[12] ;
 uc2rb_desc_12_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[12] ;
 uc2rb_desc_12_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[12] ;
 uc2rb_desc_12_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[12] ;
 uc2rb_desc_12_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[12] ;
 uc2rb_desc_12_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[12] ;
 uc2rb_desc_12_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[12] ;
 uc2rb_desc_12_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[12] ;
 uc2rb_desc_12_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[12] ;
 uc2rb_desc_12_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[12] ;
 uc2rb_desc_12_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[12] ;
 uc2rb_desc_13_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[13] ;
 uc2rb_desc_13_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[13] ;
 uc2rb_desc_13_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[13] ;
 uc2rb_desc_13_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[13] ;
 uc2rb_desc_13_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[13] ;
 uc2rb_desc_13_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[13] ;
 uc2rb_desc_13_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[13] ;
 uc2rb_desc_13_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[13] ;
 uc2rb_desc_13_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[13] ;
 uc2rb_desc_13_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[13] ;
 uc2rb_desc_13_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[13] ;
 uc2rb_desc_13_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[13] ;
 uc2rb_desc_13_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[13] ;
 uc2rb_desc_13_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[13] ;
 uc2rb_desc_13_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[13] ;
 uc2rb_desc_13_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[13] ;
 uc2rb_desc_14_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[14] ;
 uc2rb_desc_14_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[14] ;
 uc2rb_desc_14_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[14] ;
 uc2rb_desc_14_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[14] ;
 uc2rb_desc_14_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[14] ;
 uc2rb_desc_14_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[14] ;
 uc2rb_desc_14_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[14] ;
 uc2rb_desc_14_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[14] ;
 uc2rb_desc_14_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[14] ;
 uc2rb_desc_14_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[14] ;
 uc2rb_desc_14_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[14] ;
 uc2rb_desc_14_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[14] ;
 uc2rb_desc_14_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[14] ;
 uc2rb_desc_14_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[14] ;
 uc2rb_desc_14_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[14] ;
 uc2rb_desc_14_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[14] ;
 uc2rb_desc_15_xuser_0_reg <= int_reg_desc_n_xuser_0_xuser[15] ;
 uc2rb_desc_15_xuser_1_reg <= int_reg_desc_n_xuser_1_xuser[15] ;
 uc2rb_desc_15_xuser_2_reg <= int_reg_desc_n_xuser_2_xuser[15] ;
 uc2rb_desc_15_xuser_3_reg <= int_reg_desc_n_xuser_3_xuser[15] ;
 uc2rb_desc_15_xuser_4_reg <= int_reg_desc_n_xuser_4_xuser[15] ;
 uc2rb_desc_15_xuser_5_reg <= int_reg_desc_n_xuser_5_xuser[15] ;
 uc2rb_desc_15_xuser_6_reg <= int_reg_desc_n_xuser_6_xuser[15] ;
 uc2rb_desc_15_xuser_7_reg <= int_reg_desc_n_xuser_7_xuser[15] ;
 uc2rb_desc_15_xuser_8_reg <= int_reg_desc_n_xuser_8_xuser[15] ;
 uc2rb_desc_15_xuser_9_reg <= int_reg_desc_n_xuser_9_xuser[15] ;
 uc2rb_desc_15_xuser_10_reg <= int_reg_desc_n_xuser_10_xuser[15] ;
 uc2rb_desc_15_xuser_11_reg <= int_reg_desc_n_xuser_11_xuser[15] ;
 uc2rb_desc_15_xuser_12_reg <= int_reg_desc_n_xuser_12_xuser[15] ;
 uc2rb_desc_15_xuser_13_reg <= int_reg_desc_n_xuser_13_xuser[15] ;
 uc2rb_desc_15_xuser_14_reg <= int_reg_desc_n_xuser_14_xuser[15] ;
 uc2rb_desc_15_xuser_15_reg <= int_reg_desc_n_xuser_15_xuser[15] ;
end




always@(posedge axi_aclk) begin
 uc2rb_desc_0_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[0] ; 
 uc2rb_desc_0_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[0] ;
 uc2rb_desc_0_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[0] ;
 uc2rb_desc_0_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[0] ;
 uc2rb_desc_0_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[0] ;
 uc2rb_desc_0_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[0] ;
 uc2rb_desc_0_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[0] ;
 uc2rb_desc_0_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[0] ;
 uc2rb_desc_0_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[0] ;
 uc2rb_desc_0_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[0] ;
 uc2rb_desc_0_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[0] ;
 uc2rb_desc_0_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[0] ;
 uc2rb_desc_0_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[0] ;
 uc2rb_desc_0_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[0] ;
 uc2rb_desc_0_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[0] ;
 uc2rb_desc_0_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[0] ;
 uc2rb_desc_1_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[1] ;
 uc2rb_desc_1_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[1] ;
 uc2rb_desc_1_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[1] ;
 uc2rb_desc_1_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[1] ;
 uc2rb_desc_1_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[1] ;
 uc2rb_desc_1_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[1] ;
 uc2rb_desc_1_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[1] ;
 uc2rb_desc_1_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[1] ;
 uc2rb_desc_1_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[1] ;
 uc2rb_desc_1_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[1] ;
 uc2rb_desc_1_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[1] ;
 uc2rb_desc_1_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[1] ;
 uc2rb_desc_1_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[1] ;
 uc2rb_desc_1_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[1] ;
 uc2rb_desc_1_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[1] ;
 uc2rb_desc_1_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[1] ;
 uc2rb_desc_2_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[2] ;
 uc2rb_desc_2_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[2] ;
 uc2rb_desc_2_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[2] ;
 uc2rb_desc_2_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[2] ;
 uc2rb_desc_2_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[2] ;
 uc2rb_desc_2_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[2] ;
 uc2rb_desc_2_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[2] ;
 uc2rb_desc_2_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[2] ;
 uc2rb_desc_2_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[2] ;
 uc2rb_desc_2_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[2] ;
 uc2rb_desc_2_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[2] ;
 uc2rb_desc_2_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[2] ;
 uc2rb_desc_2_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[2] ;
 uc2rb_desc_2_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[2] ;
 uc2rb_desc_2_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[2] ;
 uc2rb_desc_2_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[2] ;
 uc2rb_desc_3_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[3] ;
 uc2rb_desc_3_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[3] ;
 uc2rb_desc_3_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[3] ;
 uc2rb_desc_3_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[3] ;
 uc2rb_desc_3_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[3] ;
 uc2rb_desc_3_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[3] ;
 uc2rb_desc_3_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[3] ;
 uc2rb_desc_3_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[3] ;
 uc2rb_desc_3_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[3] ;
 uc2rb_desc_3_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[3] ;
 uc2rb_desc_3_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[3] ;
 uc2rb_desc_3_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[3] ;
 uc2rb_desc_3_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[3] ;
 uc2rb_desc_3_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[3] ;
 uc2rb_desc_3_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[3] ;
 uc2rb_desc_3_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[3] ;
 uc2rb_desc_4_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[4] ;
 uc2rb_desc_4_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[4] ;
 uc2rb_desc_4_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[4] ;
 uc2rb_desc_4_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[4] ;
 uc2rb_desc_4_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[4] ;
 uc2rb_desc_4_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[4] ;
 uc2rb_desc_4_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[4] ;
 uc2rb_desc_4_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[4] ;
 uc2rb_desc_4_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[4] ;
 uc2rb_desc_4_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[4] ;
 uc2rb_desc_4_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[4] ;
 uc2rb_desc_4_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[4] ;
 uc2rb_desc_4_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[4] ;
 uc2rb_desc_4_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[4] ;
 uc2rb_desc_4_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[4] ;
 uc2rb_desc_4_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[4] ;
 uc2rb_desc_5_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[5] ;
 uc2rb_desc_5_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[5] ;
 uc2rb_desc_5_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[5] ;
 uc2rb_desc_5_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[5] ;
 uc2rb_desc_5_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[5] ;
 uc2rb_desc_5_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[5] ;
 uc2rb_desc_5_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[5] ;
 uc2rb_desc_5_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[5] ;
 uc2rb_desc_5_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[5] ;
 uc2rb_desc_5_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[5] ;
 uc2rb_desc_5_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[5] ;
 uc2rb_desc_5_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[5] ;
 uc2rb_desc_5_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[5] ;
 uc2rb_desc_5_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[5] ;
 uc2rb_desc_5_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[5] ;
 uc2rb_desc_5_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[5] ;
 uc2rb_desc_6_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[6] ;
 uc2rb_desc_6_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[6] ;
 uc2rb_desc_6_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[6] ;
 uc2rb_desc_6_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[6] ;
 uc2rb_desc_6_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[6] ;
 uc2rb_desc_6_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[6] ;
 uc2rb_desc_6_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[6] ;
 uc2rb_desc_6_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[6] ;
 uc2rb_desc_6_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[6] ;
 uc2rb_desc_6_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[6] ;
 uc2rb_desc_6_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[6] ;
 uc2rb_desc_6_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[6] ;
 uc2rb_desc_6_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[6] ;
 uc2rb_desc_6_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[6] ;
 uc2rb_desc_6_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[6] ;
 uc2rb_desc_6_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[6] ;
 uc2rb_desc_7_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[7] ;
 uc2rb_desc_7_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[7] ;
 uc2rb_desc_7_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[7] ;
 uc2rb_desc_7_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[7] ;
 uc2rb_desc_7_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[7] ;
 uc2rb_desc_7_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[7] ;
 uc2rb_desc_7_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[7] ;
 uc2rb_desc_7_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[7] ;
 uc2rb_desc_7_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[7] ;
 uc2rb_desc_7_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[7] ;
 uc2rb_desc_7_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[7] ;
 uc2rb_desc_7_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[7] ;
 uc2rb_desc_7_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[7] ;
 uc2rb_desc_7_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[7] ;
 uc2rb_desc_7_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[7] ;
 uc2rb_desc_7_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[7] ;
 uc2rb_desc_8_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[8] ;
 uc2rb_desc_8_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[8] ;
 uc2rb_desc_8_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[8] ;
 uc2rb_desc_8_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[8] ;
 uc2rb_desc_8_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[8] ;
 uc2rb_desc_8_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[8] ;
 uc2rb_desc_8_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[8] ;
 uc2rb_desc_8_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[8] ;
 uc2rb_desc_8_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[8] ;
 uc2rb_desc_8_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[8] ;
 uc2rb_desc_8_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[8] ;
 uc2rb_desc_8_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[8] ;
 uc2rb_desc_8_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[8] ;
 uc2rb_desc_8_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[8] ;
 uc2rb_desc_8_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[8] ;
 uc2rb_desc_8_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[8] ;
 uc2rb_desc_9_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[9] ;
 uc2rb_desc_9_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[9] ;
 uc2rb_desc_9_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[9] ;
 uc2rb_desc_9_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[9] ;
 uc2rb_desc_9_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[9] ;
 uc2rb_desc_9_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[9] ;
 uc2rb_desc_9_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[9] ;
 uc2rb_desc_9_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[9] ;
 uc2rb_desc_9_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[9] ;
 uc2rb_desc_9_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[9] ;
 uc2rb_desc_9_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[9] ;
 uc2rb_desc_9_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[9] ;
 uc2rb_desc_9_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[9] ;
 uc2rb_desc_9_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[9] ;
 uc2rb_desc_9_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[9] ;
 uc2rb_desc_9_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[9] ;
 uc2rb_desc_10_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[10] ;
 uc2rb_desc_10_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[10] ;
 uc2rb_desc_10_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[10] ;
 uc2rb_desc_10_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[10] ;
 uc2rb_desc_10_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[10] ;
 uc2rb_desc_10_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[10] ;
 uc2rb_desc_10_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[10] ;
 uc2rb_desc_10_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[10] ;
 uc2rb_desc_10_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[10] ;
 uc2rb_desc_10_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[10] ;
 uc2rb_desc_10_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[10] ;
 uc2rb_desc_10_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[10] ;
 uc2rb_desc_10_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[10] ;
 uc2rb_desc_10_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[10] ;
 uc2rb_desc_10_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[10] ;
 uc2rb_desc_10_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[10] ;
 uc2rb_desc_11_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[11] ;
 uc2rb_desc_11_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[11] ;
 uc2rb_desc_11_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[11] ;
 uc2rb_desc_11_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[11] ;
 uc2rb_desc_11_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[11] ;
 uc2rb_desc_11_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[11] ;
 uc2rb_desc_11_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[11] ;
 uc2rb_desc_11_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[11] ;
 uc2rb_desc_11_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[11] ;
 uc2rb_desc_11_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[11] ;
 uc2rb_desc_11_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[11] ;
 uc2rb_desc_11_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[11] ;
 uc2rb_desc_11_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[11] ;
 uc2rb_desc_11_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[11] ;
 uc2rb_desc_11_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[11] ;
 uc2rb_desc_11_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[11] ;
 uc2rb_desc_12_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[12] ;
 uc2rb_desc_12_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[12] ;
 uc2rb_desc_12_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[12] ;
 uc2rb_desc_12_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[12] ;
 uc2rb_desc_12_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[12] ;
 uc2rb_desc_12_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[12] ;
 uc2rb_desc_12_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[12] ;
 uc2rb_desc_12_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[12] ;
 uc2rb_desc_12_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[12] ;
 uc2rb_desc_12_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[12] ;
 uc2rb_desc_12_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[12] ;
 uc2rb_desc_12_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[12] ;
 uc2rb_desc_12_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[12] ;
 uc2rb_desc_12_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[12] ;
 uc2rb_desc_12_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[12] ;
 uc2rb_desc_12_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[12] ;
 uc2rb_desc_13_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[13] ;
 uc2rb_desc_13_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[13] ;
 uc2rb_desc_13_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[13] ;
 uc2rb_desc_13_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[13] ;
 uc2rb_desc_13_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[13] ;
 uc2rb_desc_13_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[13] ;
 uc2rb_desc_13_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[13] ;
 uc2rb_desc_13_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[13] ;
 uc2rb_desc_13_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[13] ;
 uc2rb_desc_13_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[13] ;
 uc2rb_desc_13_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[13] ;
 uc2rb_desc_13_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[13] ;
 uc2rb_desc_13_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[13] ;
 uc2rb_desc_13_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[13] ;
 uc2rb_desc_13_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[13] ;
 uc2rb_desc_13_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[13] ;
 uc2rb_desc_14_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[14] ;
 uc2rb_desc_14_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[14] ;
 uc2rb_desc_14_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[14] ;
 uc2rb_desc_14_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[14] ;
 uc2rb_desc_14_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[14] ;
 uc2rb_desc_14_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[14] ;
 uc2rb_desc_14_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[14] ;
 uc2rb_desc_14_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[14] ;
 uc2rb_desc_14_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[14] ;
 uc2rb_desc_14_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[14] ;
 uc2rb_desc_14_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[14] ;
 uc2rb_desc_14_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[14] ;
 uc2rb_desc_14_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[14] ;
 uc2rb_desc_14_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[14] ;
 uc2rb_desc_14_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[14] ;
 uc2rb_desc_14_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[14] ;
 uc2rb_desc_15_xuser_0_reg_we <= int_reg_desc_n_xuser_0_xuser_we[15] ;
 uc2rb_desc_15_xuser_1_reg_we <= int_reg_desc_n_xuser_1_xuser_we[15] ;
 uc2rb_desc_15_xuser_2_reg_we <= int_reg_desc_n_xuser_2_xuser_we[15] ;
 uc2rb_desc_15_xuser_3_reg_we <= int_reg_desc_n_xuser_3_xuser_we[15] ;
 uc2rb_desc_15_xuser_4_reg_we <= int_reg_desc_n_xuser_4_xuser_we[15] ;
 uc2rb_desc_15_xuser_5_reg_we <= int_reg_desc_n_xuser_5_xuser_we[15] ;
 uc2rb_desc_15_xuser_6_reg_we <= int_reg_desc_n_xuser_6_xuser_we[15] ;
 uc2rb_desc_15_xuser_7_reg_we <= int_reg_desc_n_xuser_7_xuser_we[15] ;
 uc2rb_desc_15_xuser_8_reg_we <= int_reg_desc_n_xuser_8_xuser_we[15] ;
 uc2rb_desc_15_xuser_9_reg_we <= int_reg_desc_n_xuser_9_xuser_we[15] ;
 uc2rb_desc_15_xuser_10_reg_we <= int_reg_desc_n_xuser_10_xuser_we[15] ;
 uc2rb_desc_15_xuser_11_reg_we <= int_reg_desc_n_xuser_11_xuser_we[15] ;
 uc2rb_desc_15_xuser_12_reg_we <= int_reg_desc_n_xuser_12_xuser_we[15] ;
 uc2rb_desc_15_xuser_13_reg_we <= int_reg_desc_n_xuser_13_xuser_we[15] ;
 uc2rb_desc_15_xuser_14_reg_we <= int_reg_desc_n_xuser_14_xuser_we[15] ;
 uc2rb_desc_15_xuser_15_reg_we <= int_reg_desc_n_xuser_15_xuser_we[15] ;
end

generate
 for(i=0;i<MAX_DESC;i=i+1) begin :reg_to_wire
 assign int_wire_desc_n_txn_type_wr_strb[i] = int_reg_desc_n_txn_type_wr_strb[i] ; 
 assign int_wire_desc_n_txn_type_wr_rd[i] = int_reg_desc_n_txn_type_wr_rd[i] ; 
 assign int_wire_desc_n_attr_axregion[i] = int_reg_desc_n_attr_axregion[i] ; 
 assign int_wire_desc_n_attr_axqos[i] = int_reg_desc_n_attr_axqos[i] ; 
 assign int_wire_desc_n_attr_axprot[i] = int_reg_desc_n_attr_axprot[i] ; 
 assign int_wire_desc_n_attr_axcache[i] = int_reg_desc_n_attr_axcache[i] ; 
 assign int_wire_desc_n_attr_axlock[i] = int_reg_desc_n_attr_axlock[i] ; 
 assign int_wire_desc_n_attr_axburst[i] = int_reg_desc_n_attr_axburst[i] ; 
 assign int_wire_desc_n_axid_0_axid[i] = int_reg_desc_n_axid_0_axid[i] ; 
 assign int_wire_desc_n_axid_1_axid[i] = int_reg_desc_n_axid_1_axid[i] ; 
 assign int_wire_desc_n_axid_2_axid[i] = int_reg_desc_n_axid_2_axid[i] ; 
 assign int_wire_desc_n_axid_3_axid[i] = int_reg_desc_n_axid_3_axid[i] ; 
 assign int_wire_desc_n_axuser_0_axuser[i] = int_reg_desc_n_axuser_0_axuser[i] ; 
 assign int_wire_desc_n_axuser_1_axuser[i] = int_reg_desc_n_axuser_1_axuser[i] ; 
 assign int_wire_desc_n_axuser_2_axuser[i] = int_reg_desc_n_axuser_2_axuser[i] ; 
 assign int_wire_desc_n_axuser_3_axuser[i] = int_reg_desc_n_axuser_3_axuser[i] ; 
 assign int_wire_desc_n_axuser_4_axuser[i] = int_reg_desc_n_axuser_4_axuser[i] ; 
 assign int_wire_desc_n_axuser_5_axuser[i] = int_reg_desc_n_axuser_5_axuser[i] ; 
 assign int_wire_desc_n_axuser_6_axuser[i] = int_reg_desc_n_axuser_6_axuser[i] ; 
 assign int_wire_desc_n_axuser_7_axuser[i] = int_reg_desc_n_axuser_7_axuser[i] ; 
 assign int_wire_desc_n_axuser_8_axuser[i] = int_reg_desc_n_axuser_8_axuser[i] ; 
 assign int_wire_desc_n_axuser_9_axuser[i] = int_reg_desc_n_axuser_9_axuser[i] ; 
 assign int_wire_desc_n_axuser_10_axuser[i] = int_reg_desc_n_axuser_10_axuser[i] ; 
 assign int_wire_desc_n_axuser_11_axuser[i] = int_reg_desc_n_axuser_11_axuser[i] ; 
 assign int_wire_desc_n_axuser_12_axuser[i] = int_reg_desc_n_axuser_12_axuser[i] ; 
 assign int_wire_desc_n_axuser_13_axuser[i] = int_reg_desc_n_axuser_13_axuser[i] ; 
 assign int_wire_desc_n_axuser_14_axuser[i] = int_reg_desc_n_axuser_14_axuser[i] ; 
 assign int_wire_desc_n_axuser_15_axuser[i] = int_reg_desc_n_axuser_15_axuser[i] ; 
 assign int_wire_desc_n_size_txn_size[i] = int_reg_desc_n_size_txn_size[i] ; 
 assign int_wire_desc_n_axsize_axsize[i] = int_reg_desc_n_axsize_axsize[i] ; 
 assign int_wire_desc_n_axaddr_0_addr[i] = int_reg_desc_n_axaddr_0_addr[i] ; 
 assign int_wire_desc_n_axaddr_1_addr[i] = int_reg_desc_n_axaddr_1_addr[i] ; 
 assign int_wire_desc_n_axaddr_2_addr[i] = int_reg_desc_n_axaddr_2_addr[i] ; 
 assign int_wire_desc_n_axaddr_3_addr[i] = int_reg_desc_n_axaddr_3_addr[i] ; 
 assign int_wire_desc_n_data_offset_addr[i] = int_reg_desc_n_data_offset_addr[i] ; 
 assign int_wire_desc_n_wuser_0_wuser[i] = int_reg_desc_n_wuser_0_wuser[i] ; 
 assign int_wire_desc_n_wuser_1_wuser[i] = int_reg_desc_n_wuser_1_wuser[i] ; 
 assign int_wire_desc_n_wuser_2_wuser[i] = int_reg_desc_n_wuser_2_wuser[i] ; 
 assign int_wire_desc_n_wuser_3_wuser[i] = int_reg_desc_n_wuser_3_wuser[i] ; 
 assign int_wire_desc_n_wuser_4_wuser[i] = int_reg_desc_n_wuser_4_wuser[i] ; 
 assign int_wire_desc_n_wuser_5_wuser[i] = int_reg_desc_n_wuser_5_wuser[i] ; 
 assign int_wire_desc_n_wuser_6_wuser[i] = int_reg_desc_n_wuser_6_wuser[i] ; 
 assign int_wire_desc_n_wuser_7_wuser[i] = int_reg_desc_n_wuser_7_wuser[i] ; 
 assign int_wire_desc_n_wuser_8_wuser[i] = int_reg_desc_n_wuser_8_wuser[i] ; 
 assign int_wire_desc_n_wuser_9_wuser[i] = int_reg_desc_n_wuser_9_wuser[i] ; 
 assign int_wire_desc_n_wuser_10_wuser[i] = int_reg_desc_n_wuser_10_wuser[i] ; 
 assign int_wire_desc_n_wuser_11_wuser[i] = int_reg_desc_n_wuser_11_wuser[i] ; 
 assign int_wire_desc_n_wuser_12_wuser[i] = int_reg_desc_n_wuser_12_wuser[i] ; 
 assign int_wire_desc_n_wuser_13_wuser[i] = int_reg_desc_n_wuser_13_wuser[i] ; 
 assign int_wire_desc_n_wuser_14_wuser[i] = int_reg_desc_n_wuser_14_wuser[i] ; 
 assign int_wire_desc_n_wuser_15_wuser[i] = int_reg_desc_n_wuser_15_wuser[i] ; 
 end //for

endgenerate

