/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */

,input [13:0] int_rd_resp_desc_0_data_offset_addr
 ,input [31:0] int_rd_resp_desc_0_data_size_size
 ,input [31:0] int_rd_resp_desc_0_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_0_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_0_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_0_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_0_resp_resp
 ,input [31:0] int_rd_resp_desc_0_xid_0_xid
 ,input [31:0] int_rd_resp_desc_0_xid_1_xid
 ,input [31:0] int_rd_resp_desc_0_xid_2_xid
 ,input [31:0] int_rd_resp_desc_0_xid_3_xid
 ,input [31:0] int_rd_resp_desc_0_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_0_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_0_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_0_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_0_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_0_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_0_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_0_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_0_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_0_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_0_resp_resp
 ,input [31:0] int_wr_resp_desc_0_xid_0_xid
 ,input [31:0] int_wr_resp_desc_0_xid_1_xid
 ,input [31:0] int_wr_resp_desc_0_xid_2_xid
 ,input [31:0] int_wr_resp_desc_0_xid_3_xid
 ,input [31:0] int_wr_resp_desc_0_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_0_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_0_attr_acsnoop
 ,input [2:0] int_sn_req_desc_0_attr_acprot
 ,input [31:0] int_sn_req_desc_0_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_0_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_0_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_0_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_1_data_offset_addr
 ,input [31:0] int_rd_resp_desc_1_data_size_size
 ,input [31:0] int_rd_resp_desc_1_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_1_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_1_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_1_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_1_resp_resp
 ,input [31:0] int_rd_resp_desc_1_xid_0_xid
 ,input [31:0] int_rd_resp_desc_1_xid_1_xid
 ,input [31:0] int_rd_resp_desc_1_xid_2_xid
 ,input [31:0] int_rd_resp_desc_1_xid_3_xid
 ,input [31:0] int_rd_resp_desc_1_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_1_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_1_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_1_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_1_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_1_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_1_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_1_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_1_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_1_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_1_resp_resp
 ,input [31:0] int_wr_resp_desc_1_xid_0_xid
 ,input [31:0] int_wr_resp_desc_1_xid_1_xid
 ,input [31:0] int_wr_resp_desc_1_xid_2_xid
 ,input [31:0] int_wr_resp_desc_1_xid_3_xid
 ,input [31:0] int_wr_resp_desc_1_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_1_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_1_attr_acsnoop
 ,input [2:0] int_sn_req_desc_1_attr_acprot
 ,input [31:0] int_sn_req_desc_1_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_1_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_1_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_1_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_2_data_offset_addr
 ,input [31:0] int_rd_resp_desc_2_data_size_size
 ,input [31:0] int_rd_resp_desc_2_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_2_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_2_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_2_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_2_resp_resp
 ,input [31:0] int_rd_resp_desc_2_xid_0_xid
 ,input [31:0] int_rd_resp_desc_2_xid_1_xid
 ,input [31:0] int_rd_resp_desc_2_xid_2_xid
 ,input [31:0] int_rd_resp_desc_2_xid_3_xid
 ,input [31:0] int_rd_resp_desc_2_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_2_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_2_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_2_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_2_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_2_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_2_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_2_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_2_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_2_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_2_resp_resp
 ,input [31:0] int_wr_resp_desc_2_xid_0_xid
 ,input [31:0] int_wr_resp_desc_2_xid_1_xid
 ,input [31:0] int_wr_resp_desc_2_xid_2_xid
 ,input [31:0] int_wr_resp_desc_2_xid_3_xid
 ,input [31:0] int_wr_resp_desc_2_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_2_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_2_attr_acsnoop
 ,input [2:0] int_sn_req_desc_2_attr_acprot
 ,input [31:0] int_sn_req_desc_2_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_2_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_2_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_2_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_3_data_offset_addr
 ,input [31:0] int_rd_resp_desc_3_data_size_size
 ,input [31:0] int_rd_resp_desc_3_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_3_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_3_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_3_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_3_resp_resp
 ,input [31:0] int_rd_resp_desc_3_xid_0_xid
 ,input [31:0] int_rd_resp_desc_3_xid_1_xid
 ,input [31:0] int_rd_resp_desc_3_xid_2_xid
 ,input [31:0] int_rd_resp_desc_3_xid_3_xid
 ,input [31:0] int_rd_resp_desc_3_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_3_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_3_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_3_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_3_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_3_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_3_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_3_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_3_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_3_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_3_resp_resp
 ,input [31:0] int_wr_resp_desc_3_xid_0_xid
 ,input [31:0] int_wr_resp_desc_3_xid_1_xid
 ,input [31:0] int_wr_resp_desc_3_xid_2_xid
 ,input [31:0] int_wr_resp_desc_3_xid_3_xid
 ,input [31:0] int_wr_resp_desc_3_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_3_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_3_attr_acsnoop
 ,input [2:0] int_sn_req_desc_3_attr_acprot
 ,input [31:0] int_sn_req_desc_3_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_3_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_3_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_3_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_4_data_offset_addr
 ,input [31:0] int_rd_resp_desc_4_data_size_size
 ,input [31:0] int_rd_resp_desc_4_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_4_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_4_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_4_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_4_resp_resp
 ,input [31:0] int_rd_resp_desc_4_xid_0_xid
 ,input [31:0] int_rd_resp_desc_4_xid_1_xid
 ,input [31:0] int_rd_resp_desc_4_xid_2_xid
 ,input [31:0] int_rd_resp_desc_4_xid_3_xid
 ,input [31:0] int_rd_resp_desc_4_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_4_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_4_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_4_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_4_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_4_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_4_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_4_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_4_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_4_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_4_resp_resp
 ,input [31:0] int_wr_resp_desc_4_xid_0_xid
 ,input [31:0] int_wr_resp_desc_4_xid_1_xid
 ,input [31:0] int_wr_resp_desc_4_xid_2_xid
 ,input [31:0] int_wr_resp_desc_4_xid_3_xid
 ,input [31:0] int_wr_resp_desc_4_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_4_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_4_attr_acsnoop
 ,input [2:0] int_sn_req_desc_4_attr_acprot
 ,input [31:0] int_sn_req_desc_4_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_4_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_4_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_4_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_5_data_offset_addr
 ,input [31:0] int_rd_resp_desc_5_data_size_size
 ,input [31:0] int_rd_resp_desc_5_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_5_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_5_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_5_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_5_resp_resp
 ,input [31:0] int_rd_resp_desc_5_xid_0_xid
 ,input [31:0] int_rd_resp_desc_5_xid_1_xid
 ,input [31:0] int_rd_resp_desc_5_xid_2_xid
 ,input [31:0] int_rd_resp_desc_5_xid_3_xid
 ,input [31:0] int_rd_resp_desc_5_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_5_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_5_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_5_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_5_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_5_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_5_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_5_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_5_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_5_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_5_resp_resp
 ,input [31:0] int_wr_resp_desc_5_xid_0_xid
 ,input [31:0] int_wr_resp_desc_5_xid_1_xid
 ,input [31:0] int_wr_resp_desc_5_xid_2_xid
 ,input [31:0] int_wr_resp_desc_5_xid_3_xid
 ,input [31:0] int_wr_resp_desc_5_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_5_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_5_attr_acsnoop
 ,input [2:0] int_sn_req_desc_5_attr_acprot
 ,input [31:0] int_sn_req_desc_5_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_5_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_5_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_5_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_6_data_offset_addr
 ,input [31:0] int_rd_resp_desc_6_data_size_size
 ,input [31:0] int_rd_resp_desc_6_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_6_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_6_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_6_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_6_resp_resp
 ,input [31:0] int_rd_resp_desc_6_xid_0_xid
 ,input [31:0] int_rd_resp_desc_6_xid_1_xid
 ,input [31:0] int_rd_resp_desc_6_xid_2_xid
 ,input [31:0] int_rd_resp_desc_6_xid_3_xid
 ,input [31:0] int_rd_resp_desc_6_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_6_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_6_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_6_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_6_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_6_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_6_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_6_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_6_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_6_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_6_resp_resp
 ,input [31:0] int_wr_resp_desc_6_xid_0_xid
 ,input [31:0] int_wr_resp_desc_6_xid_1_xid
 ,input [31:0] int_wr_resp_desc_6_xid_2_xid
 ,input [31:0] int_wr_resp_desc_6_xid_3_xid
 ,input [31:0] int_wr_resp_desc_6_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_6_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_6_attr_acsnoop
 ,input [2:0] int_sn_req_desc_6_attr_acprot
 ,input [31:0] int_sn_req_desc_6_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_6_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_6_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_6_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_7_data_offset_addr
 ,input [31:0] int_rd_resp_desc_7_data_size_size
 ,input [31:0] int_rd_resp_desc_7_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_7_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_7_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_7_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_7_resp_resp
 ,input [31:0] int_rd_resp_desc_7_xid_0_xid
 ,input [31:0] int_rd_resp_desc_7_xid_1_xid
 ,input [31:0] int_rd_resp_desc_7_xid_2_xid
 ,input [31:0] int_rd_resp_desc_7_xid_3_xid
 ,input [31:0] int_rd_resp_desc_7_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_7_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_7_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_7_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_7_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_7_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_7_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_7_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_7_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_7_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_7_resp_resp
 ,input [31:0] int_wr_resp_desc_7_xid_0_xid
 ,input [31:0] int_wr_resp_desc_7_xid_1_xid
 ,input [31:0] int_wr_resp_desc_7_xid_2_xid
 ,input [31:0] int_wr_resp_desc_7_xid_3_xid
 ,input [31:0] int_wr_resp_desc_7_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_7_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_7_attr_acsnoop
 ,input [2:0] int_sn_req_desc_7_attr_acprot
 ,input [31:0] int_sn_req_desc_7_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_7_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_7_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_7_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_8_data_offset_addr
 ,input [31:0] int_rd_resp_desc_8_data_size_size
 ,input [31:0] int_rd_resp_desc_8_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_8_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_8_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_8_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_8_resp_resp
 ,input [31:0] int_rd_resp_desc_8_xid_0_xid
 ,input [31:0] int_rd_resp_desc_8_xid_1_xid
 ,input [31:0] int_rd_resp_desc_8_xid_2_xid
 ,input [31:0] int_rd_resp_desc_8_xid_3_xid
 ,input [31:0] int_rd_resp_desc_8_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_8_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_8_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_8_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_8_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_8_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_8_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_8_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_8_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_8_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_8_resp_resp
 ,input [31:0] int_wr_resp_desc_8_xid_0_xid
 ,input [31:0] int_wr_resp_desc_8_xid_1_xid
 ,input [31:0] int_wr_resp_desc_8_xid_2_xid
 ,input [31:0] int_wr_resp_desc_8_xid_3_xid
 ,input [31:0] int_wr_resp_desc_8_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_8_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_8_attr_acsnoop
 ,input [2:0] int_sn_req_desc_8_attr_acprot
 ,input [31:0] int_sn_req_desc_8_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_8_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_8_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_8_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_9_data_offset_addr
 ,input [31:0] int_rd_resp_desc_9_data_size_size
 ,input [31:0] int_rd_resp_desc_9_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_9_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_9_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_9_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_9_resp_resp
 ,input [31:0] int_rd_resp_desc_9_xid_0_xid
 ,input [31:0] int_rd_resp_desc_9_xid_1_xid
 ,input [31:0] int_rd_resp_desc_9_xid_2_xid
 ,input [31:0] int_rd_resp_desc_9_xid_3_xid
 ,input [31:0] int_rd_resp_desc_9_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_9_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_9_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_9_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_9_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_9_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_9_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_9_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_9_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_9_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_9_resp_resp
 ,input [31:0] int_wr_resp_desc_9_xid_0_xid
 ,input [31:0] int_wr_resp_desc_9_xid_1_xid
 ,input [31:0] int_wr_resp_desc_9_xid_2_xid
 ,input [31:0] int_wr_resp_desc_9_xid_3_xid
 ,input [31:0] int_wr_resp_desc_9_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_9_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_9_attr_acsnoop
 ,input [2:0] int_sn_req_desc_9_attr_acprot
 ,input [31:0] int_sn_req_desc_9_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_9_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_9_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_9_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_a_data_offset_addr
 ,input [31:0] int_rd_resp_desc_a_data_size_size
 ,input [31:0] int_rd_resp_desc_a_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_a_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_a_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_a_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_a_resp_resp
 ,input [31:0] int_rd_resp_desc_a_xid_0_xid
 ,input [31:0] int_rd_resp_desc_a_xid_1_xid
 ,input [31:0] int_rd_resp_desc_a_xid_2_xid
 ,input [31:0] int_rd_resp_desc_a_xid_3_xid
 ,input [31:0] int_rd_resp_desc_a_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_a_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_a_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_a_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_a_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_a_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_a_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_a_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_a_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_a_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_a_resp_resp
 ,input [31:0] int_wr_resp_desc_a_xid_0_xid
 ,input [31:0] int_wr_resp_desc_a_xid_1_xid
 ,input [31:0] int_wr_resp_desc_a_xid_2_xid
 ,input [31:0] int_wr_resp_desc_a_xid_3_xid
 ,input [31:0] int_wr_resp_desc_a_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_a_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_a_attr_acsnoop
 ,input [2:0] int_sn_req_desc_a_attr_acprot
 ,input [31:0] int_sn_req_desc_a_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_a_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_a_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_a_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_b_data_offset_addr
 ,input [31:0] int_rd_resp_desc_b_data_size_size
 ,input [31:0] int_rd_resp_desc_b_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_b_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_b_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_b_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_b_resp_resp
 ,input [31:0] int_rd_resp_desc_b_xid_0_xid
 ,input [31:0] int_rd_resp_desc_b_xid_1_xid
 ,input [31:0] int_rd_resp_desc_b_xid_2_xid
 ,input [31:0] int_rd_resp_desc_b_xid_3_xid
 ,input [31:0] int_rd_resp_desc_b_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_b_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_b_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_b_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_b_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_b_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_b_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_b_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_b_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_b_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_b_resp_resp
 ,input [31:0] int_wr_resp_desc_b_xid_0_xid
 ,input [31:0] int_wr_resp_desc_b_xid_1_xid
 ,input [31:0] int_wr_resp_desc_b_xid_2_xid
 ,input [31:0] int_wr_resp_desc_b_xid_3_xid
 ,input [31:0] int_wr_resp_desc_b_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_b_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_b_attr_acsnoop
 ,input [2:0] int_sn_req_desc_b_attr_acprot
 ,input [31:0] int_sn_req_desc_b_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_b_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_b_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_b_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_c_data_offset_addr
 ,input [31:0] int_rd_resp_desc_c_data_size_size
 ,input [31:0] int_rd_resp_desc_c_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_c_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_c_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_c_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_c_resp_resp
 ,input [31:0] int_rd_resp_desc_c_xid_0_xid
 ,input [31:0] int_rd_resp_desc_c_xid_1_xid
 ,input [31:0] int_rd_resp_desc_c_xid_2_xid
 ,input [31:0] int_rd_resp_desc_c_xid_3_xid
 ,input [31:0] int_rd_resp_desc_c_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_c_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_c_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_c_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_c_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_c_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_c_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_c_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_c_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_c_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_c_resp_resp
 ,input [31:0] int_wr_resp_desc_c_xid_0_xid
 ,input [31:0] int_wr_resp_desc_c_xid_1_xid
 ,input [31:0] int_wr_resp_desc_c_xid_2_xid
 ,input [31:0] int_wr_resp_desc_c_xid_3_xid
 ,input [31:0] int_wr_resp_desc_c_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_c_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_c_attr_acsnoop
 ,input [2:0] int_sn_req_desc_c_attr_acprot
 ,input [31:0] int_sn_req_desc_c_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_c_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_c_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_c_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_d_data_offset_addr
 ,input [31:0] int_rd_resp_desc_d_data_size_size
 ,input [31:0] int_rd_resp_desc_d_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_d_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_d_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_d_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_d_resp_resp
 ,input [31:0] int_rd_resp_desc_d_xid_0_xid
 ,input [31:0] int_rd_resp_desc_d_xid_1_xid
 ,input [31:0] int_rd_resp_desc_d_xid_2_xid
 ,input [31:0] int_rd_resp_desc_d_xid_3_xid
 ,input [31:0] int_rd_resp_desc_d_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_d_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_d_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_d_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_d_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_d_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_d_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_d_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_d_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_d_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_d_resp_resp
 ,input [31:0] int_wr_resp_desc_d_xid_0_xid
 ,input [31:0] int_wr_resp_desc_d_xid_1_xid
 ,input [31:0] int_wr_resp_desc_d_xid_2_xid
 ,input [31:0] int_wr_resp_desc_d_xid_3_xid
 ,input [31:0] int_wr_resp_desc_d_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_d_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_d_attr_acsnoop
 ,input [2:0] int_sn_req_desc_d_attr_acprot
 ,input [31:0] int_sn_req_desc_d_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_d_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_d_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_d_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_e_data_offset_addr
 ,input [31:0] int_rd_resp_desc_e_data_size_size
 ,input [31:0] int_rd_resp_desc_e_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_e_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_e_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_e_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_e_resp_resp
 ,input [31:0] int_rd_resp_desc_e_xid_0_xid
 ,input [31:0] int_rd_resp_desc_e_xid_1_xid
 ,input [31:0] int_rd_resp_desc_e_xid_2_xid
 ,input [31:0] int_rd_resp_desc_e_xid_3_xid
 ,input [31:0] int_rd_resp_desc_e_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_e_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_e_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_e_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_e_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_e_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_e_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_e_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_e_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_e_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_e_resp_resp
 ,input [31:0] int_wr_resp_desc_e_xid_0_xid
 ,input [31:0] int_wr_resp_desc_e_xid_1_xid
 ,input [31:0] int_wr_resp_desc_e_xid_2_xid
 ,input [31:0] int_wr_resp_desc_e_xid_3_xid
 ,input [31:0] int_wr_resp_desc_e_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_e_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_e_attr_acsnoop
 ,input [2:0] int_sn_req_desc_e_attr_acprot
 ,input [31:0] int_sn_req_desc_e_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_e_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_e_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_e_acaddr_3_addr
 ,input [13:0] int_rd_resp_desc_f_data_offset_addr
 ,input [31:0] int_rd_resp_desc_f_data_size_size
 ,input [31:0] int_rd_resp_desc_f_data_host_addr_0_addr
 ,input [31:0] int_rd_resp_desc_f_data_host_addr_1_addr
 ,input [31:0] int_rd_resp_desc_f_data_host_addr_2_addr
 ,input [31:0] int_rd_resp_desc_f_data_host_addr_3_addr
 ,input [4:0] int_rd_resp_desc_f_resp_resp
 ,input [31:0] int_rd_resp_desc_f_xid_0_xid
 ,input [31:0] int_rd_resp_desc_f_xid_1_xid
 ,input [31:0] int_rd_resp_desc_f_xid_2_xid
 ,input [31:0] int_rd_resp_desc_f_xid_3_xid
 ,input [31:0] int_rd_resp_desc_f_xuser_0_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_1_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_2_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_3_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_4_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_5_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_6_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_7_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_8_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_9_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_10_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_11_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_12_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_13_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_14_xuser
 ,input [31:0] int_rd_resp_desc_f_xuser_15_xuser
 ,input [31:0] int_wr_req_desc_f_data_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_f_data_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_f_data_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_f_data_host_addr_3_addr
 ,input [31:0] int_wr_req_desc_f_wstrb_host_addr_0_addr
 ,input [31:0] int_wr_req_desc_f_wstrb_host_addr_1_addr
 ,input [31:0] int_wr_req_desc_f_wstrb_host_addr_2_addr
 ,input [31:0] int_wr_req_desc_f_wstrb_host_addr_3_addr
 ,input [4:0] int_wr_resp_desc_f_resp_resp
 ,input [31:0] int_wr_resp_desc_f_xid_0_xid
 ,input [31:0] int_wr_resp_desc_f_xid_1_xid
 ,input [31:0] int_wr_resp_desc_f_xid_2_xid
 ,input [31:0] int_wr_resp_desc_f_xid_3_xid
 ,input [31:0] int_wr_resp_desc_f_xuser_0_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_1_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_2_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_3_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_4_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_5_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_6_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_7_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_8_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_9_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_10_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_11_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_12_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_13_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_14_xuser
 ,input [31:0] int_wr_resp_desc_f_xuser_15_xuser
 ,input [3:0] int_sn_req_desc_f_attr_acsnoop
 ,input [2:0] int_sn_req_desc_f_attr_acprot
 ,input [31:0] int_sn_req_desc_f_acaddr_0_addr
 ,input [31:0] int_sn_req_desc_f_acaddr_1_addr
 ,input [31:0] int_sn_req_desc_f_acaddr_2_addr
 ,input [31:0] int_sn_req_desc_f_acaddr_3_addr
 ,output [31:0] int_rd_req_desc_0_size_txn_size
 ,output [2:0] int_rd_req_desc_0_axsize_axsize
 ,output [3:0] int_rd_req_desc_0_attr_axsnoop
 ,output [1:0] int_rd_req_desc_0_attr_axdomain
 ,output [1:0] int_rd_req_desc_0_attr_axbar
 ,output [3:0] int_rd_req_desc_0_attr_axregion
 ,output [3:0] int_rd_req_desc_0_attr_axqos
 ,output [2:0] int_rd_req_desc_0_attr_axprot
 ,output [3:0] int_rd_req_desc_0_attr_axcache
 ,output [0:0] int_rd_req_desc_0_attr_axlock
 ,output [1:0] int_rd_req_desc_0_attr_axburst
 ,output [31:0] int_rd_req_desc_0_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_0_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_0_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_0_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_0_axid_0_axid
 ,output [31:0] int_rd_req_desc_0_axid_1_axid
 ,output [31:0] int_rd_req_desc_0_axid_2_axid
 ,output [31:0] int_rd_req_desc_0_axid_3_axid
 ,output [31:0] int_rd_req_desc_0_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_0_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_0_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_0_size_txn_size
 ,output [13:0] int_wr_req_desc_0_data_offset_addr
 ,output [2:0] int_wr_req_desc_0_axsize_axsize
 ,output [3:0] int_wr_req_desc_0_attr_axsnoop
 ,output [1:0] int_wr_req_desc_0_attr_axdomain
 ,output [1:0] int_wr_req_desc_0_attr_axbar
 ,output [0:0] int_wr_req_desc_0_attr_awunique
 ,output [3:0] int_wr_req_desc_0_attr_axregion
 ,output [3:0] int_wr_req_desc_0_attr_axqos
 ,output [2:0] int_wr_req_desc_0_attr_axprot
 ,output [3:0] int_wr_req_desc_0_attr_axcache
 ,output [0:0] int_wr_req_desc_0_attr_axlock
 ,output [1:0] int_wr_req_desc_0_attr_axburst
 ,output [31:0] int_wr_req_desc_0_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_0_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_0_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_0_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_0_axid_0_axid
 ,output [31:0] int_wr_req_desc_0_axid_1_axid
 ,output [31:0] int_wr_req_desc_0_axid_2_axid
 ,output [31:0] int_wr_req_desc_0_axid_3_axid
 ,output [31:0] int_wr_req_desc_0_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_0_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_0_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_0_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_0_resp_resp
 ,output [31:0] int_rd_req_desc_1_size_txn_size
 ,output [2:0] int_rd_req_desc_1_axsize_axsize
 ,output [3:0] int_rd_req_desc_1_attr_axsnoop
 ,output [1:0] int_rd_req_desc_1_attr_axdomain
 ,output [1:0] int_rd_req_desc_1_attr_axbar
 ,output [3:0] int_rd_req_desc_1_attr_axregion
 ,output [3:0] int_rd_req_desc_1_attr_axqos
 ,output [2:0] int_rd_req_desc_1_attr_axprot
 ,output [3:0] int_rd_req_desc_1_attr_axcache
 ,output [0:0] int_rd_req_desc_1_attr_axlock
 ,output [1:0] int_rd_req_desc_1_attr_axburst
 ,output [31:0] int_rd_req_desc_1_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_1_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_1_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_1_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_1_axid_0_axid
 ,output [31:0] int_rd_req_desc_1_axid_1_axid
 ,output [31:0] int_rd_req_desc_1_axid_2_axid
 ,output [31:0] int_rd_req_desc_1_axid_3_axid
 ,output [31:0] int_rd_req_desc_1_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_1_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_1_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_1_size_txn_size
 ,output [13:0] int_wr_req_desc_1_data_offset_addr
 ,output [2:0] int_wr_req_desc_1_axsize_axsize
 ,output [3:0] int_wr_req_desc_1_attr_axsnoop
 ,output [1:0] int_wr_req_desc_1_attr_axdomain
 ,output [1:0] int_wr_req_desc_1_attr_axbar
 ,output [0:0] int_wr_req_desc_1_attr_awunique
 ,output [3:0] int_wr_req_desc_1_attr_axregion
 ,output [3:0] int_wr_req_desc_1_attr_axqos
 ,output [2:0] int_wr_req_desc_1_attr_axprot
 ,output [3:0] int_wr_req_desc_1_attr_axcache
 ,output [0:0] int_wr_req_desc_1_attr_axlock
 ,output [1:0] int_wr_req_desc_1_attr_axburst
 ,output [31:0] int_wr_req_desc_1_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_1_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_1_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_1_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_1_axid_0_axid
 ,output [31:0] int_wr_req_desc_1_axid_1_axid
 ,output [31:0] int_wr_req_desc_1_axid_2_axid
 ,output [31:0] int_wr_req_desc_1_axid_3_axid
 ,output [31:0] int_wr_req_desc_1_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_1_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_1_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_1_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_1_resp_resp
 ,output [31:0] int_rd_req_desc_2_size_txn_size
 ,output [2:0] int_rd_req_desc_2_axsize_axsize
 ,output [3:0] int_rd_req_desc_2_attr_axsnoop
 ,output [1:0] int_rd_req_desc_2_attr_axdomain
 ,output [1:0] int_rd_req_desc_2_attr_axbar
 ,output [3:0] int_rd_req_desc_2_attr_axregion
 ,output [3:0] int_rd_req_desc_2_attr_axqos
 ,output [2:0] int_rd_req_desc_2_attr_axprot
 ,output [3:0] int_rd_req_desc_2_attr_axcache
 ,output [0:0] int_rd_req_desc_2_attr_axlock
 ,output [1:0] int_rd_req_desc_2_attr_axburst
 ,output [31:0] int_rd_req_desc_2_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_2_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_2_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_2_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_2_axid_0_axid
 ,output [31:0] int_rd_req_desc_2_axid_1_axid
 ,output [31:0] int_rd_req_desc_2_axid_2_axid
 ,output [31:0] int_rd_req_desc_2_axid_3_axid
 ,output [31:0] int_rd_req_desc_2_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_2_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_2_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_2_size_txn_size
 ,output [13:0] int_wr_req_desc_2_data_offset_addr
 ,output [2:0] int_wr_req_desc_2_axsize_axsize
 ,output [3:0] int_wr_req_desc_2_attr_axsnoop
 ,output [1:0] int_wr_req_desc_2_attr_axdomain
 ,output [1:0] int_wr_req_desc_2_attr_axbar
 ,output [0:0] int_wr_req_desc_2_attr_awunique
 ,output [3:0] int_wr_req_desc_2_attr_axregion
 ,output [3:0] int_wr_req_desc_2_attr_axqos
 ,output [2:0] int_wr_req_desc_2_attr_axprot
 ,output [3:0] int_wr_req_desc_2_attr_axcache
 ,output [0:0] int_wr_req_desc_2_attr_axlock
 ,output [1:0] int_wr_req_desc_2_attr_axburst
 ,output [31:0] int_wr_req_desc_2_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_2_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_2_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_2_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_2_axid_0_axid
 ,output [31:0] int_wr_req_desc_2_axid_1_axid
 ,output [31:0] int_wr_req_desc_2_axid_2_axid
 ,output [31:0] int_wr_req_desc_2_axid_3_axid
 ,output [31:0] int_wr_req_desc_2_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_2_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_2_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_2_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_2_resp_resp
 ,output [31:0] int_rd_req_desc_3_size_txn_size
 ,output [2:0] int_rd_req_desc_3_axsize_axsize
 ,output [3:0] int_rd_req_desc_3_attr_axsnoop
 ,output [1:0] int_rd_req_desc_3_attr_axdomain
 ,output [1:0] int_rd_req_desc_3_attr_axbar
 ,output [3:0] int_rd_req_desc_3_attr_axregion
 ,output [3:0] int_rd_req_desc_3_attr_axqos
 ,output [2:0] int_rd_req_desc_3_attr_axprot
 ,output [3:0] int_rd_req_desc_3_attr_axcache
 ,output [0:0] int_rd_req_desc_3_attr_axlock
 ,output [1:0] int_rd_req_desc_3_attr_axburst
 ,output [31:0] int_rd_req_desc_3_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_3_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_3_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_3_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_3_axid_0_axid
 ,output [31:0] int_rd_req_desc_3_axid_1_axid
 ,output [31:0] int_rd_req_desc_3_axid_2_axid
 ,output [31:0] int_rd_req_desc_3_axid_3_axid
 ,output [31:0] int_rd_req_desc_3_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_3_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_3_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_3_size_txn_size
 ,output [13:0] int_wr_req_desc_3_data_offset_addr
 ,output [2:0] int_wr_req_desc_3_axsize_axsize
 ,output [3:0] int_wr_req_desc_3_attr_axsnoop
 ,output [1:0] int_wr_req_desc_3_attr_axdomain
 ,output [1:0] int_wr_req_desc_3_attr_axbar
 ,output [0:0] int_wr_req_desc_3_attr_awunique
 ,output [3:0] int_wr_req_desc_3_attr_axregion
 ,output [3:0] int_wr_req_desc_3_attr_axqos
 ,output [2:0] int_wr_req_desc_3_attr_axprot
 ,output [3:0] int_wr_req_desc_3_attr_axcache
 ,output [0:0] int_wr_req_desc_3_attr_axlock
 ,output [1:0] int_wr_req_desc_3_attr_axburst
 ,output [31:0] int_wr_req_desc_3_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_3_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_3_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_3_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_3_axid_0_axid
 ,output [31:0] int_wr_req_desc_3_axid_1_axid
 ,output [31:0] int_wr_req_desc_3_axid_2_axid
 ,output [31:0] int_wr_req_desc_3_axid_3_axid
 ,output [31:0] int_wr_req_desc_3_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_3_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_3_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_3_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_3_resp_resp
 ,output [31:0] int_rd_req_desc_4_size_txn_size
 ,output [2:0] int_rd_req_desc_4_axsize_axsize
 ,output [3:0] int_rd_req_desc_4_attr_axsnoop
 ,output [1:0] int_rd_req_desc_4_attr_axdomain
 ,output [1:0] int_rd_req_desc_4_attr_axbar
 ,output [3:0] int_rd_req_desc_4_attr_axregion
 ,output [3:0] int_rd_req_desc_4_attr_axqos
 ,output [2:0] int_rd_req_desc_4_attr_axprot
 ,output [3:0] int_rd_req_desc_4_attr_axcache
 ,output [0:0] int_rd_req_desc_4_attr_axlock
 ,output [1:0] int_rd_req_desc_4_attr_axburst
 ,output [31:0] int_rd_req_desc_4_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_4_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_4_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_4_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_4_axid_0_axid
 ,output [31:0] int_rd_req_desc_4_axid_1_axid
 ,output [31:0] int_rd_req_desc_4_axid_2_axid
 ,output [31:0] int_rd_req_desc_4_axid_3_axid
 ,output [31:0] int_rd_req_desc_4_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_4_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_4_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_4_size_txn_size
 ,output [13:0] int_wr_req_desc_4_data_offset_addr
 ,output [2:0] int_wr_req_desc_4_axsize_axsize
 ,output [3:0] int_wr_req_desc_4_attr_axsnoop
 ,output [1:0] int_wr_req_desc_4_attr_axdomain
 ,output [1:0] int_wr_req_desc_4_attr_axbar
 ,output [0:0] int_wr_req_desc_4_attr_awunique
 ,output [3:0] int_wr_req_desc_4_attr_axregion
 ,output [3:0] int_wr_req_desc_4_attr_axqos
 ,output [2:0] int_wr_req_desc_4_attr_axprot
 ,output [3:0] int_wr_req_desc_4_attr_axcache
 ,output [0:0] int_wr_req_desc_4_attr_axlock
 ,output [1:0] int_wr_req_desc_4_attr_axburst
 ,output [31:0] int_wr_req_desc_4_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_4_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_4_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_4_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_4_axid_0_axid
 ,output [31:0] int_wr_req_desc_4_axid_1_axid
 ,output [31:0] int_wr_req_desc_4_axid_2_axid
 ,output [31:0] int_wr_req_desc_4_axid_3_axid
 ,output [31:0] int_wr_req_desc_4_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_4_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_4_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_4_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_4_resp_resp
 ,output [31:0] int_rd_req_desc_5_size_txn_size
 ,output [2:0] int_rd_req_desc_5_axsize_axsize
 ,output [3:0] int_rd_req_desc_5_attr_axsnoop
 ,output [1:0] int_rd_req_desc_5_attr_axdomain
 ,output [1:0] int_rd_req_desc_5_attr_axbar
 ,output [3:0] int_rd_req_desc_5_attr_axregion
 ,output [3:0] int_rd_req_desc_5_attr_axqos
 ,output [2:0] int_rd_req_desc_5_attr_axprot
 ,output [3:0] int_rd_req_desc_5_attr_axcache
 ,output [0:0] int_rd_req_desc_5_attr_axlock
 ,output [1:0] int_rd_req_desc_5_attr_axburst
 ,output [31:0] int_rd_req_desc_5_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_5_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_5_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_5_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_5_axid_0_axid
 ,output [31:0] int_rd_req_desc_5_axid_1_axid
 ,output [31:0] int_rd_req_desc_5_axid_2_axid
 ,output [31:0] int_rd_req_desc_5_axid_3_axid
 ,output [31:0] int_rd_req_desc_5_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_5_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_5_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_5_size_txn_size
 ,output [13:0] int_wr_req_desc_5_data_offset_addr
 ,output [2:0] int_wr_req_desc_5_axsize_axsize
 ,output [3:0] int_wr_req_desc_5_attr_axsnoop
 ,output [1:0] int_wr_req_desc_5_attr_axdomain
 ,output [1:0] int_wr_req_desc_5_attr_axbar
 ,output [0:0] int_wr_req_desc_5_attr_awunique
 ,output [3:0] int_wr_req_desc_5_attr_axregion
 ,output [3:0] int_wr_req_desc_5_attr_axqos
 ,output [2:0] int_wr_req_desc_5_attr_axprot
 ,output [3:0] int_wr_req_desc_5_attr_axcache
 ,output [0:0] int_wr_req_desc_5_attr_axlock
 ,output [1:0] int_wr_req_desc_5_attr_axburst
 ,output [31:0] int_wr_req_desc_5_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_5_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_5_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_5_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_5_axid_0_axid
 ,output [31:0] int_wr_req_desc_5_axid_1_axid
 ,output [31:0] int_wr_req_desc_5_axid_2_axid
 ,output [31:0] int_wr_req_desc_5_axid_3_axid
 ,output [31:0] int_wr_req_desc_5_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_5_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_5_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_5_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_5_resp_resp
 ,output [31:0] int_rd_req_desc_6_size_txn_size
 ,output [2:0] int_rd_req_desc_6_axsize_axsize
 ,output [3:0] int_rd_req_desc_6_attr_axsnoop
 ,output [1:0] int_rd_req_desc_6_attr_axdomain
 ,output [1:0] int_rd_req_desc_6_attr_axbar
 ,output [3:0] int_rd_req_desc_6_attr_axregion
 ,output [3:0] int_rd_req_desc_6_attr_axqos
 ,output [2:0] int_rd_req_desc_6_attr_axprot
 ,output [3:0] int_rd_req_desc_6_attr_axcache
 ,output [0:0] int_rd_req_desc_6_attr_axlock
 ,output [1:0] int_rd_req_desc_6_attr_axburst
 ,output [31:0] int_rd_req_desc_6_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_6_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_6_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_6_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_6_axid_0_axid
 ,output [31:0] int_rd_req_desc_6_axid_1_axid
 ,output [31:0] int_rd_req_desc_6_axid_2_axid
 ,output [31:0] int_rd_req_desc_6_axid_3_axid
 ,output [31:0] int_rd_req_desc_6_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_6_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_6_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_6_size_txn_size
 ,output [13:0] int_wr_req_desc_6_data_offset_addr
 ,output [2:0] int_wr_req_desc_6_axsize_axsize
 ,output [3:0] int_wr_req_desc_6_attr_axsnoop
 ,output [1:0] int_wr_req_desc_6_attr_axdomain
 ,output [1:0] int_wr_req_desc_6_attr_axbar
 ,output [0:0] int_wr_req_desc_6_attr_awunique
 ,output [3:0] int_wr_req_desc_6_attr_axregion
 ,output [3:0] int_wr_req_desc_6_attr_axqos
 ,output [2:0] int_wr_req_desc_6_attr_axprot
 ,output [3:0] int_wr_req_desc_6_attr_axcache
 ,output [0:0] int_wr_req_desc_6_attr_axlock
 ,output [1:0] int_wr_req_desc_6_attr_axburst
 ,output [31:0] int_wr_req_desc_6_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_6_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_6_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_6_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_6_axid_0_axid
 ,output [31:0] int_wr_req_desc_6_axid_1_axid
 ,output [31:0] int_wr_req_desc_6_axid_2_axid
 ,output [31:0] int_wr_req_desc_6_axid_3_axid
 ,output [31:0] int_wr_req_desc_6_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_6_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_6_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_6_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_6_resp_resp
 ,output [31:0] int_rd_req_desc_7_size_txn_size
 ,output [2:0] int_rd_req_desc_7_axsize_axsize
 ,output [3:0] int_rd_req_desc_7_attr_axsnoop
 ,output [1:0] int_rd_req_desc_7_attr_axdomain
 ,output [1:0] int_rd_req_desc_7_attr_axbar
 ,output [3:0] int_rd_req_desc_7_attr_axregion
 ,output [3:0] int_rd_req_desc_7_attr_axqos
 ,output [2:0] int_rd_req_desc_7_attr_axprot
 ,output [3:0] int_rd_req_desc_7_attr_axcache
 ,output [0:0] int_rd_req_desc_7_attr_axlock
 ,output [1:0] int_rd_req_desc_7_attr_axburst
 ,output [31:0] int_rd_req_desc_7_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_7_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_7_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_7_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_7_axid_0_axid
 ,output [31:0] int_rd_req_desc_7_axid_1_axid
 ,output [31:0] int_rd_req_desc_7_axid_2_axid
 ,output [31:0] int_rd_req_desc_7_axid_3_axid
 ,output [31:0] int_rd_req_desc_7_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_7_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_7_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_7_size_txn_size
 ,output [13:0] int_wr_req_desc_7_data_offset_addr
 ,output [2:0] int_wr_req_desc_7_axsize_axsize
 ,output [3:0] int_wr_req_desc_7_attr_axsnoop
 ,output [1:0] int_wr_req_desc_7_attr_axdomain
 ,output [1:0] int_wr_req_desc_7_attr_axbar
 ,output [0:0] int_wr_req_desc_7_attr_awunique
 ,output [3:0] int_wr_req_desc_7_attr_axregion
 ,output [3:0] int_wr_req_desc_7_attr_axqos
 ,output [2:0] int_wr_req_desc_7_attr_axprot
 ,output [3:0] int_wr_req_desc_7_attr_axcache
 ,output [0:0] int_wr_req_desc_7_attr_axlock
 ,output [1:0] int_wr_req_desc_7_attr_axburst
 ,output [31:0] int_wr_req_desc_7_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_7_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_7_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_7_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_7_axid_0_axid
 ,output [31:0] int_wr_req_desc_7_axid_1_axid
 ,output [31:0] int_wr_req_desc_7_axid_2_axid
 ,output [31:0] int_wr_req_desc_7_axid_3_axid
 ,output [31:0] int_wr_req_desc_7_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_7_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_7_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_7_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_7_resp_resp
 ,output [31:0] int_rd_req_desc_8_size_txn_size
 ,output [2:0] int_rd_req_desc_8_axsize_axsize
 ,output [3:0] int_rd_req_desc_8_attr_axsnoop
 ,output [1:0] int_rd_req_desc_8_attr_axdomain
 ,output [1:0] int_rd_req_desc_8_attr_axbar
 ,output [3:0] int_rd_req_desc_8_attr_axregion
 ,output [3:0] int_rd_req_desc_8_attr_axqos
 ,output [2:0] int_rd_req_desc_8_attr_axprot
 ,output [3:0] int_rd_req_desc_8_attr_axcache
 ,output [0:0] int_rd_req_desc_8_attr_axlock
 ,output [1:0] int_rd_req_desc_8_attr_axburst
 ,output [31:0] int_rd_req_desc_8_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_8_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_8_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_8_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_8_axid_0_axid
 ,output [31:0] int_rd_req_desc_8_axid_1_axid
 ,output [31:0] int_rd_req_desc_8_axid_2_axid
 ,output [31:0] int_rd_req_desc_8_axid_3_axid
 ,output [31:0] int_rd_req_desc_8_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_8_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_8_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_8_size_txn_size
 ,output [13:0] int_wr_req_desc_8_data_offset_addr
 ,output [2:0] int_wr_req_desc_8_axsize_axsize
 ,output [3:0] int_wr_req_desc_8_attr_axsnoop
 ,output [1:0] int_wr_req_desc_8_attr_axdomain
 ,output [1:0] int_wr_req_desc_8_attr_axbar
 ,output [0:0] int_wr_req_desc_8_attr_awunique
 ,output [3:0] int_wr_req_desc_8_attr_axregion
 ,output [3:0] int_wr_req_desc_8_attr_axqos
 ,output [2:0] int_wr_req_desc_8_attr_axprot
 ,output [3:0] int_wr_req_desc_8_attr_axcache
 ,output [0:0] int_wr_req_desc_8_attr_axlock
 ,output [1:0] int_wr_req_desc_8_attr_axburst
 ,output [31:0] int_wr_req_desc_8_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_8_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_8_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_8_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_8_axid_0_axid
 ,output [31:0] int_wr_req_desc_8_axid_1_axid
 ,output [31:0] int_wr_req_desc_8_axid_2_axid
 ,output [31:0] int_wr_req_desc_8_axid_3_axid
 ,output [31:0] int_wr_req_desc_8_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_8_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_8_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_8_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_8_resp_resp
 ,output [31:0] int_rd_req_desc_9_size_txn_size
 ,output [2:0] int_rd_req_desc_9_axsize_axsize
 ,output [3:0] int_rd_req_desc_9_attr_axsnoop
 ,output [1:0] int_rd_req_desc_9_attr_axdomain
 ,output [1:0] int_rd_req_desc_9_attr_axbar
 ,output [3:0] int_rd_req_desc_9_attr_axregion
 ,output [3:0] int_rd_req_desc_9_attr_axqos
 ,output [2:0] int_rd_req_desc_9_attr_axprot
 ,output [3:0] int_rd_req_desc_9_attr_axcache
 ,output [0:0] int_rd_req_desc_9_attr_axlock
 ,output [1:0] int_rd_req_desc_9_attr_axburst
 ,output [31:0] int_rd_req_desc_9_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_9_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_9_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_9_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_9_axid_0_axid
 ,output [31:0] int_rd_req_desc_9_axid_1_axid
 ,output [31:0] int_rd_req_desc_9_axid_2_axid
 ,output [31:0] int_rd_req_desc_9_axid_3_axid
 ,output [31:0] int_rd_req_desc_9_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_9_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_9_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_9_size_txn_size
 ,output [13:0] int_wr_req_desc_9_data_offset_addr
 ,output [2:0] int_wr_req_desc_9_axsize_axsize
 ,output [3:0] int_wr_req_desc_9_attr_axsnoop
 ,output [1:0] int_wr_req_desc_9_attr_axdomain
 ,output [1:0] int_wr_req_desc_9_attr_axbar
 ,output [0:0] int_wr_req_desc_9_attr_awunique
 ,output [3:0] int_wr_req_desc_9_attr_axregion
 ,output [3:0] int_wr_req_desc_9_attr_axqos
 ,output [2:0] int_wr_req_desc_9_attr_axprot
 ,output [3:0] int_wr_req_desc_9_attr_axcache
 ,output [0:0] int_wr_req_desc_9_attr_axlock
 ,output [1:0] int_wr_req_desc_9_attr_axburst
 ,output [31:0] int_wr_req_desc_9_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_9_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_9_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_9_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_9_axid_0_axid
 ,output [31:0] int_wr_req_desc_9_axid_1_axid
 ,output [31:0] int_wr_req_desc_9_axid_2_axid
 ,output [31:0] int_wr_req_desc_9_axid_3_axid
 ,output [31:0] int_wr_req_desc_9_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_9_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_9_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_9_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_9_resp_resp
 ,output [31:0] int_rd_req_desc_a_size_txn_size
 ,output [2:0] int_rd_req_desc_a_axsize_axsize
 ,output [3:0] int_rd_req_desc_a_attr_axsnoop
 ,output [1:0] int_rd_req_desc_a_attr_axdomain
 ,output [1:0] int_rd_req_desc_a_attr_axbar
 ,output [3:0] int_rd_req_desc_a_attr_axregion
 ,output [3:0] int_rd_req_desc_a_attr_axqos
 ,output [2:0] int_rd_req_desc_a_attr_axprot
 ,output [3:0] int_rd_req_desc_a_attr_axcache
 ,output [0:0] int_rd_req_desc_a_attr_axlock
 ,output [1:0] int_rd_req_desc_a_attr_axburst
 ,output [31:0] int_rd_req_desc_a_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_a_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_a_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_a_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_a_axid_0_axid
 ,output [31:0] int_rd_req_desc_a_axid_1_axid
 ,output [31:0] int_rd_req_desc_a_axid_2_axid
 ,output [31:0] int_rd_req_desc_a_axid_3_axid
 ,output [31:0] int_rd_req_desc_a_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_a_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_a_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_a_size_txn_size
 ,output [13:0] int_wr_req_desc_a_data_offset_addr
 ,output [2:0] int_wr_req_desc_a_axsize_axsize
 ,output [3:0] int_wr_req_desc_a_attr_axsnoop
 ,output [1:0] int_wr_req_desc_a_attr_axdomain
 ,output [1:0] int_wr_req_desc_a_attr_axbar
 ,output [0:0] int_wr_req_desc_a_attr_awunique
 ,output [3:0] int_wr_req_desc_a_attr_axregion
 ,output [3:0] int_wr_req_desc_a_attr_axqos
 ,output [2:0] int_wr_req_desc_a_attr_axprot
 ,output [3:0] int_wr_req_desc_a_attr_axcache
 ,output [0:0] int_wr_req_desc_a_attr_axlock
 ,output [1:0] int_wr_req_desc_a_attr_axburst
 ,output [31:0] int_wr_req_desc_a_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_a_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_a_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_a_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_a_axid_0_axid
 ,output [31:0] int_wr_req_desc_a_axid_1_axid
 ,output [31:0] int_wr_req_desc_a_axid_2_axid
 ,output [31:0] int_wr_req_desc_a_axid_3_axid
 ,output [31:0] int_wr_req_desc_a_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_a_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_a_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_a_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_a_resp_resp
 ,output [31:0] int_rd_req_desc_b_size_txn_size
 ,output [2:0] int_rd_req_desc_b_axsize_axsize
 ,output [3:0] int_rd_req_desc_b_attr_axsnoop
 ,output [1:0] int_rd_req_desc_b_attr_axdomain
 ,output [1:0] int_rd_req_desc_b_attr_axbar
 ,output [3:0] int_rd_req_desc_b_attr_axregion
 ,output [3:0] int_rd_req_desc_b_attr_axqos
 ,output [2:0] int_rd_req_desc_b_attr_axprot
 ,output [3:0] int_rd_req_desc_b_attr_axcache
 ,output [0:0] int_rd_req_desc_b_attr_axlock
 ,output [1:0] int_rd_req_desc_b_attr_axburst
 ,output [31:0] int_rd_req_desc_b_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_b_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_b_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_b_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_b_axid_0_axid
 ,output [31:0] int_rd_req_desc_b_axid_1_axid
 ,output [31:0] int_rd_req_desc_b_axid_2_axid
 ,output [31:0] int_rd_req_desc_b_axid_3_axid
 ,output [31:0] int_rd_req_desc_b_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_b_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_b_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_b_size_txn_size
 ,output [13:0] int_wr_req_desc_b_data_offset_addr
 ,output [2:0] int_wr_req_desc_b_axsize_axsize
 ,output [3:0] int_wr_req_desc_b_attr_axsnoop
 ,output [1:0] int_wr_req_desc_b_attr_axdomain
 ,output [1:0] int_wr_req_desc_b_attr_axbar
 ,output [0:0] int_wr_req_desc_b_attr_awunique
 ,output [3:0] int_wr_req_desc_b_attr_axregion
 ,output [3:0] int_wr_req_desc_b_attr_axqos
 ,output [2:0] int_wr_req_desc_b_attr_axprot
 ,output [3:0] int_wr_req_desc_b_attr_axcache
 ,output [0:0] int_wr_req_desc_b_attr_axlock
 ,output [1:0] int_wr_req_desc_b_attr_axburst
 ,output [31:0] int_wr_req_desc_b_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_b_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_b_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_b_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_b_axid_0_axid
 ,output [31:0] int_wr_req_desc_b_axid_1_axid
 ,output [31:0] int_wr_req_desc_b_axid_2_axid
 ,output [31:0] int_wr_req_desc_b_axid_3_axid
 ,output [31:0] int_wr_req_desc_b_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_b_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_b_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_b_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_b_resp_resp
 ,output [31:0] int_rd_req_desc_c_size_txn_size
 ,output [2:0] int_rd_req_desc_c_axsize_axsize
 ,output [3:0] int_rd_req_desc_c_attr_axsnoop
 ,output [1:0] int_rd_req_desc_c_attr_axdomain
 ,output [1:0] int_rd_req_desc_c_attr_axbar
 ,output [3:0] int_rd_req_desc_c_attr_axregion
 ,output [3:0] int_rd_req_desc_c_attr_axqos
 ,output [2:0] int_rd_req_desc_c_attr_axprot
 ,output [3:0] int_rd_req_desc_c_attr_axcache
 ,output [0:0] int_rd_req_desc_c_attr_axlock
 ,output [1:0] int_rd_req_desc_c_attr_axburst
 ,output [31:0] int_rd_req_desc_c_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_c_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_c_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_c_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_c_axid_0_axid
 ,output [31:0] int_rd_req_desc_c_axid_1_axid
 ,output [31:0] int_rd_req_desc_c_axid_2_axid
 ,output [31:0] int_rd_req_desc_c_axid_3_axid
 ,output [31:0] int_rd_req_desc_c_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_c_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_c_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_c_size_txn_size
 ,output [13:0] int_wr_req_desc_c_data_offset_addr
 ,output [2:0] int_wr_req_desc_c_axsize_axsize
 ,output [3:0] int_wr_req_desc_c_attr_axsnoop
 ,output [1:0] int_wr_req_desc_c_attr_axdomain
 ,output [1:0] int_wr_req_desc_c_attr_axbar
 ,output [0:0] int_wr_req_desc_c_attr_awunique
 ,output [3:0] int_wr_req_desc_c_attr_axregion
 ,output [3:0] int_wr_req_desc_c_attr_axqos
 ,output [2:0] int_wr_req_desc_c_attr_axprot
 ,output [3:0] int_wr_req_desc_c_attr_axcache
 ,output [0:0] int_wr_req_desc_c_attr_axlock
 ,output [1:0] int_wr_req_desc_c_attr_axburst
 ,output [31:0] int_wr_req_desc_c_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_c_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_c_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_c_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_c_axid_0_axid
 ,output [31:0] int_wr_req_desc_c_axid_1_axid
 ,output [31:0] int_wr_req_desc_c_axid_2_axid
 ,output [31:0] int_wr_req_desc_c_axid_3_axid
 ,output [31:0] int_wr_req_desc_c_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_c_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_c_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_c_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_c_resp_resp
 ,output [31:0] int_rd_req_desc_d_size_txn_size
 ,output [2:0] int_rd_req_desc_d_axsize_axsize
 ,output [3:0] int_rd_req_desc_d_attr_axsnoop
 ,output [1:0] int_rd_req_desc_d_attr_axdomain
 ,output [1:0] int_rd_req_desc_d_attr_axbar
 ,output [3:0] int_rd_req_desc_d_attr_axregion
 ,output [3:0] int_rd_req_desc_d_attr_axqos
 ,output [2:0] int_rd_req_desc_d_attr_axprot
 ,output [3:0] int_rd_req_desc_d_attr_axcache
 ,output [0:0] int_rd_req_desc_d_attr_axlock
 ,output [1:0] int_rd_req_desc_d_attr_axburst
 ,output [31:0] int_rd_req_desc_d_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_d_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_d_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_d_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_d_axid_0_axid
 ,output [31:0] int_rd_req_desc_d_axid_1_axid
 ,output [31:0] int_rd_req_desc_d_axid_2_axid
 ,output [31:0] int_rd_req_desc_d_axid_3_axid
 ,output [31:0] int_rd_req_desc_d_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_d_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_d_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_d_size_txn_size
 ,output [13:0] int_wr_req_desc_d_data_offset_addr
 ,output [2:0] int_wr_req_desc_d_axsize_axsize
 ,output [3:0] int_wr_req_desc_d_attr_axsnoop
 ,output [1:0] int_wr_req_desc_d_attr_axdomain
 ,output [1:0] int_wr_req_desc_d_attr_axbar
 ,output [0:0] int_wr_req_desc_d_attr_awunique
 ,output [3:0] int_wr_req_desc_d_attr_axregion
 ,output [3:0] int_wr_req_desc_d_attr_axqos
 ,output [2:0] int_wr_req_desc_d_attr_axprot
 ,output [3:0] int_wr_req_desc_d_attr_axcache
 ,output [0:0] int_wr_req_desc_d_attr_axlock
 ,output [1:0] int_wr_req_desc_d_attr_axburst
 ,output [31:0] int_wr_req_desc_d_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_d_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_d_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_d_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_d_axid_0_axid
 ,output [31:0] int_wr_req_desc_d_axid_1_axid
 ,output [31:0] int_wr_req_desc_d_axid_2_axid
 ,output [31:0] int_wr_req_desc_d_axid_3_axid
 ,output [31:0] int_wr_req_desc_d_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_d_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_d_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_d_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_d_resp_resp
 ,output [31:0] int_rd_req_desc_e_size_txn_size
 ,output [2:0] int_rd_req_desc_e_axsize_axsize
 ,output [3:0] int_rd_req_desc_e_attr_axsnoop
 ,output [1:0] int_rd_req_desc_e_attr_axdomain
 ,output [1:0] int_rd_req_desc_e_attr_axbar
 ,output [3:0] int_rd_req_desc_e_attr_axregion
 ,output [3:0] int_rd_req_desc_e_attr_axqos
 ,output [2:0] int_rd_req_desc_e_attr_axprot
 ,output [3:0] int_rd_req_desc_e_attr_axcache
 ,output [0:0] int_rd_req_desc_e_attr_axlock
 ,output [1:0] int_rd_req_desc_e_attr_axburst
 ,output [31:0] int_rd_req_desc_e_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_e_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_e_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_e_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_e_axid_0_axid
 ,output [31:0] int_rd_req_desc_e_axid_1_axid
 ,output [31:0] int_rd_req_desc_e_axid_2_axid
 ,output [31:0] int_rd_req_desc_e_axid_3_axid
 ,output [31:0] int_rd_req_desc_e_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_e_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_e_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_e_size_txn_size
 ,output [13:0] int_wr_req_desc_e_data_offset_addr
 ,output [2:0] int_wr_req_desc_e_axsize_axsize
 ,output [3:0] int_wr_req_desc_e_attr_axsnoop
 ,output [1:0] int_wr_req_desc_e_attr_axdomain
 ,output [1:0] int_wr_req_desc_e_attr_axbar
 ,output [0:0] int_wr_req_desc_e_attr_awunique
 ,output [3:0] int_wr_req_desc_e_attr_axregion
 ,output [3:0] int_wr_req_desc_e_attr_axqos
 ,output [2:0] int_wr_req_desc_e_attr_axprot
 ,output [3:0] int_wr_req_desc_e_attr_axcache
 ,output [0:0] int_wr_req_desc_e_attr_axlock
 ,output [1:0] int_wr_req_desc_e_attr_axburst
 ,output [31:0] int_wr_req_desc_e_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_e_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_e_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_e_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_e_axid_0_axid
 ,output [31:0] int_wr_req_desc_e_axid_1_axid
 ,output [31:0] int_wr_req_desc_e_axid_2_axid
 ,output [31:0] int_wr_req_desc_e_axid_3_axid
 ,output [31:0] int_wr_req_desc_e_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_e_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_e_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_e_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_e_resp_resp
 ,output [31:0] int_rd_req_desc_f_size_txn_size
 ,output [2:0] int_rd_req_desc_f_axsize_axsize
 ,output [3:0] int_rd_req_desc_f_attr_axsnoop
 ,output [1:0] int_rd_req_desc_f_attr_axdomain
 ,output [1:0] int_rd_req_desc_f_attr_axbar
 ,output [3:0] int_rd_req_desc_f_attr_axregion
 ,output [3:0] int_rd_req_desc_f_attr_axqos
 ,output [2:0] int_rd_req_desc_f_attr_axprot
 ,output [3:0] int_rd_req_desc_f_attr_axcache
 ,output [0:0] int_rd_req_desc_f_attr_axlock
 ,output [1:0] int_rd_req_desc_f_attr_axburst
 ,output [31:0] int_rd_req_desc_f_axaddr_0_addr
 ,output [31:0] int_rd_req_desc_f_axaddr_1_addr
 ,output [31:0] int_rd_req_desc_f_axaddr_2_addr
 ,output [31:0] int_rd_req_desc_f_axaddr_3_addr
 ,output [31:0] int_rd_req_desc_f_axid_0_axid
 ,output [31:0] int_rd_req_desc_f_axid_1_axid
 ,output [31:0] int_rd_req_desc_f_axid_2_axid
 ,output [31:0] int_rd_req_desc_f_axid_3_axid
 ,output [31:0] int_rd_req_desc_f_axuser_0_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_1_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_2_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_3_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_4_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_5_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_6_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_7_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_8_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_9_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_10_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_11_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_12_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_13_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_14_axuser
 ,output [31:0] int_rd_req_desc_f_axuser_15_axuser
 ,output [0:0] int_wr_req_desc_f_txn_type_wr_strb
 ,output [31:0] int_wr_req_desc_f_size_txn_size
 ,output [13:0] int_wr_req_desc_f_data_offset_addr
 ,output [2:0] int_wr_req_desc_f_axsize_axsize
 ,output [3:0] int_wr_req_desc_f_attr_axsnoop
 ,output [1:0] int_wr_req_desc_f_attr_axdomain
 ,output [1:0] int_wr_req_desc_f_attr_axbar
 ,output [0:0] int_wr_req_desc_f_attr_awunique
 ,output [3:0] int_wr_req_desc_f_attr_axregion
 ,output [3:0] int_wr_req_desc_f_attr_axqos
 ,output [2:0] int_wr_req_desc_f_attr_axprot
 ,output [3:0] int_wr_req_desc_f_attr_axcache
 ,output [0:0] int_wr_req_desc_f_attr_axlock
 ,output [1:0] int_wr_req_desc_f_attr_axburst
 ,output [31:0] int_wr_req_desc_f_axaddr_0_addr
 ,output [31:0] int_wr_req_desc_f_axaddr_1_addr
 ,output [31:0] int_wr_req_desc_f_axaddr_2_addr
 ,output [31:0] int_wr_req_desc_f_axaddr_3_addr
 ,output [31:0] int_wr_req_desc_f_axid_0_axid
 ,output [31:0] int_wr_req_desc_f_axid_1_axid
 ,output [31:0] int_wr_req_desc_f_axid_2_axid
 ,output [31:0] int_wr_req_desc_f_axid_3_axid
 ,output [31:0] int_wr_req_desc_f_axuser_0_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_1_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_2_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_3_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_4_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_5_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_6_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_7_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_8_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_9_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_10_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_11_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_12_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_13_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_14_axuser
 ,output [31:0] int_wr_req_desc_f_axuser_15_axuser
 ,output [31:0] int_wr_req_desc_f_wuser_0_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_1_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_2_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_3_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_4_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_5_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_6_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_7_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_8_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_9_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_10_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_11_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_12_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_13_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_14_wuser
 ,output [31:0] int_wr_req_desc_f_wuser_15_wuser
 ,output [4:0] int_sn_resp_desc_f_resp_resp

