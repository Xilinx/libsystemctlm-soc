/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Alok Mistry.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 *
 * Description: 
 *   User Master Control is wrapper on top of axi_master_control.
 *
 *
 */

`include "defines_common.vh"
module user_master_control #(
                             parameter M_AXI_USR_ADDR_WIDTH         =    64,    
                             parameter M_AXI_USR_DATA_WIDTH         =    128, //Allowed values : 32,64,128
                             parameter M_AXI_USR_ID_WIDTH           =    16,  //Allowed values : 1-16
			     parameter M_AXI_USR_AWUSER_WIDTH         =    32, //Allowed values : 1-32
			     parameter M_AXI_USR_WUSER_WIDTH         =    32, //Allowed values : 1-32
			     parameter M_AXI_USR_BUSER_WIDTH         =    32, //Allowed values : 1-32
			     parameter M_AXI_USR_ARUSER_WIDTH         =    32, //Allowed values : 1-32
			     parameter M_AXI_USR_RUSER_WIDTH         =    32, //Allowed values : 1-32
                             parameter RAM_SIZE                     =   16384, // Size of RAM in Bytes
                             parameter MAX_DESC                     =   16,                  							 
			     parameter EN_INTFM_AXI4  = 1,
			     parameter EN_INTFM_AXI4LITE = 0,
			     parameter EN_INTFM_AXI3 = 0

                             )
   (



    input 						     axi_aclk,
    input 						     axi_aresetn,
   
    // Data Ram Interface 
    //read port of WR DataRam
    output [(`CLOG2(RAM_SIZE/(M_AXI_USR_DATA_WIDTH/8)))-1:0] uc2rb_rd_addr, //Currently, [10:0]
    input [M_AXI_USR_DATA_WIDTH-1:0] 			     rb2uc_rd_data,
    input [(M_AXI_USR_DATA_WIDTH/8 -1):0] 		     rb2uc_rd_wstrb, 
    // Write port of RD DataRam
    output 						     uc2rb_wr_we, 
    output [(M_AXI_USR_DATA_WIDTH/8 -1):0] 		     uc2rb_wr_bwe, 
    //    output [(`CLOG2(RAM_SIZE/(M_AXI_USR_DATA_WIDTH/8)))-1:0] uc2rb_wr_addr, //Currently, [10:0]
    output [(`CLOG2(RAM_SIZE/(M_AXI_USR_DATA_WIDTH/8)))-1:0] uc2rb_wr_addr, //Currently, [10:0]
    output [M_AXI_USR_DATA_WIDTH-1:0] 			     uc2rb_wr_data, 

    //Host Master Interface (Mode 1)
    output [15:0] 					     uc2hm_trig,
    input [15:0] 					     hm2uc_done,
   
    // Registers from Block
    input [31:0] 					     version_reg ,
    input [31:0] 					     bridge_type_reg ,
    input [31:0] 					     mode_select_reg ,
    input [31:0] 					     reset_reg ,
    input [31:0] 					     intr_h2c_0_reg ,
    input [31:0] 					     intr_h2c_1_reg ,
    input [31:0] 					     intr_c2h_0_status_reg ,
    input [31:0] 					     intr_c2h_1_status_reg ,
    input [31:0] 					     c2h_gpio_0_status_reg ,
    input [31:0] 					     c2h_gpio_1_status_reg ,
    input [31:0] 					     c2h_gpio_2_status_reg ,
    input [31:0] 					     c2h_gpio_3_status_reg ,
    input [31:0] 					     c2h_gpio_4_status_reg ,
    input [31:0] 					     c2h_gpio_5_status_reg ,
    input [31:0] 					     c2h_gpio_6_status_reg ,
    input [31:0] 					     c2h_gpio_7_status_reg ,
    input [31:0] 					     c2h_gpio_8_status_reg ,
    input [31:0] 					     c2h_gpio_9_status_reg ,
    input [31:0] 					     c2h_gpio_10_status_reg ,
    input [31:0] 					     c2h_gpio_11_status_reg ,
    input [31:0] 					     c2h_gpio_12_status_reg ,
    input [31:0] 					     c2h_gpio_13_status_reg ,
    input [31:0] 					     c2h_gpio_14_status_reg ,
    input [31:0] 					     c2h_gpio_15_status_reg ,
    input [31:0] 					     axi_bridge_config_reg ,
    input [31:0] 					     axi_max_desc_reg ,
    input [31:0] 					     intr_status_reg ,
    input [31:0] 					     intr_error_status_reg ,
    input [31:0] 					     intr_error_clear_reg ,
    input [31:0] 					     intr_error_enable_reg ,
    input [31:0] 					     ownership_reg ,
    input [31:0] 					     ownership_flip_reg ,
    input [31:0] 					     status_resp_reg ,
    input [31:0] 					     intr_comp_status_reg ,
    input [31:0] 					     intr_comp_clear_reg ,
    input [31:0] 					     intr_comp_enable_reg ,
    input [31:0] 					     desc_0_txn_type_reg ,
    input [31:0] 					     desc_0_size_reg ,
    input [31:0] 					     desc_0_data_offset_reg ,
    input [31:0] 					     desc_0_data_host_addr_0_reg ,
    input [31:0] 					     desc_0_data_host_addr_1_reg ,
    input [31:0] 					     desc_0_data_host_addr_2_reg ,
    input [31:0] 					     desc_0_data_host_addr_3_reg ,
    input [31:0] 					     desc_0_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_0_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_0_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_0_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_0_axsize_reg ,
    input [31:0] 					     desc_0_attr_reg ,
    input [31:0] 					     desc_0_axaddr_0_reg ,
    input [31:0] 					     desc_0_axaddr_1_reg ,
    input [31:0] 					     desc_0_axaddr_2_reg ,
    input [31:0] 					     desc_0_axaddr_3_reg ,
    input [31:0] 					     desc_0_axid_0_reg ,
    input [31:0] 					     desc_0_axid_1_reg ,
    input [31:0] 					     desc_0_axid_2_reg ,
    input [31:0] 					     desc_0_axid_3_reg ,
    input [31:0] 					     desc_0_axuser_0_reg ,
    input [31:0] 					     desc_0_axuser_1_reg ,
    input [31:0] 					     desc_0_axuser_2_reg ,
    input [31:0] 					     desc_0_axuser_3_reg ,
    input [31:0] 					     desc_0_axuser_4_reg ,
    input [31:0] 					     desc_0_axuser_5_reg ,
    input [31:0] 					     desc_0_axuser_6_reg ,
    input [31:0] 					     desc_0_axuser_7_reg ,
    input [31:0] 					     desc_0_axuser_8_reg ,
    input [31:0] 					     desc_0_axuser_9_reg ,
    input [31:0] 					     desc_0_axuser_10_reg ,
    input [31:0] 					     desc_0_axuser_11_reg ,
    input [31:0] 					     desc_0_axuser_12_reg ,
    input [31:0] 					     desc_0_axuser_13_reg ,
    input [31:0] 					     desc_0_axuser_14_reg ,
    input [31:0] 					     desc_0_axuser_15_reg ,
    input [31:0] 					     desc_0_xuser_0_reg ,
    input [31:0] 					     desc_0_xuser_1_reg ,
    input [31:0] 					     desc_0_xuser_2_reg ,
    input [31:0] 					     desc_0_xuser_3_reg ,
    input [31:0] 					     desc_0_xuser_4_reg ,
    input [31:0] 					     desc_0_xuser_5_reg ,
    input [31:0] 					     desc_0_xuser_6_reg ,
    input [31:0] 					     desc_0_xuser_7_reg ,
    input [31:0] 					     desc_0_xuser_8_reg ,
    input [31:0] 					     desc_0_xuser_9_reg ,
    input [31:0] 					     desc_0_xuser_10_reg ,
    input [31:0] 					     desc_0_xuser_11_reg ,
    input [31:0] 					     desc_0_xuser_12_reg ,
    input [31:0] 					     desc_0_xuser_13_reg ,
    input [31:0] 					     desc_0_xuser_14_reg ,
    input [31:0] 					     desc_0_xuser_15_reg ,
    input [31:0] 					     desc_0_wuser_0_reg ,
    input [31:0] 					     desc_0_wuser_1_reg ,
    input [31:0] 					     desc_0_wuser_2_reg ,
    input [31:0] 					     desc_0_wuser_3_reg ,
    input [31:0] 					     desc_0_wuser_4_reg ,
    input [31:0] 					     desc_0_wuser_5_reg ,
    input [31:0] 					     desc_0_wuser_6_reg ,
    input [31:0] 					     desc_0_wuser_7_reg ,
    input [31:0] 					     desc_0_wuser_8_reg ,
    input [31:0] 					     desc_0_wuser_9_reg ,
    input [31:0] 					     desc_0_wuser_10_reg ,
    input [31:0] 					     desc_0_wuser_11_reg ,
    input [31:0] 					     desc_0_wuser_12_reg ,
    input [31:0] 					     desc_0_wuser_13_reg ,
    input [31:0] 					     desc_0_wuser_14_reg ,
    input [31:0] 					     desc_0_wuser_15_reg ,
    input [31:0] 					     desc_1_txn_type_reg ,
    input [31:0] 					     desc_1_size_reg ,
    input [31:0] 					     desc_1_data_offset_reg ,
    input [31:0] 					     desc_1_data_host_addr_0_reg ,
    input [31:0] 					     desc_1_data_host_addr_1_reg ,
    input [31:0] 					     desc_1_data_host_addr_2_reg ,
    input [31:0] 					     desc_1_data_host_addr_3_reg ,
    input [31:0] 					     desc_1_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_1_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_1_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_1_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_1_axsize_reg ,
    input [31:0] 					     desc_1_attr_reg ,
    input [31:0] 					     desc_1_axaddr_0_reg ,
    input [31:0] 					     desc_1_axaddr_1_reg ,
    input [31:0] 					     desc_1_axaddr_2_reg ,
    input [31:0] 					     desc_1_axaddr_3_reg ,
    input [31:0] 					     desc_1_axid_0_reg ,
    input [31:0] 					     desc_1_axid_1_reg ,
    input [31:0] 					     desc_1_axid_2_reg ,
    input [31:0] 					     desc_1_axid_3_reg ,
    input [31:0] 					     desc_1_axuser_0_reg ,
    input [31:0] 					     desc_1_axuser_1_reg ,
    input [31:0] 					     desc_1_axuser_2_reg ,
    input [31:0] 					     desc_1_axuser_3_reg ,
    input [31:0] 					     desc_1_axuser_4_reg ,
    input [31:0] 					     desc_1_axuser_5_reg ,
    input [31:0] 					     desc_1_axuser_6_reg ,
    input [31:0] 					     desc_1_axuser_7_reg ,
    input [31:0] 					     desc_1_axuser_8_reg ,
    input [31:0] 					     desc_1_axuser_9_reg ,
    input [31:0] 					     desc_1_axuser_10_reg ,
    input [31:0] 					     desc_1_axuser_11_reg ,
    input [31:0] 					     desc_1_axuser_12_reg ,
    input [31:0] 					     desc_1_axuser_13_reg ,
    input [31:0] 					     desc_1_axuser_14_reg ,
    input [31:0] 					     desc_1_axuser_15_reg ,
    input [31:0] 					     desc_1_xuser_0_reg ,
    input [31:0] 					     desc_1_xuser_1_reg ,
    input [31:0] 					     desc_1_xuser_2_reg ,
    input [31:0] 					     desc_1_xuser_3_reg ,
    input [31:0] 					     desc_1_xuser_4_reg ,
    input [31:0] 					     desc_1_xuser_5_reg ,
    input [31:0] 					     desc_1_xuser_6_reg ,
    input [31:0] 					     desc_1_xuser_7_reg ,
    input [31:0] 					     desc_1_xuser_8_reg ,
    input [31:0] 					     desc_1_xuser_9_reg ,
    input [31:0] 					     desc_1_xuser_10_reg ,
    input [31:0] 					     desc_1_xuser_11_reg ,
    input [31:0] 					     desc_1_xuser_12_reg ,
    input [31:0] 					     desc_1_xuser_13_reg ,
    input [31:0] 					     desc_1_xuser_14_reg ,
    input [31:0] 					     desc_1_xuser_15_reg ,
    input [31:0] 					     desc_1_wuser_0_reg ,
    input [31:0] 					     desc_1_wuser_1_reg ,
    input [31:0] 					     desc_1_wuser_2_reg ,
    input [31:0] 					     desc_1_wuser_3_reg ,
    input [31:0] 					     desc_1_wuser_4_reg ,
    input [31:0] 					     desc_1_wuser_5_reg ,
    input [31:0] 					     desc_1_wuser_6_reg ,
    input [31:0] 					     desc_1_wuser_7_reg ,
    input [31:0] 					     desc_1_wuser_8_reg ,
    input [31:0] 					     desc_1_wuser_9_reg ,
    input [31:0] 					     desc_1_wuser_10_reg ,
    input [31:0] 					     desc_1_wuser_11_reg ,
    input [31:0] 					     desc_1_wuser_12_reg ,
    input [31:0] 					     desc_1_wuser_13_reg ,
    input [31:0] 					     desc_1_wuser_14_reg ,
    input [31:0] 					     desc_1_wuser_15_reg ,
    input [31:0] 					     desc_2_txn_type_reg ,
    input [31:0] 					     desc_2_size_reg ,
    input [31:0] 					     desc_2_data_offset_reg ,
    input [31:0] 					     desc_2_data_host_addr_0_reg ,
    input [31:0] 					     desc_2_data_host_addr_1_reg ,
    input [31:0] 					     desc_2_data_host_addr_2_reg ,
    input [31:0] 					     desc_2_data_host_addr_3_reg ,
    input [31:0] 					     desc_2_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_2_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_2_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_2_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_2_axsize_reg ,
    input [31:0] 					     desc_2_attr_reg ,
    input [31:0] 					     desc_2_axaddr_0_reg ,
    input [31:0] 					     desc_2_axaddr_1_reg ,
    input [31:0] 					     desc_2_axaddr_2_reg ,
    input [31:0] 					     desc_2_axaddr_3_reg ,
    input [31:0] 					     desc_2_axid_0_reg ,
    input [31:0] 					     desc_2_axid_1_reg ,
    input [31:0] 					     desc_2_axid_2_reg ,
    input [31:0] 					     desc_2_axid_3_reg ,
    input [31:0] 					     desc_2_axuser_0_reg ,
    input [31:0] 					     desc_2_axuser_1_reg ,
    input [31:0] 					     desc_2_axuser_2_reg ,
    input [31:0] 					     desc_2_axuser_3_reg ,
    input [31:0] 					     desc_2_axuser_4_reg ,
    input [31:0] 					     desc_2_axuser_5_reg ,
    input [31:0] 					     desc_2_axuser_6_reg ,
    input [31:0] 					     desc_2_axuser_7_reg ,
    input [31:0] 					     desc_2_axuser_8_reg ,
    input [31:0] 					     desc_2_axuser_9_reg ,
    input [31:0] 					     desc_2_axuser_10_reg ,
    input [31:0] 					     desc_2_axuser_11_reg ,
    input [31:0] 					     desc_2_axuser_12_reg ,
    input [31:0] 					     desc_2_axuser_13_reg ,
    input [31:0] 					     desc_2_axuser_14_reg ,
    input [31:0] 					     desc_2_axuser_15_reg ,
    input [31:0] 					     desc_2_xuser_0_reg ,
    input [31:0] 					     desc_2_xuser_1_reg ,
    input [31:0] 					     desc_2_xuser_2_reg ,
    input [31:0] 					     desc_2_xuser_3_reg ,
    input [31:0] 					     desc_2_xuser_4_reg ,
    input [31:0] 					     desc_2_xuser_5_reg ,
    input [31:0] 					     desc_2_xuser_6_reg ,
    input [31:0] 					     desc_2_xuser_7_reg ,
    input [31:0] 					     desc_2_xuser_8_reg ,
    input [31:0] 					     desc_2_xuser_9_reg ,
    input [31:0] 					     desc_2_xuser_10_reg ,
    input [31:0] 					     desc_2_xuser_11_reg ,
    input [31:0] 					     desc_2_xuser_12_reg ,
    input [31:0] 					     desc_2_xuser_13_reg ,
    input [31:0] 					     desc_2_xuser_14_reg ,
    input [31:0] 					     desc_2_xuser_15_reg ,
    input [31:0] 					     desc_2_wuser_0_reg ,
    input [31:0] 					     desc_2_wuser_1_reg ,
    input [31:0] 					     desc_2_wuser_2_reg ,
    input [31:0] 					     desc_2_wuser_3_reg ,
    input [31:0] 					     desc_2_wuser_4_reg ,
    input [31:0] 					     desc_2_wuser_5_reg ,
    input [31:0] 					     desc_2_wuser_6_reg ,
    input [31:0] 					     desc_2_wuser_7_reg ,
    input [31:0] 					     desc_2_wuser_8_reg ,
    input [31:0] 					     desc_2_wuser_9_reg ,
    input [31:0] 					     desc_2_wuser_10_reg ,
    input [31:0] 					     desc_2_wuser_11_reg ,
    input [31:0] 					     desc_2_wuser_12_reg ,
    input [31:0] 					     desc_2_wuser_13_reg ,
    input [31:0] 					     desc_2_wuser_14_reg ,
    input [31:0] 					     desc_2_wuser_15_reg ,
    input [31:0] 					     desc_3_txn_type_reg ,
    input [31:0] 					     desc_3_size_reg ,
    input [31:0] 					     desc_3_data_offset_reg ,
    input [31:0] 					     desc_3_data_host_addr_0_reg ,
    input [31:0] 					     desc_3_data_host_addr_1_reg ,
    input [31:0] 					     desc_3_data_host_addr_2_reg ,
    input [31:0] 					     desc_3_data_host_addr_3_reg ,
    input [31:0] 					     desc_3_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_3_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_3_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_3_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_3_axsize_reg ,
    input [31:0] 					     desc_3_attr_reg ,
    input [31:0] 					     desc_3_axaddr_0_reg ,
    input [31:0] 					     desc_3_axaddr_1_reg ,
    input [31:0] 					     desc_3_axaddr_2_reg ,
    input [31:0] 					     desc_3_axaddr_3_reg ,
    input [31:0] 					     desc_3_axid_0_reg ,
    input [31:0] 					     desc_3_axid_1_reg ,
    input [31:0] 					     desc_3_axid_2_reg ,
    input [31:0] 					     desc_3_axid_3_reg ,
    input [31:0] 					     desc_3_axuser_0_reg ,
    input [31:0] 					     desc_3_axuser_1_reg ,
    input [31:0] 					     desc_3_axuser_2_reg ,
    input [31:0] 					     desc_3_axuser_3_reg ,
    input [31:0] 					     desc_3_axuser_4_reg ,
    input [31:0] 					     desc_3_axuser_5_reg ,
    input [31:0] 					     desc_3_axuser_6_reg ,
    input [31:0] 					     desc_3_axuser_7_reg ,
    input [31:0] 					     desc_3_axuser_8_reg ,
    input [31:0] 					     desc_3_axuser_9_reg ,
    input [31:0] 					     desc_3_axuser_10_reg ,
    input [31:0] 					     desc_3_axuser_11_reg ,
    input [31:0] 					     desc_3_axuser_12_reg ,
    input [31:0] 					     desc_3_axuser_13_reg ,
    input [31:0] 					     desc_3_axuser_14_reg ,
    input [31:0] 					     desc_3_axuser_15_reg ,
    input [31:0] 					     desc_3_xuser_0_reg ,
    input [31:0] 					     desc_3_xuser_1_reg ,
    input [31:0] 					     desc_3_xuser_2_reg ,
    input [31:0] 					     desc_3_xuser_3_reg ,
    input [31:0] 					     desc_3_xuser_4_reg ,
    input [31:0] 					     desc_3_xuser_5_reg ,
    input [31:0] 					     desc_3_xuser_6_reg ,
    input [31:0] 					     desc_3_xuser_7_reg ,
    input [31:0] 					     desc_3_xuser_8_reg ,
    input [31:0] 					     desc_3_xuser_9_reg ,
    input [31:0] 					     desc_3_xuser_10_reg ,
    input [31:0] 					     desc_3_xuser_11_reg ,
    input [31:0] 					     desc_3_xuser_12_reg ,
    input [31:0] 					     desc_3_xuser_13_reg ,
    input [31:0] 					     desc_3_xuser_14_reg ,
    input [31:0] 					     desc_3_xuser_15_reg ,
    input [31:0] 					     desc_3_wuser_0_reg ,
    input [31:0] 					     desc_3_wuser_1_reg ,
    input [31:0] 					     desc_3_wuser_2_reg ,
    input [31:0] 					     desc_3_wuser_3_reg ,
    input [31:0] 					     desc_3_wuser_4_reg ,
    input [31:0] 					     desc_3_wuser_5_reg ,
    input [31:0] 					     desc_3_wuser_6_reg ,
    input [31:0] 					     desc_3_wuser_7_reg ,
    input [31:0] 					     desc_3_wuser_8_reg ,
    input [31:0] 					     desc_3_wuser_9_reg ,
    input [31:0] 					     desc_3_wuser_10_reg ,
    input [31:0] 					     desc_3_wuser_11_reg ,
    input [31:0] 					     desc_3_wuser_12_reg ,
    input [31:0] 					     desc_3_wuser_13_reg ,
    input [31:0] 					     desc_3_wuser_14_reg ,
    input [31:0] 					     desc_3_wuser_15_reg ,
    input [31:0] 					     desc_4_txn_type_reg ,
    input [31:0] 					     desc_4_size_reg ,
    input [31:0] 					     desc_4_data_offset_reg ,
    input [31:0] 					     desc_4_data_host_addr_0_reg ,
    input [31:0] 					     desc_4_data_host_addr_1_reg ,
    input [31:0] 					     desc_4_data_host_addr_2_reg ,
    input [31:0] 					     desc_4_data_host_addr_3_reg ,
    input [31:0] 					     desc_4_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_4_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_4_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_4_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_4_axsize_reg ,
    input [31:0] 					     desc_4_attr_reg ,
    input [31:0] 					     desc_4_axaddr_0_reg ,
    input [31:0] 					     desc_4_axaddr_1_reg ,
    input [31:0] 					     desc_4_axaddr_2_reg ,
    input [31:0] 					     desc_4_axaddr_3_reg ,
    input [31:0] 					     desc_4_axid_0_reg ,
    input [31:0] 					     desc_4_axid_1_reg ,
    input [31:0] 					     desc_4_axid_2_reg ,
    input [31:0] 					     desc_4_axid_3_reg ,
    input [31:0] 					     desc_4_axuser_0_reg ,
    input [31:0] 					     desc_4_axuser_1_reg ,
    input [31:0] 					     desc_4_axuser_2_reg ,
    input [31:0] 					     desc_4_axuser_3_reg ,
    input [31:0] 					     desc_4_axuser_4_reg ,
    input [31:0] 					     desc_4_axuser_5_reg ,
    input [31:0] 					     desc_4_axuser_6_reg ,
    input [31:0] 					     desc_4_axuser_7_reg ,
    input [31:0] 					     desc_4_axuser_8_reg ,
    input [31:0] 					     desc_4_axuser_9_reg ,
    input [31:0] 					     desc_4_axuser_10_reg ,
    input [31:0] 					     desc_4_axuser_11_reg ,
    input [31:0] 					     desc_4_axuser_12_reg ,
    input [31:0] 					     desc_4_axuser_13_reg ,
    input [31:0] 					     desc_4_axuser_14_reg ,
    input [31:0] 					     desc_4_axuser_15_reg ,
    input [31:0] 					     desc_4_xuser_0_reg ,
    input [31:0] 					     desc_4_xuser_1_reg ,
    input [31:0] 					     desc_4_xuser_2_reg ,
    input [31:0] 					     desc_4_xuser_3_reg ,
    input [31:0] 					     desc_4_xuser_4_reg ,
    input [31:0] 					     desc_4_xuser_5_reg ,
    input [31:0] 					     desc_4_xuser_6_reg ,
    input [31:0] 					     desc_4_xuser_7_reg ,
    input [31:0] 					     desc_4_xuser_8_reg ,
    input [31:0] 					     desc_4_xuser_9_reg ,
    input [31:0] 					     desc_4_xuser_10_reg ,
    input [31:0] 					     desc_4_xuser_11_reg ,
    input [31:0] 					     desc_4_xuser_12_reg ,
    input [31:0] 					     desc_4_xuser_13_reg ,
    input [31:0] 					     desc_4_xuser_14_reg ,
    input [31:0] 					     desc_4_xuser_15_reg ,
    input [31:0] 					     desc_4_wuser_0_reg ,
    input [31:0] 					     desc_4_wuser_1_reg ,
    input [31:0] 					     desc_4_wuser_2_reg ,
    input [31:0] 					     desc_4_wuser_3_reg ,
    input [31:0] 					     desc_4_wuser_4_reg ,
    input [31:0] 					     desc_4_wuser_5_reg ,
    input [31:0] 					     desc_4_wuser_6_reg ,
    input [31:0] 					     desc_4_wuser_7_reg ,
    input [31:0] 					     desc_4_wuser_8_reg ,
    input [31:0] 					     desc_4_wuser_9_reg ,
    input [31:0] 					     desc_4_wuser_10_reg ,
    input [31:0] 					     desc_4_wuser_11_reg ,
    input [31:0] 					     desc_4_wuser_12_reg ,
    input [31:0] 					     desc_4_wuser_13_reg ,
    input [31:0] 					     desc_4_wuser_14_reg ,
    input [31:0] 					     desc_4_wuser_15_reg ,
    input [31:0] 					     desc_5_txn_type_reg ,
    input [31:0] 					     desc_5_size_reg ,
    input [31:0] 					     desc_5_data_offset_reg ,
    input [31:0] 					     desc_5_data_host_addr_0_reg ,
    input [31:0] 					     desc_5_data_host_addr_1_reg ,
    input [31:0] 					     desc_5_data_host_addr_2_reg ,
    input [31:0] 					     desc_5_data_host_addr_3_reg ,
    input [31:0] 					     desc_5_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_5_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_5_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_5_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_5_axsize_reg ,
    input [31:0] 					     desc_5_attr_reg ,
    input [31:0] 					     desc_5_axaddr_0_reg ,
    input [31:0] 					     desc_5_axaddr_1_reg ,
    input [31:0] 					     desc_5_axaddr_2_reg ,
    input [31:0] 					     desc_5_axaddr_3_reg ,
    input [31:0] 					     desc_5_axid_0_reg ,
    input [31:0] 					     desc_5_axid_1_reg ,
    input [31:0] 					     desc_5_axid_2_reg ,
    input [31:0] 					     desc_5_axid_3_reg ,
    input [31:0] 					     desc_5_axuser_0_reg ,
    input [31:0] 					     desc_5_axuser_1_reg ,
    input [31:0] 					     desc_5_axuser_2_reg ,
    input [31:0] 					     desc_5_axuser_3_reg ,
    input [31:0] 					     desc_5_axuser_4_reg ,
    input [31:0] 					     desc_5_axuser_5_reg ,
    input [31:0] 					     desc_5_axuser_6_reg ,
    input [31:0] 					     desc_5_axuser_7_reg ,
    input [31:0] 					     desc_5_axuser_8_reg ,
    input [31:0] 					     desc_5_axuser_9_reg ,
    input [31:0] 					     desc_5_axuser_10_reg ,
    input [31:0] 					     desc_5_axuser_11_reg ,
    input [31:0] 					     desc_5_axuser_12_reg ,
    input [31:0] 					     desc_5_axuser_13_reg ,
    input [31:0] 					     desc_5_axuser_14_reg ,
    input [31:0] 					     desc_5_axuser_15_reg ,
    input [31:0] 					     desc_5_xuser_0_reg ,
    input [31:0] 					     desc_5_xuser_1_reg ,
    input [31:0] 					     desc_5_xuser_2_reg ,
    input [31:0] 					     desc_5_xuser_3_reg ,
    input [31:0] 					     desc_5_xuser_4_reg ,
    input [31:0] 					     desc_5_xuser_5_reg ,
    input [31:0] 					     desc_5_xuser_6_reg ,
    input [31:0] 					     desc_5_xuser_7_reg ,
    input [31:0] 					     desc_5_xuser_8_reg ,
    input [31:0] 					     desc_5_xuser_9_reg ,
    input [31:0] 					     desc_5_xuser_10_reg ,
    input [31:0] 					     desc_5_xuser_11_reg ,
    input [31:0] 					     desc_5_xuser_12_reg ,
    input [31:0] 					     desc_5_xuser_13_reg ,
    input [31:0] 					     desc_5_xuser_14_reg ,
    input [31:0] 					     desc_5_xuser_15_reg ,
    input [31:0] 					     desc_5_wuser_0_reg ,
    input [31:0] 					     desc_5_wuser_1_reg ,
    input [31:0] 					     desc_5_wuser_2_reg ,
    input [31:0] 					     desc_5_wuser_3_reg ,
    input [31:0] 					     desc_5_wuser_4_reg ,
    input [31:0] 					     desc_5_wuser_5_reg ,
    input [31:0] 					     desc_5_wuser_6_reg ,
    input [31:0] 					     desc_5_wuser_7_reg ,
    input [31:0] 					     desc_5_wuser_8_reg ,
    input [31:0] 					     desc_5_wuser_9_reg ,
    input [31:0] 					     desc_5_wuser_10_reg ,
    input [31:0] 					     desc_5_wuser_11_reg ,
    input [31:0] 					     desc_5_wuser_12_reg ,
    input [31:0] 					     desc_5_wuser_13_reg ,
    input [31:0] 					     desc_5_wuser_14_reg ,
    input [31:0] 					     desc_5_wuser_15_reg ,
    input [31:0] 					     desc_6_txn_type_reg ,
    input [31:0] 					     desc_6_size_reg ,
    input [31:0] 					     desc_6_data_offset_reg ,
    input [31:0] 					     desc_6_data_host_addr_0_reg ,
    input [31:0] 					     desc_6_data_host_addr_1_reg ,
    input [31:0] 					     desc_6_data_host_addr_2_reg ,
    input [31:0] 					     desc_6_data_host_addr_3_reg ,
    input [31:0] 					     desc_6_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_6_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_6_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_6_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_6_axsize_reg ,
    input [31:0] 					     desc_6_attr_reg ,
    input [31:0] 					     desc_6_axaddr_0_reg ,
    input [31:0] 					     desc_6_axaddr_1_reg ,
    input [31:0] 					     desc_6_axaddr_2_reg ,
    input [31:0] 					     desc_6_axaddr_3_reg ,
    input [31:0] 					     desc_6_axid_0_reg ,
    input [31:0] 					     desc_6_axid_1_reg ,
    input [31:0] 					     desc_6_axid_2_reg ,
    input [31:0] 					     desc_6_axid_3_reg ,
    input [31:0] 					     desc_6_axuser_0_reg ,
    input [31:0] 					     desc_6_axuser_1_reg ,
    input [31:0] 					     desc_6_axuser_2_reg ,
    input [31:0] 					     desc_6_axuser_3_reg ,
    input [31:0] 					     desc_6_axuser_4_reg ,
    input [31:0] 					     desc_6_axuser_5_reg ,
    input [31:0] 					     desc_6_axuser_6_reg ,
    input [31:0] 					     desc_6_axuser_7_reg ,
    input [31:0] 					     desc_6_axuser_8_reg ,
    input [31:0] 					     desc_6_axuser_9_reg ,
    input [31:0] 					     desc_6_axuser_10_reg ,
    input [31:0] 					     desc_6_axuser_11_reg ,
    input [31:0] 					     desc_6_axuser_12_reg ,
    input [31:0] 					     desc_6_axuser_13_reg ,
    input [31:0] 					     desc_6_axuser_14_reg ,
    input [31:0] 					     desc_6_axuser_15_reg ,
    input [31:0] 					     desc_6_xuser_0_reg ,
    input [31:0] 					     desc_6_xuser_1_reg ,
    input [31:0] 					     desc_6_xuser_2_reg ,
    input [31:0] 					     desc_6_xuser_3_reg ,
    input [31:0] 					     desc_6_xuser_4_reg ,
    input [31:0] 					     desc_6_xuser_5_reg ,
    input [31:0] 					     desc_6_xuser_6_reg ,
    input [31:0] 					     desc_6_xuser_7_reg ,
    input [31:0] 					     desc_6_xuser_8_reg ,
    input [31:0] 					     desc_6_xuser_9_reg ,
    input [31:0] 					     desc_6_xuser_10_reg ,
    input [31:0] 					     desc_6_xuser_11_reg ,
    input [31:0] 					     desc_6_xuser_12_reg ,
    input [31:0] 					     desc_6_xuser_13_reg ,
    input [31:0] 					     desc_6_xuser_14_reg ,
    input [31:0] 					     desc_6_xuser_15_reg ,
    input [31:0] 					     desc_6_wuser_0_reg ,
    input [31:0] 					     desc_6_wuser_1_reg ,
    input [31:0] 					     desc_6_wuser_2_reg ,
    input [31:0] 					     desc_6_wuser_3_reg ,
    input [31:0] 					     desc_6_wuser_4_reg ,
    input [31:0] 					     desc_6_wuser_5_reg ,
    input [31:0] 					     desc_6_wuser_6_reg ,
    input [31:0] 					     desc_6_wuser_7_reg ,
    input [31:0] 					     desc_6_wuser_8_reg ,
    input [31:0] 					     desc_6_wuser_9_reg ,
    input [31:0] 					     desc_6_wuser_10_reg ,
    input [31:0] 					     desc_6_wuser_11_reg ,
    input [31:0] 					     desc_6_wuser_12_reg ,
    input [31:0] 					     desc_6_wuser_13_reg ,
    input [31:0] 					     desc_6_wuser_14_reg ,
    input [31:0] 					     desc_6_wuser_15_reg ,
    input [31:0] 					     desc_7_txn_type_reg ,
    input [31:0] 					     desc_7_size_reg ,
    input [31:0] 					     desc_7_data_offset_reg ,
    input [31:0] 					     desc_7_data_host_addr_0_reg ,
    input [31:0] 					     desc_7_data_host_addr_1_reg ,
    input [31:0] 					     desc_7_data_host_addr_2_reg ,
    input [31:0] 					     desc_7_data_host_addr_3_reg ,
    input [31:0] 					     desc_7_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_7_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_7_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_7_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_7_axsize_reg ,
    input [31:0] 					     desc_7_attr_reg ,
    input [31:0] 					     desc_7_axaddr_0_reg ,
    input [31:0] 					     desc_7_axaddr_1_reg ,
    input [31:0] 					     desc_7_axaddr_2_reg ,
    input [31:0] 					     desc_7_axaddr_3_reg ,
    input [31:0] 					     desc_7_axid_0_reg ,
    input [31:0] 					     desc_7_axid_1_reg ,
    input [31:0] 					     desc_7_axid_2_reg ,
    input [31:0] 					     desc_7_axid_3_reg ,
    input [31:0] 					     desc_7_axuser_0_reg ,
    input [31:0] 					     desc_7_axuser_1_reg ,
    input [31:0] 					     desc_7_axuser_2_reg ,
    input [31:0] 					     desc_7_axuser_3_reg ,
    input [31:0] 					     desc_7_axuser_4_reg ,
    input [31:0] 					     desc_7_axuser_5_reg ,
    input [31:0] 					     desc_7_axuser_6_reg ,
    input [31:0] 					     desc_7_axuser_7_reg ,
    input [31:0] 					     desc_7_axuser_8_reg ,
    input [31:0] 					     desc_7_axuser_9_reg ,
    input [31:0] 					     desc_7_axuser_10_reg ,
    input [31:0] 					     desc_7_axuser_11_reg ,
    input [31:0] 					     desc_7_axuser_12_reg ,
    input [31:0] 					     desc_7_axuser_13_reg ,
    input [31:0] 					     desc_7_axuser_14_reg ,
    input [31:0] 					     desc_7_axuser_15_reg ,
    input [31:0] 					     desc_7_xuser_0_reg ,
    input [31:0] 					     desc_7_xuser_1_reg ,
    input [31:0] 					     desc_7_xuser_2_reg ,
    input [31:0] 					     desc_7_xuser_3_reg ,
    input [31:0] 					     desc_7_xuser_4_reg ,
    input [31:0] 					     desc_7_xuser_5_reg ,
    input [31:0] 					     desc_7_xuser_6_reg ,
    input [31:0] 					     desc_7_xuser_7_reg ,
    input [31:0] 					     desc_7_xuser_8_reg ,
    input [31:0] 					     desc_7_xuser_9_reg ,
    input [31:0] 					     desc_7_xuser_10_reg ,
    input [31:0] 					     desc_7_xuser_11_reg ,
    input [31:0] 					     desc_7_xuser_12_reg ,
    input [31:0] 					     desc_7_xuser_13_reg ,
    input [31:0] 					     desc_7_xuser_14_reg ,
    input [31:0] 					     desc_7_xuser_15_reg ,
    input [31:0] 					     desc_7_wuser_0_reg ,
    input [31:0] 					     desc_7_wuser_1_reg ,
    input [31:0] 					     desc_7_wuser_2_reg ,
    input [31:0] 					     desc_7_wuser_3_reg ,
    input [31:0] 					     desc_7_wuser_4_reg ,
    input [31:0] 					     desc_7_wuser_5_reg ,
    input [31:0] 					     desc_7_wuser_6_reg ,
    input [31:0] 					     desc_7_wuser_7_reg ,
    input [31:0] 					     desc_7_wuser_8_reg ,
    input [31:0] 					     desc_7_wuser_9_reg ,
    input [31:0] 					     desc_7_wuser_10_reg ,
    input [31:0] 					     desc_7_wuser_11_reg ,
    input [31:0] 					     desc_7_wuser_12_reg ,
    input [31:0] 					     desc_7_wuser_13_reg ,
    input [31:0] 					     desc_7_wuser_14_reg ,
    input [31:0] 					     desc_7_wuser_15_reg ,
    input [31:0] 					     desc_8_txn_type_reg ,
    input [31:0] 					     desc_8_size_reg ,
    input [31:0] 					     desc_8_data_offset_reg ,
    input [31:0] 					     desc_8_data_host_addr_0_reg ,
    input [31:0] 					     desc_8_data_host_addr_1_reg ,
    input [31:0] 					     desc_8_data_host_addr_2_reg ,
    input [31:0] 					     desc_8_data_host_addr_3_reg ,
    input [31:0] 					     desc_8_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_8_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_8_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_8_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_8_axsize_reg ,
    input [31:0] 					     desc_8_attr_reg ,
    input [31:0] 					     desc_8_axaddr_0_reg ,
    input [31:0] 					     desc_8_axaddr_1_reg ,
    input [31:0] 					     desc_8_axaddr_2_reg ,
    input [31:0] 					     desc_8_axaddr_3_reg ,
    input [31:0] 					     desc_8_axid_0_reg ,
    input [31:0] 					     desc_8_axid_1_reg ,
    input [31:0] 					     desc_8_axid_2_reg ,
    input [31:0] 					     desc_8_axid_3_reg ,
    input [31:0] 					     desc_8_axuser_0_reg ,
    input [31:0] 					     desc_8_axuser_1_reg ,
    input [31:0] 					     desc_8_axuser_2_reg ,
    input [31:0] 					     desc_8_axuser_3_reg ,
    input [31:0] 					     desc_8_axuser_4_reg ,
    input [31:0] 					     desc_8_axuser_5_reg ,
    input [31:0] 					     desc_8_axuser_6_reg ,
    input [31:0] 					     desc_8_axuser_7_reg ,
    input [31:0] 					     desc_8_axuser_8_reg ,
    input [31:0] 					     desc_8_axuser_9_reg ,
    input [31:0] 					     desc_8_axuser_10_reg ,
    input [31:0] 					     desc_8_axuser_11_reg ,
    input [31:0] 					     desc_8_axuser_12_reg ,
    input [31:0] 					     desc_8_axuser_13_reg ,
    input [31:0] 					     desc_8_axuser_14_reg ,
    input [31:0] 					     desc_8_axuser_15_reg ,
    input [31:0] 					     desc_8_xuser_0_reg ,
    input [31:0] 					     desc_8_xuser_1_reg ,
    input [31:0] 					     desc_8_xuser_2_reg ,
    input [31:0] 					     desc_8_xuser_3_reg ,
    input [31:0] 					     desc_8_xuser_4_reg ,
    input [31:0] 					     desc_8_xuser_5_reg ,
    input [31:0] 					     desc_8_xuser_6_reg ,
    input [31:0] 					     desc_8_xuser_7_reg ,
    input [31:0] 					     desc_8_xuser_8_reg ,
    input [31:0] 					     desc_8_xuser_9_reg ,
    input [31:0] 					     desc_8_xuser_10_reg ,
    input [31:0] 					     desc_8_xuser_11_reg ,
    input [31:0] 					     desc_8_xuser_12_reg ,
    input [31:0] 					     desc_8_xuser_13_reg ,
    input [31:0] 					     desc_8_xuser_14_reg ,
    input [31:0] 					     desc_8_xuser_15_reg ,
    input [31:0] 					     desc_8_wuser_0_reg ,
    input [31:0] 					     desc_8_wuser_1_reg ,
    input [31:0] 					     desc_8_wuser_2_reg ,
    input [31:0] 					     desc_8_wuser_3_reg ,
    input [31:0] 					     desc_8_wuser_4_reg ,
    input [31:0] 					     desc_8_wuser_5_reg ,
    input [31:0] 					     desc_8_wuser_6_reg ,
    input [31:0] 					     desc_8_wuser_7_reg ,
    input [31:0] 					     desc_8_wuser_8_reg ,
    input [31:0] 					     desc_8_wuser_9_reg ,
    input [31:0] 					     desc_8_wuser_10_reg ,
    input [31:0] 					     desc_8_wuser_11_reg ,
    input [31:0] 					     desc_8_wuser_12_reg ,
    input [31:0] 					     desc_8_wuser_13_reg ,
    input [31:0] 					     desc_8_wuser_14_reg ,
    input [31:0] 					     desc_8_wuser_15_reg ,
    input [31:0] 					     desc_9_txn_type_reg ,
    input [31:0] 					     desc_9_size_reg ,
    input [31:0] 					     desc_9_data_offset_reg ,
    input [31:0] 					     desc_9_data_host_addr_0_reg ,
    input [31:0] 					     desc_9_data_host_addr_1_reg ,
    input [31:0] 					     desc_9_data_host_addr_2_reg ,
    input [31:0] 					     desc_9_data_host_addr_3_reg ,
    input [31:0] 					     desc_9_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_9_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_9_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_9_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_9_axsize_reg ,
    input [31:0] 					     desc_9_attr_reg ,
    input [31:0] 					     desc_9_axaddr_0_reg ,
    input [31:0] 					     desc_9_axaddr_1_reg ,
    input [31:0] 					     desc_9_axaddr_2_reg ,
    input [31:0] 					     desc_9_axaddr_3_reg ,
    input [31:0] 					     desc_9_axid_0_reg ,
    input [31:0] 					     desc_9_axid_1_reg ,
    input [31:0] 					     desc_9_axid_2_reg ,
    input [31:0] 					     desc_9_axid_3_reg ,
    input [31:0] 					     desc_9_axuser_0_reg ,
    input [31:0] 					     desc_9_axuser_1_reg ,
    input [31:0] 					     desc_9_axuser_2_reg ,
    input [31:0] 					     desc_9_axuser_3_reg ,
    input [31:0] 					     desc_9_axuser_4_reg ,
    input [31:0] 					     desc_9_axuser_5_reg ,
    input [31:0] 					     desc_9_axuser_6_reg ,
    input [31:0] 					     desc_9_axuser_7_reg ,
    input [31:0] 					     desc_9_axuser_8_reg ,
    input [31:0] 					     desc_9_axuser_9_reg ,
    input [31:0] 					     desc_9_axuser_10_reg ,
    input [31:0] 					     desc_9_axuser_11_reg ,
    input [31:0] 					     desc_9_axuser_12_reg ,
    input [31:0] 					     desc_9_axuser_13_reg ,
    input [31:0] 					     desc_9_axuser_14_reg ,
    input [31:0] 					     desc_9_axuser_15_reg ,
    input [31:0] 					     desc_9_xuser_0_reg ,
    input [31:0] 					     desc_9_xuser_1_reg ,
    input [31:0] 					     desc_9_xuser_2_reg ,
    input [31:0] 					     desc_9_xuser_3_reg ,
    input [31:0] 					     desc_9_xuser_4_reg ,
    input [31:0] 					     desc_9_xuser_5_reg ,
    input [31:0] 					     desc_9_xuser_6_reg ,
    input [31:0] 					     desc_9_xuser_7_reg ,
    input [31:0] 					     desc_9_xuser_8_reg ,
    input [31:0] 					     desc_9_xuser_9_reg ,
    input [31:0] 					     desc_9_xuser_10_reg ,
    input [31:0] 					     desc_9_xuser_11_reg ,
    input [31:0] 					     desc_9_xuser_12_reg ,
    input [31:0] 					     desc_9_xuser_13_reg ,
    input [31:0] 					     desc_9_xuser_14_reg ,
    input [31:0] 					     desc_9_xuser_15_reg ,
    input [31:0] 					     desc_9_wuser_0_reg ,
    input [31:0] 					     desc_9_wuser_1_reg ,
    input [31:0] 					     desc_9_wuser_2_reg ,
    input [31:0] 					     desc_9_wuser_3_reg ,
    input [31:0] 					     desc_9_wuser_4_reg ,
    input [31:0] 					     desc_9_wuser_5_reg ,
    input [31:0] 					     desc_9_wuser_6_reg ,
    input [31:0] 					     desc_9_wuser_7_reg ,
    input [31:0] 					     desc_9_wuser_8_reg ,
    input [31:0] 					     desc_9_wuser_9_reg ,
    input [31:0] 					     desc_9_wuser_10_reg ,
    input [31:0] 					     desc_9_wuser_11_reg ,
    input [31:0] 					     desc_9_wuser_12_reg ,
    input [31:0] 					     desc_9_wuser_13_reg ,
    input [31:0] 					     desc_9_wuser_14_reg ,
    input [31:0] 					     desc_9_wuser_15_reg ,
    input [31:0] 					     desc_10_txn_type_reg ,
    input [31:0] 					     desc_10_size_reg ,
    input [31:0] 					     desc_10_data_offset_reg ,
    input [31:0] 					     desc_10_data_host_addr_0_reg ,
    input [31:0] 					     desc_10_data_host_addr_1_reg ,
    input [31:0] 					     desc_10_data_host_addr_2_reg ,
    input [31:0] 					     desc_10_data_host_addr_3_reg ,
    input [31:0] 					     desc_10_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_10_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_10_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_10_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_10_axsize_reg ,
    input [31:0] 					     desc_10_attr_reg ,
    input [31:0] 					     desc_10_axaddr_0_reg ,
    input [31:0] 					     desc_10_axaddr_1_reg ,
    input [31:0] 					     desc_10_axaddr_2_reg ,
    input [31:0] 					     desc_10_axaddr_3_reg ,
    input [31:0] 					     desc_10_axid_0_reg ,
    input [31:0] 					     desc_10_axid_1_reg ,
    input [31:0] 					     desc_10_axid_2_reg ,
    input [31:0] 					     desc_10_axid_3_reg ,
    input [31:0] 					     desc_10_axuser_0_reg ,
    input [31:0] 					     desc_10_axuser_1_reg ,
    input [31:0] 					     desc_10_axuser_2_reg ,
    input [31:0] 					     desc_10_axuser_3_reg ,
    input [31:0] 					     desc_10_axuser_4_reg ,
    input [31:0] 					     desc_10_axuser_5_reg ,
    input [31:0] 					     desc_10_axuser_6_reg ,
    input [31:0] 					     desc_10_axuser_7_reg ,
    input [31:0] 					     desc_10_axuser_8_reg ,
    input [31:0] 					     desc_10_axuser_9_reg ,
    input [31:0] 					     desc_10_axuser_10_reg ,
    input [31:0] 					     desc_10_axuser_11_reg ,
    input [31:0] 					     desc_10_axuser_12_reg ,
    input [31:0] 					     desc_10_axuser_13_reg ,
    input [31:0] 					     desc_10_axuser_14_reg ,
    input [31:0] 					     desc_10_axuser_15_reg ,
    input [31:0] 					     desc_10_xuser_0_reg ,
    input [31:0] 					     desc_10_xuser_1_reg ,
    input [31:0] 					     desc_10_xuser_2_reg ,
    input [31:0] 					     desc_10_xuser_3_reg ,
    input [31:0] 					     desc_10_xuser_4_reg ,
    input [31:0] 					     desc_10_xuser_5_reg ,
    input [31:0] 					     desc_10_xuser_6_reg ,
    input [31:0] 					     desc_10_xuser_7_reg ,
    input [31:0] 					     desc_10_xuser_8_reg ,
    input [31:0] 					     desc_10_xuser_9_reg ,
    input [31:0] 					     desc_10_xuser_10_reg ,
    input [31:0] 					     desc_10_xuser_11_reg ,
    input [31:0] 					     desc_10_xuser_12_reg ,
    input [31:0] 					     desc_10_xuser_13_reg ,
    input [31:0] 					     desc_10_xuser_14_reg ,
    input [31:0] 					     desc_10_xuser_15_reg ,
    input [31:0] 					     desc_10_wuser_0_reg ,
    input [31:0] 					     desc_10_wuser_1_reg ,
    input [31:0] 					     desc_10_wuser_2_reg ,
    input [31:0] 					     desc_10_wuser_3_reg ,
    input [31:0] 					     desc_10_wuser_4_reg ,
    input [31:0] 					     desc_10_wuser_5_reg ,
    input [31:0] 					     desc_10_wuser_6_reg ,
    input [31:0] 					     desc_10_wuser_7_reg ,
    input [31:0] 					     desc_10_wuser_8_reg ,
    input [31:0] 					     desc_10_wuser_9_reg ,
    input [31:0] 					     desc_10_wuser_10_reg ,
    input [31:0] 					     desc_10_wuser_11_reg ,
    input [31:0] 					     desc_10_wuser_12_reg ,
    input [31:0] 					     desc_10_wuser_13_reg ,
    input [31:0] 					     desc_10_wuser_14_reg ,
    input [31:0] 					     desc_10_wuser_15_reg ,
    input [31:0] 					     desc_11_txn_type_reg ,
    input [31:0] 					     desc_11_size_reg ,
    input [31:0] 					     desc_11_data_offset_reg ,
    input [31:0] 					     desc_11_data_host_addr_0_reg ,
    input [31:0] 					     desc_11_data_host_addr_1_reg ,
    input [31:0] 					     desc_11_data_host_addr_2_reg ,
    input [31:0] 					     desc_11_data_host_addr_3_reg ,
    input [31:0] 					     desc_11_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_11_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_11_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_11_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_11_axsize_reg ,
    input [31:0] 					     desc_11_attr_reg ,
    input [31:0] 					     desc_11_axaddr_0_reg ,
    input [31:0] 					     desc_11_axaddr_1_reg ,
    input [31:0] 					     desc_11_axaddr_2_reg ,
    input [31:0] 					     desc_11_axaddr_3_reg ,
    input [31:0] 					     desc_11_axid_0_reg ,
    input [31:0] 					     desc_11_axid_1_reg ,
    input [31:0] 					     desc_11_axid_2_reg ,
    input [31:0] 					     desc_11_axid_3_reg ,
    input [31:0] 					     desc_11_axuser_0_reg ,
    input [31:0] 					     desc_11_axuser_1_reg ,
    input [31:0] 					     desc_11_axuser_2_reg ,
    input [31:0] 					     desc_11_axuser_3_reg ,
    input [31:0] 					     desc_11_axuser_4_reg ,
    input [31:0] 					     desc_11_axuser_5_reg ,
    input [31:0] 					     desc_11_axuser_6_reg ,
    input [31:0] 					     desc_11_axuser_7_reg ,
    input [31:0] 					     desc_11_axuser_8_reg ,
    input [31:0] 					     desc_11_axuser_9_reg ,
    input [31:0] 					     desc_11_axuser_10_reg ,
    input [31:0] 					     desc_11_axuser_11_reg ,
    input [31:0] 					     desc_11_axuser_12_reg ,
    input [31:0] 					     desc_11_axuser_13_reg ,
    input [31:0] 					     desc_11_axuser_14_reg ,
    input [31:0] 					     desc_11_axuser_15_reg ,
    input [31:0] 					     desc_11_xuser_0_reg ,
    input [31:0] 					     desc_11_xuser_1_reg ,
    input [31:0] 					     desc_11_xuser_2_reg ,
    input [31:0] 					     desc_11_xuser_3_reg ,
    input [31:0] 					     desc_11_xuser_4_reg ,
    input [31:0] 					     desc_11_xuser_5_reg ,
    input [31:0] 					     desc_11_xuser_6_reg ,
    input [31:0] 					     desc_11_xuser_7_reg ,
    input [31:0] 					     desc_11_xuser_8_reg ,
    input [31:0] 					     desc_11_xuser_9_reg ,
    input [31:0] 					     desc_11_xuser_10_reg ,
    input [31:0] 					     desc_11_xuser_11_reg ,
    input [31:0] 					     desc_11_xuser_12_reg ,
    input [31:0] 					     desc_11_xuser_13_reg ,
    input [31:0] 					     desc_11_xuser_14_reg ,
    input [31:0] 					     desc_11_xuser_15_reg ,
    input [31:0] 					     desc_11_wuser_0_reg ,
    input [31:0] 					     desc_11_wuser_1_reg ,
    input [31:0] 					     desc_11_wuser_2_reg ,
    input [31:0] 					     desc_11_wuser_3_reg ,
    input [31:0] 					     desc_11_wuser_4_reg ,
    input [31:0] 					     desc_11_wuser_5_reg ,
    input [31:0] 					     desc_11_wuser_6_reg ,
    input [31:0] 					     desc_11_wuser_7_reg ,
    input [31:0] 					     desc_11_wuser_8_reg ,
    input [31:0] 					     desc_11_wuser_9_reg ,
    input [31:0] 					     desc_11_wuser_10_reg ,
    input [31:0] 					     desc_11_wuser_11_reg ,
    input [31:0] 					     desc_11_wuser_12_reg ,
    input [31:0] 					     desc_11_wuser_13_reg ,
    input [31:0] 					     desc_11_wuser_14_reg ,
    input [31:0] 					     desc_11_wuser_15_reg ,
    input [31:0] 					     desc_12_txn_type_reg ,
    input [31:0] 					     desc_12_size_reg ,
    input [31:0] 					     desc_12_data_offset_reg ,
    input [31:0] 					     desc_12_data_host_addr_0_reg ,
    input [31:0] 					     desc_12_data_host_addr_1_reg ,
    input [31:0] 					     desc_12_data_host_addr_2_reg ,
    input [31:0] 					     desc_12_data_host_addr_3_reg ,
    input [31:0] 					     desc_12_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_12_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_12_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_12_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_12_axsize_reg ,
    input [31:0] 					     desc_12_attr_reg ,
    input [31:0] 					     desc_12_axaddr_0_reg ,
    input [31:0] 					     desc_12_axaddr_1_reg ,
    input [31:0] 					     desc_12_axaddr_2_reg ,
    input [31:0] 					     desc_12_axaddr_3_reg ,
    input [31:0] 					     desc_12_axid_0_reg ,
    input [31:0] 					     desc_12_axid_1_reg ,
    input [31:0] 					     desc_12_axid_2_reg ,
    input [31:0] 					     desc_12_axid_3_reg ,
    input [31:0] 					     desc_12_axuser_0_reg ,
    input [31:0] 					     desc_12_axuser_1_reg ,
    input [31:0] 					     desc_12_axuser_2_reg ,
    input [31:0] 					     desc_12_axuser_3_reg ,
    input [31:0] 					     desc_12_axuser_4_reg ,
    input [31:0] 					     desc_12_axuser_5_reg ,
    input [31:0] 					     desc_12_axuser_6_reg ,
    input [31:0] 					     desc_12_axuser_7_reg ,
    input [31:0] 					     desc_12_axuser_8_reg ,
    input [31:0] 					     desc_12_axuser_9_reg ,
    input [31:0] 					     desc_12_axuser_10_reg ,
    input [31:0] 					     desc_12_axuser_11_reg ,
    input [31:0] 					     desc_12_axuser_12_reg ,
    input [31:0] 					     desc_12_axuser_13_reg ,
    input [31:0] 					     desc_12_axuser_14_reg ,
    input [31:0] 					     desc_12_axuser_15_reg ,
    input [31:0] 					     desc_12_xuser_0_reg ,
    input [31:0] 					     desc_12_xuser_1_reg ,
    input [31:0] 					     desc_12_xuser_2_reg ,
    input [31:0] 					     desc_12_xuser_3_reg ,
    input [31:0] 					     desc_12_xuser_4_reg ,
    input [31:0] 					     desc_12_xuser_5_reg ,
    input [31:0] 					     desc_12_xuser_6_reg ,
    input [31:0] 					     desc_12_xuser_7_reg ,
    input [31:0] 					     desc_12_xuser_8_reg ,
    input [31:0] 					     desc_12_xuser_9_reg ,
    input [31:0] 					     desc_12_xuser_10_reg ,
    input [31:0] 					     desc_12_xuser_11_reg ,
    input [31:0] 					     desc_12_xuser_12_reg ,
    input [31:0] 					     desc_12_xuser_13_reg ,
    input [31:0] 					     desc_12_xuser_14_reg ,
    input [31:0] 					     desc_12_xuser_15_reg ,
    input [31:0] 					     desc_12_wuser_0_reg ,
    input [31:0] 					     desc_12_wuser_1_reg ,
    input [31:0] 					     desc_12_wuser_2_reg ,
    input [31:0] 					     desc_12_wuser_3_reg ,
    input [31:0] 					     desc_12_wuser_4_reg ,
    input [31:0] 					     desc_12_wuser_5_reg ,
    input [31:0] 					     desc_12_wuser_6_reg ,
    input [31:0] 					     desc_12_wuser_7_reg ,
    input [31:0] 					     desc_12_wuser_8_reg ,
    input [31:0] 					     desc_12_wuser_9_reg ,
    input [31:0] 					     desc_12_wuser_10_reg ,
    input [31:0] 					     desc_12_wuser_11_reg ,
    input [31:0] 					     desc_12_wuser_12_reg ,
    input [31:0] 					     desc_12_wuser_13_reg ,
    input [31:0] 					     desc_12_wuser_14_reg ,
    input [31:0] 					     desc_12_wuser_15_reg ,
    input [31:0] 					     desc_13_txn_type_reg ,
    input [31:0] 					     desc_13_size_reg ,
    input [31:0] 					     desc_13_data_offset_reg ,
    input [31:0] 					     desc_13_data_host_addr_0_reg ,
    input [31:0] 					     desc_13_data_host_addr_1_reg ,
    input [31:0] 					     desc_13_data_host_addr_2_reg ,
    input [31:0] 					     desc_13_data_host_addr_3_reg ,
    input [31:0] 					     desc_13_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_13_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_13_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_13_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_13_axsize_reg ,
    input [31:0] 					     desc_13_attr_reg ,
    input [31:0] 					     desc_13_axaddr_0_reg ,
    input [31:0] 					     desc_13_axaddr_1_reg ,
    input [31:0] 					     desc_13_axaddr_2_reg ,
    input [31:0] 					     desc_13_axaddr_3_reg ,
    input [31:0] 					     desc_13_axid_0_reg ,
    input [31:0] 					     desc_13_axid_1_reg ,
    input [31:0] 					     desc_13_axid_2_reg ,
    input [31:0] 					     desc_13_axid_3_reg ,
    input [31:0] 					     desc_13_axuser_0_reg ,
    input [31:0] 					     desc_13_axuser_1_reg ,
    input [31:0] 					     desc_13_axuser_2_reg ,
    input [31:0] 					     desc_13_axuser_3_reg ,
    input [31:0] 					     desc_13_axuser_4_reg ,
    input [31:0] 					     desc_13_axuser_5_reg ,
    input [31:0] 					     desc_13_axuser_6_reg ,
    input [31:0] 					     desc_13_axuser_7_reg ,
    input [31:0] 					     desc_13_axuser_8_reg ,
    input [31:0] 					     desc_13_axuser_9_reg ,
    input [31:0] 					     desc_13_axuser_10_reg ,
    input [31:0] 					     desc_13_axuser_11_reg ,
    input [31:0] 					     desc_13_axuser_12_reg ,
    input [31:0] 					     desc_13_axuser_13_reg ,
    input [31:0] 					     desc_13_axuser_14_reg ,
    input [31:0] 					     desc_13_axuser_15_reg ,
    input [31:0] 					     desc_13_xuser_0_reg ,
    input [31:0] 					     desc_13_xuser_1_reg ,
    input [31:0] 					     desc_13_xuser_2_reg ,
    input [31:0] 					     desc_13_xuser_3_reg ,
    input [31:0] 					     desc_13_xuser_4_reg ,
    input [31:0] 					     desc_13_xuser_5_reg ,
    input [31:0] 					     desc_13_xuser_6_reg ,
    input [31:0] 					     desc_13_xuser_7_reg ,
    input [31:0] 					     desc_13_xuser_8_reg ,
    input [31:0] 					     desc_13_xuser_9_reg ,
    input [31:0] 					     desc_13_xuser_10_reg ,
    input [31:0] 					     desc_13_xuser_11_reg ,
    input [31:0] 					     desc_13_xuser_12_reg ,
    input [31:0] 					     desc_13_xuser_13_reg ,
    input [31:0] 					     desc_13_xuser_14_reg ,
    input [31:0] 					     desc_13_xuser_15_reg ,
    input [31:0] 					     desc_13_wuser_0_reg ,
    input [31:0] 					     desc_13_wuser_1_reg ,
    input [31:0] 					     desc_13_wuser_2_reg ,
    input [31:0] 					     desc_13_wuser_3_reg ,
    input [31:0] 					     desc_13_wuser_4_reg ,
    input [31:0] 					     desc_13_wuser_5_reg ,
    input [31:0] 					     desc_13_wuser_6_reg ,
    input [31:0] 					     desc_13_wuser_7_reg ,
    input [31:0] 					     desc_13_wuser_8_reg ,
    input [31:0] 					     desc_13_wuser_9_reg ,
    input [31:0] 					     desc_13_wuser_10_reg ,
    input [31:0] 					     desc_13_wuser_11_reg ,
    input [31:0] 					     desc_13_wuser_12_reg ,
    input [31:0] 					     desc_13_wuser_13_reg ,
    input [31:0] 					     desc_13_wuser_14_reg ,
    input [31:0] 					     desc_13_wuser_15_reg ,
    input [31:0] 					     desc_14_txn_type_reg ,
    input [31:0] 					     desc_14_size_reg ,
    input [31:0] 					     desc_14_data_offset_reg ,
    input [31:0] 					     desc_14_data_host_addr_0_reg ,
    input [31:0] 					     desc_14_data_host_addr_1_reg ,
    input [31:0] 					     desc_14_data_host_addr_2_reg ,
    input [31:0] 					     desc_14_data_host_addr_3_reg ,
    input [31:0] 					     desc_14_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_14_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_14_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_14_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_14_axsize_reg ,
    input [31:0] 					     desc_14_attr_reg ,
    input [31:0] 					     desc_14_axaddr_0_reg ,
    input [31:0] 					     desc_14_axaddr_1_reg ,
    input [31:0] 					     desc_14_axaddr_2_reg ,
    input [31:0] 					     desc_14_axaddr_3_reg ,
    input [31:0] 					     desc_14_axid_0_reg ,
    input [31:0] 					     desc_14_axid_1_reg ,
    input [31:0] 					     desc_14_axid_2_reg ,
    input [31:0] 					     desc_14_axid_3_reg ,
    input [31:0] 					     desc_14_axuser_0_reg ,
    input [31:0] 					     desc_14_axuser_1_reg ,
    input [31:0] 					     desc_14_axuser_2_reg ,
    input [31:0] 					     desc_14_axuser_3_reg ,
    input [31:0] 					     desc_14_axuser_4_reg ,
    input [31:0] 					     desc_14_axuser_5_reg ,
    input [31:0] 					     desc_14_axuser_6_reg ,
    input [31:0] 					     desc_14_axuser_7_reg ,
    input [31:0] 					     desc_14_axuser_8_reg ,
    input [31:0] 					     desc_14_axuser_9_reg ,
    input [31:0] 					     desc_14_axuser_10_reg ,
    input [31:0] 					     desc_14_axuser_11_reg ,
    input [31:0] 					     desc_14_axuser_12_reg ,
    input [31:0] 					     desc_14_axuser_13_reg ,
    input [31:0] 					     desc_14_axuser_14_reg ,
    input [31:0] 					     desc_14_axuser_15_reg ,
    input [31:0] 					     desc_14_xuser_0_reg ,
    input [31:0] 					     desc_14_xuser_1_reg ,
    input [31:0] 					     desc_14_xuser_2_reg ,
    input [31:0] 					     desc_14_xuser_3_reg ,
    input [31:0] 					     desc_14_xuser_4_reg ,
    input [31:0] 					     desc_14_xuser_5_reg ,
    input [31:0] 					     desc_14_xuser_6_reg ,
    input [31:0] 					     desc_14_xuser_7_reg ,
    input [31:0] 					     desc_14_xuser_8_reg ,
    input [31:0] 					     desc_14_xuser_9_reg ,
    input [31:0] 					     desc_14_xuser_10_reg ,
    input [31:0] 					     desc_14_xuser_11_reg ,
    input [31:0] 					     desc_14_xuser_12_reg ,
    input [31:0] 					     desc_14_xuser_13_reg ,
    input [31:0] 					     desc_14_xuser_14_reg ,
    input [31:0] 					     desc_14_xuser_15_reg ,
    input [31:0] 					     desc_14_wuser_0_reg ,
    input [31:0] 					     desc_14_wuser_1_reg ,
    input [31:0] 					     desc_14_wuser_2_reg ,
    input [31:0] 					     desc_14_wuser_3_reg ,
    input [31:0] 					     desc_14_wuser_4_reg ,
    input [31:0] 					     desc_14_wuser_5_reg ,
    input [31:0] 					     desc_14_wuser_6_reg ,
    input [31:0] 					     desc_14_wuser_7_reg ,
    input [31:0] 					     desc_14_wuser_8_reg ,
    input [31:0] 					     desc_14_wuser_9_reg ,
    input [31:0] 					     desc_14_wuser_10_reg ,
    input [31:0] 					     desc_14_wuser_11_reg ,
    input [31:0] 					     desc_14_wuser_12_reg ,
    input [31:0] 					     desc_14_wuser_13_reg ,
    input [31:0] 					     desc_14_wuser_14_reg ,
    input [31:0] 					     desc_14_wuser_15_reg ,
    input [31:0] 					     desc_15_txn_type_reg ,
    input [31:0] 					     desc_15_size_reg ,
    input [31:0] 					     desc_15_data_offset_reg ,
    input [31:0] 					     desc_15_data_host_addr_0_reg ,
    input [31:0] 					     desc_15_data_host_addr_1_reg ,
    input [31:0] 					     desc_15_data_host_addr_2_reg ,
    input [31:0] 					     desc_15_data_host_addr_3_reg ,
    input [31:0] 					     desc_15_wstrb_host_addr_0_reg ,
    input [31:0] 					     desc_15_wstrb_host_addr_1_reg ,
    input [31:0] 					     desc_15_wstrb_host_addr_2_reg ,
    input [31:0] 					     desc_15_wstrb_host_addr_3_reg ,
    input [31:0] 					     desc_15_axsize_reg ,
    input [31:0] 					     desc_15_attr_reg ,
    input [31:0] 					     desc_15_axaddr_0_reg ,
    input [31:0] 					     desc_15_axaddr_1_reg ,
    input [31:0] 					     desc_15_axaddr_2_reg ,
    input [31:0] 					     desc_15_axaddr_3_reg ,
    input [31:0] 					     desc_15_axid_0_reg ,
    input [31:0] 					     desc_15_axid_1_reg ,
    input [31:0] 					     desc_15_axid_2_reg ,
    input [31:0] 					     desc_15_axid_3_reg ,
    input [31:0] 					     desc_15_axuser_0_reg ,
    input [31:0] 					     desc_15_axuser_1_reg ,
    input [31:0] 					     desc_15_axuser_2_reg ,
    input [31:0] 					     desc_15_axuser_3_reg ,
    input [31:0] 					     desc_15_axuser_4_reg ,
    input [31:0] 					     desc_15_axuser_5_reg ,
    input [31:0] 					     desc_15_axuser_6_reg ,
    input [31:0] 					     desc_15_axuser_7_reg ,
    input [31:0] 					     desc_15_axuser_8_reg ,
    input [31:0] 					     desc_15_axuser_9_reg ,
    input [31:0] 					     desc_15_axuser_10_reg ,
    input [31:0] 					     desc_15_axuser_11_reg ,
    input [31:0] 					     desc_15_axuser_12_reg ,
    input [31:0] 					     desc_15_axuser_13_reg ,
    input [31:0] 					     desc_15_axuser_14_reg ,
    input [31:0] 					     desc_15_axuser_15_reg ,
    input [31:0] 					     desc_15_xuser_0_reg ,
    input [31:0] 					     desc_15_xuser_1_reg ,
    input [31:0] 					     desc_15_xuser_2_reg ,
    input [31:0] 					     desc_15_xuser_3_reg ,
    input [31:0] 					     desc_15_xuser_4_reg ,
    input [31:0] 					     desc_15_xuser_5_reg ,
    input [31:0] 					     desc_15_xuser_6_reg ,
    input [31:0] 					     desc_15_xuser_7_reg ,
    input [31:0] 					     desc_15_xuser_8_reg ,
    input [31:0] 					     desc_15_xuser_9_reg ,
    input [31:0] 					     desc_15_xuser_10_reg ,
    input [31:0] 					     desc_15_xuser_11_reg ,
    input [31:0] 					     desc_15_xuser_12_reg ,
    input [31:0] 					     desc_15_xuser_13_reg ,
    input [31:0] 					     desc_15_xuser_14_reg ,
    input [31:0] 					     desc_15_xuser_15_reg ,
    input [31:0] 					     desc_15_wuser_0_reg ,
    input [31:0] 					     desc_15_wuser_1_reg ,
    input [31:0] 					     desc_15_wuser_2_reg ,
    input [31:0] 					     desc_15_wuser_3_reg ,
    input [31:0] 					     desc_15_wuser_4_reg ,
    input [31:0] 					     desc_15_wuser_5_reg ,
    input [31:0] 					     desc_15_wuser_6_reg ,
    input [31:0] 					     desc_15_wuser_7_reg ,
    input [31:0] 					     desc_15_wuser_8_reg ,
    input [31:0] 					     desc_15_wuser_9_reg ,
    input [31:0] 					     desc_15_wuser_10_reg ,
    input [31:0] 					     desc_15_wuser_11_reg ,
    input [31:0] 					     desc_15_wuser_12_reg ,
    input [31:0] 					     desc_15_wuser_13_reg ,
    input [31:0] 					     desc_15_wuser_14_reg ,
    input [31:0] 					     desc_15_wuser_15_reg ,
  
    output [31:0] 					     uc2rb_intr_error_status_reg ,
    output [31:0] 					     uc2rb_ownership_reg ,
    output [31:0] 					     uc2rb_intr_comp_status_reg ,
    output [31:0] 					     uc2rb_status_resp_reg ,
    output [31:0] 					     uc2rb_status_busy_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_0_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_1_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_2_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_3_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_4_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_5_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_6_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_7_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_8_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_9_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_10_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_11_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_12_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_13_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_14_xuser_15_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_0_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_1_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_2_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_3_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_4_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_5_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_6_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_7_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_8_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_9_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_10_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_11_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_12_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_13_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_14_reg ,
    output [31:0] 					     uc2rb_desc_15_xuser_15_reg ,

    output [31:0] 					     uc2rb_intr_error_status_reg_we ,
    output [31:0] 					     uc2rb_ownership_reg_we ,
    output [31:0] 					     uc2rb_intr_comp_status_reg_we ,
    output [31:0] 					     uc2rb_status_resp_reg_we ,
    output [31:0] 					     uc2rb_status_busy_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_0_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_1_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_2_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_3_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_4_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_5_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_6_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_7_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_8_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_9_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_10_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_11_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_12_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_13_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_14_xuser_15_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_0_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_1_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_2_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_3_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_4_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_5_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_6_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_7_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_8_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_9_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_10_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_11_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_12_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_13_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_14_reg_we ,
    output [31:0] 					     uc2rb_desc_15_xuser_15_reg_we ,


    //M_AXI_USR
//`ifdef USER_AXI4        
    output [M_AXI_USR_ID_WIDTH-1:0] 			     m_axi_usr_awid, 
    output [M_AXI_USR_ADDR_WIDTH-1:0] 			     m_axi_usr_awaddr, 
    output [7:0] 					     m_axi_usr_awlen, 
    output [2:0] 					     m_axi_usr_awsize, 
    output [1:0] 					     m_axi_usr_awburst, 
    output [1:0] 					     m_axi_usr_awlock, 
    output [3:0] 					     m_axi_usr_awcache, 
    output [2:0] 					     m_axi_usr_awprot, 
    output [3:0] 					     m_axi_usr_awqos, 
    output [3:0] 					     m_axi_usr_awregion, 
    output [M_AXI_USR_AWUSER_WIDTH-1:0] 		     m_axi_usr_awuser, 
    output 						     m_axi_usr_awvalid, 
    input 						     m_axi_usr_awready, 
    output [M_AXI_USR_DATA_WIDTH-1:0] 			     m_axi_usr_wdata, 
    output [(M_AXI_USR_DATA_WIDTH/8)-1:0] 		     m_axi_usr_wstrb,
    output 						     m_axi_usr_wlast, 
    output [M_AXI_USR_WUSER_WIDTH-1:0] 			     m_axi_usr_wuser, 
    output 						     m_axi_usr_wvalid, 
    input 						     m_axi_usr_wready, 
    input [M_AXI_USR_ID_WIDTH-1:0] 			     m_axi_usr_bid, 
    input [1:0] 					     m_axi_usr_bresp, 
    input [M_AXI_USR_BUSER_WIDTH-1:0] 			     m_axi_usr_buser, 
    input 						     m_axi_usr_bvalid, 
    output 						     m_axi_usr_bready, 
    output [M_AXI_USR_ID_WIDTH-1:0] 			     m_axi_usr_arid, 
    output [M_AXI_USR_ADDR_WIDTH-1:0] 			     m_axi_usr_araddr, 
    output [7:0] 					     m_axi_usr_arlen, 
    output [2:0] 					     m_axi_usr_arsize, 
    output [1:0] 					     m_axi_usr_arburst, 
    output [1:0] 					     m_axi_usr_arlock, 
    output [3:0] 					     m_axi_usr_arcache, 
    output [2:0] 					     m_axi_usr_arprot, 
    output [3:0] 					     m_axi_usr_arqos, 
    output [3:0] 					     m_axi_usr_arregion, 
    output [M_AXI_USR_ARUSER_WIDTH-1:0] 		     m_axi_usr_aruser, 
    output 						     m_axi_usr_arvalid, 
    input 						     m_axi_usr_arready, 
    input [M_AXI_USR_ID_WIDTH-1:0] 			     m_axi_usr_rid, 
    input [M_AXI_USR_DATA_WIDTH-1:0] 			     m_axi_usr_rdata, 
    input [1:0] 					     m_axi_usr_rresp, 
    input 						     m_axi_usr_rlast, 
    input [M_AXI_USR_RUSER_WIDTH-1:0] 			     m_axi_usr_ruser, 
    input 						     m_axi_usr_rvalid, 
    output 						     m_axi_usr_rready, 

	
    output [M_AXI_USR_ID_WIDTH-1:0] 			     m_axi_usr_wid

    /*AUTOARG*/);

   wire [(`CLOG2(MAX_DESC))-1:0] 			     uc2rb_wr_desc_id;

   

   localparam M_AXI_USR_LEN_WIDTH = (EN_INTFM_AXI4==1) ? 8 : 4;
   
   
   axi_master_control  #(/*AutoInstParam*/
			 // Parameters
			 .M_AXI_USR_ADDR_WIDTH	(M_AXI_USR_ADDR_WIDTH),
			 .M_AXI_USR_DATA_WIDTH	(M_AXI_USR_DATA_WIDTH),
			 .M_AXI_USR_ID_WIDTH	(M_AXI_USR_ID_WIDTH),
			 .M_AXI_USR_AWUSER_WIDTH (M_AXI_USR_AWUSER_WIDTH),
			 .M_AXI_USR_ARUSER_WIDTH (M_AXI_USR_ARUSER_WIDTH),
			 .M_AXI_USR_WUSER_WIDTH  (M_AXI_USR_WUSER_WIDTH),
			 .M_AXI_USR_RUSER_WIDTH  (M_AXI_USR_RUSER_WIDTH),
			 .M_AXI_USR_BUSER_WIDTH  (M_AXI_USR_BUSER_WIDTH),
			 .M_AXI_USR_LEN_WIDTH	(M_AXI_USR_LEN_WIDTH),
			 .RAM_SIZE				(RAM_SIZE),
			 .MAX_DESC				(MAX_DESC),
			 .RTL_USE_MODE			(0), //Used as User Master 
			 .UC_AXI_DATA_WIDTH		(M_AXI_USR_DATA_WIDTH),
			 .EN_INTFM_AXI4 (EN_INTFM_AXI4),
			 .EN_INTFM_AXI3 (EN_INTFM_AXI3),
			 .EN_INTFM_AXI4LITE (EN_INTFM_AXI4LITE))
   
   axi_master_inst 
     ( /*AUTOINST*/
       // Outputs
       .uc2rb_rd_addr					(uc2rb_rd_addr[(`CLOG2(RAM_SIZE/(M_AXI_USR_DATA_WIDTH/8)))-1:0] ),
       .uc2rb_wr_we						(uc2rb_wr_we),
       .uc2rb_wr_bwe						(uc2rb_wr_bwe[(M_AXI_USR_DATA_WIDTH/8-1):0]),
       .uc2rb_wr_addr					(uc2rb_wr_addr[(`CLOG2(RAM_SIZE/(M_AXI_USR_DATA_WIDTH/8)))-1:0]),
       .uc2rb_wr_data					(uc2rb_wr_data[M_AXI_USR_DATA_WIDTH-1:0]),
       .uc2rb_wr_desc_id					(uc2rb_wr_desc_id[(`CLOG2(MAX_DESC))-1:0]),
       .uc2hm_trig						(uc2hm_trig[15:0]),
       .uc2rb_intr_error_status_reg		(uc2rb_intr_error_status_reg[31:0]),
       .uc2rb_ownership_reg				(uc2rb_ownership_reg[31:0]),
       .uc2rb_intr_comp_status_reg		(uc2rb_intr_comp_status_reg[31:0]),
       .uc2rb_status_resp_reg			(uc2rb_status_resp_reg[31:0]),
       .uc2rb_status_busy_reg			(uc2rb_status_busy_reg[31:0]),
       .uc2rb_desc_0_xuser_0_reg			(uc2rb_desc_0_xuser_0_reg[31:0]),
       .uc2rb_desc_0_xuser_1_reg			(uc2rb_desc_0_xuser_1_reg[31:0]),
       .uc2rb_desc_0_xuser_2_reg			(uc2rb_desc_0_xuser_2_reg[31:0]),
       .uc2rb_desc_0_xuser_3_reg			(uc2rb_desc_0_xuser_3_reg[31:0]),
       .uc2rb_desc_0_xuser_4_reg			(uc2rb_desc_0_xuser_4_reg[31:0]),
       .uc2rb_desc_0_xuser_5_reg			(uc2rb_desc_0_xuser_5_reg[31:0]),
       .uc2rb_desc_0_xuser_6_reg			(uc2rb_desc_0_xuser_6_reg[31:0]),
       .uc2rb_desc_0_xuser_7_reg			(uc2rb_desc_0_xuser_7_reg[31:0]),
       .uc2rb_desc_0_xuser_8_reg			(uc2rb_desc_0_xuser_8_reg[31:0]),
       .uc2rb_desc_0_xuser_9_reg			(uc2rb_desc_0_xuser_9_reg[31:0]),
       .uc2rb_desc_0_xuser_10_reg		(uc2rb_desc_0_xuser_10_reg[31:0]),
       .uc2rb_desc_0_xuser_11_reg		(uc2rb_desc_0_xuser_11_reg[31:0]),
       .uc2rb_desc_0_xuser_12_reg		(uc2rb_desc_0_xuser_12_reg[31:0]),
       .uc2rb_desc_0_xuser_13_reg		(uc2rb_desc_0_xuser_13_reg[31:0]),
       .uc2rb_desc_0_xuser_14_reg		(uc2rb_desc_0_xuser_14_reg[31:0]),
       .uc2rb_desc_0_xuser_15_reg		(uc2rb_desc_0_xuser_15_reg[31:0]),
       .uc2rb_desc_1_xuser_0_reg			(uc2rb_desc_1_xuser_0_reg[31:0]),
       .uc2rb_desc_1_xuser_1_reg			(uc2rb_desc_1_xuser_1_reg[31:0]),
       .uc2rb_desc_1_xuser_2_reg			(uc2rb_desc_1_xuser_2_reg[31:0]),
       .uc2rb_desc_1_xuser_3_reg			(uc2rb_desc_1_xuser_3_reg[31:0]),
       .uc2rb_desc_1_xuser_4_reg			(uc2rb_desc_1_xuser_4_reg[31:0]),
       .uc2rb_desc_1_xuser_5_reg			(uc2rb_desc_1_xuser_5_reg[31:0]),
       .uc2rb_desc_1_xuser_6_reg			(uc2rb_desc_1_xuser_6_reg[31:0]),
       .uc2rb_desc_1_xuser_7_reg			(uc2rb_desc_1_xuser_7_reg[31:0]),
       .uc2rb_desc_1_xuser_8_reg			(uc2rb_desc_1_xuser_8_reg[31:0]),
       .uc2rb_desc_1_xuser_9_reg			(uc2rb_desc_1_xuser_9_reg[31:0]),
       .uc2rb_desc_1_xuser_10_reg		(uc2rb_desc_1_xuser_10_reg[31:0]),
       .uc2rb_desc_1_xuser_11_reg		(uc2rb_desc_1_xuser_11_reg[31:0]),
       .uc2rb_desc_1_xuser_12_reg		(uc2rb_desc_1_xuser_12_reg[31:0]),
       .uc2rb_desc_1_xuser_13_reg		(uc2rb_desc_1_xuser_13_reg[31:0]),
       .uc2rb_desc_1_xuser_14_reg		(uc2rb_desc_1_xuser_14_reg[31:0]),
       .uc2rb_desc_1_xuser_15_reg		(uc2rb_desc_1_xuser_15_reg[31:0]),
       .uc2rb_desc_2_xuser_0_reg			(uc2rb_desc_2_xuser_0_reg[31:0]),
       .uc2rb_desc_2_xuser_1_reg			(uc2rb_desc_2_xuser_1_reg[31:0]),
       .uc2rb_desc_2_xuser_2_reg			(uc2rb_desc_2_xuser_2_reg[31:0]),
       .uc2rb_desc_2_xuser_3_reg			(uc2rb_desc_2_xuser_3_reg[31:0]),
       .uc2rb_desc_2_xuser_4_reg			(uc2rb_desc_2_xuser_4_reg[31:0]),
       .uc2rb_desc_2_xuser_5_reg			(uc2rb_desc_2_xuser_5_reg[31:0]),
       .uc2rb_desc_2_xuser_6_reg			(uc2rb_desc_2_xuser_6_reg[31:0]),
       .uc2rb_desc_2_xuser_7_reg			(uc2rb_desc_2_xuser_7_reg[31:0]),
       .uc2rb_desc_2_xuser_8_reg			(uc2rb_desc_2_xuser_8_reg[31:0]),
       .uc2rb_desc_2_xuser_9_reg			(uc2rb_desc_2_xuser_9_reg[31:0]),
       .uc2rb_desc_2_xuser_10_reg		(uc2rb_desc_2_xuser_10_reg[31:0]),
       .uc2rb_desc_2_xuser_11_reg		(uc2rb_desc_2_xuser_11_reg[31:0]),
       .uc2rb_desc_2_xuser_12_reg		(uc2rb_desc_2_xuser_12_reg[31:0]),
       .uc2rb_desc_2_xuser_13_reg		(uc2rb_desc_2_xuser_13_reg[31:0]),
       .uc2rb_desc_2_xuser_14_reg		(uc2rb_desc_2_xuser_14_reg[31:0]),
       .uc2rb_desc_2_xuser_15_reg		(uc2rb_desc_2_xuser_15_reg[31:0]),
       .uc2rb_desc_3_xuser_0_reg			(uc2rb_desc_3_xuser_0_reg[31:0]),
       .uc2rb_desc_3_xuser_1_reg			(uc2rb_desc_3_xuser_1_reg[31:0]),
       .uc2rb_desc_3_xuser_2_reg			(uc2rb_desc_3_xuser_2_reg[31:0]),
       .uc2rb_desc_3_xuser_3_reg			(uc2rb_desc_3_xuser_3_reg[31:0]),
       .uc2rb_desc_3_xuser_4_reg			(uc2rb_desc_3_xuser_4_reg[31:0]),
       .uc2rb_desc_3_xuser_5_reg			(uc2rb_desc_3_xuser_5_reg[31:0]),
       .uc2rb_desc_3_xuser_6_reg			(uc2rb_desc_3_xuser_6_reg[31:0]),
       .uc2rb_desc_3_xuser_7_reg			(uc2rb_desc_3_xuser_7_reg[31:0]),
       .uc2rb_desc_3_xuser_8_reg			(uc2rb_desc_3_xuser_8_reg[31:0]),
       .uc2rb_desc_3_xuser_9_reg			(uc2rb_desc_3_xuser_9_reg[31:0]),
       .uc2rb_desc_3_xuser_10_reg		(uc2rb_desc_3_xuser_10_reg[31:0]),
       .uc2rb_desc_3_xuser_11_reg		(uc2rb_desc_3_xuser_11_reg[31:0]),
       .uc2rb_desc_3_xuser_12_reg		(uc2rb_desc_3_xuser_12_reg[31:0]),
       .uc2rb_desc_3_xuser_13_reg		(uc2rb_desc_3_xuser_13_reg[31:0]),
       .uc2rb_desc_3_xuser_14_reg		(uc2rb_desc_3_xuser_14_reg[31:0]),
       .uc2rb_desc_3_xuser_15_reg		(uc2rb_desc_3_xuser_15_reg[31:0]),
       .uc2rb_desc_4_xuser_0_reg			(uc2rb_desc_4_xuser_0_reg[31:0]),
       .uc2rb_desc_4_xuser_1_reg			(uc2rb_desc_4_xuser_1_reg[31:0]),
       .uc2rb_desc_4_xuser_2_reg			(uc2rb_desc_4_xuser_2_reg[31:0]),
       .uc2rb_desc_4_xuser_3_reg			(uc2rb_desc_4_xuser_3_reg[31:0]),
       .uc2rb_desc_4_xuser_4_reg			(uc2rb_desc_4_xuser_4_reg[31:0]),
       .uc2rb_desc_4_xuser_5_reg			(uc2rb_desc_4_xuser_5_reg[31:0]),
       .uc2rb_desc_4_xuser_6_reg			(uc2rb_desc_4_xuser_6_reg[31:0]),
       .uc2rb_desc_4_xuser_7_reg			(uc2rb_desc_4_xuser_7_reg[31:0]),
       .uc2rb_desc_4_xuser_8_reg			(uc2rb_desc_4_xuser_8_reg[31:0]),
       .uc2rb_desc_4_xuser_9_reg			(uc2rb_desc_4_xuser_9_reg[31:0]),
       .uc2rb_desc_4_xuser_10_reg		(uc2rb_desc_4_xuser_10_reg[31:0]),
       .uc2rb_desc_4_xuser_11_reg		(uc2rb_desc_4_xuser_11_reg[31:0]),
       .uc2rb_desc_4_xuser_12_reg		(uc2rb_desc_4_xuser_12_reg[31:0]),
       .uc2rb_desc_4_xuser_13_reg		(uc2rb_desc_4_xuser_13_reg[31:0]),
       .uc2rb_desc_4_xuser_14_reg		(uc2rb_desc_4_xuser_14_reg[31:0]),
       .uc2rb_desc_4_xuser_15_reg		(uc2rb_desc_4_xuser_15_reg[31:0]),
       .uc2rb_desc_5_xuser_0_reg			(uc2rb_desc_5_xuser_0_reg[31:0]),
       .uc2rb_desc_5_xuser_1_reg			(uc2rb_desc_5_xuser_1_reg[31:0]),
       .uc2rb_desc_5_xuser_2_reg			(uc2rb_desc_5_xuser_2_reg[31:0]),
       .uc2rb_desc_5_xuser_3_reg			(uc2rb_desc_5_xuser_3_reg[31:0]),
       .uc2rb_desc_5_xuser_4_reg			(uc2rb_desc_5_xuser_4_reg[31:0]),
       .uc2rb_desc_5_xuser_5_reg			(uc2rb_desc_5_xuser_5_reg[31:0]),
       .uc2rb_desc_5_xuser_6_reg			(uc2rb_desc_5_xuser_6_reg[31:0]),
       .uc2rb_desc_5_xuser_7_reg			(uc2rb_desc_5_xuser_7_reg[31:0]),
       .uc2rb_desc_5_xuser_8_reg			(uc2rb_desc_5_xuser_8_reg[31:0]),
       .uc2rb_desc_5_xuser_9_reg			(uc2rb_desc_5_xuser_9_reg[31:0]),
       .uc2rb_desc_5_xuser_10_reg		(uc2rb_desc_5_xuser_10_reg[31:0]),
       .uc2rb_desc_5_xuser_11_reg		(uc2rb_desc_5_xuser_11_reg[31:0]),
       .uc2rb_desc_5_xuser_12_reg		(uc2rb_desc_5_xuser_12_reg[31:0]),
       .uc2rb_desc_5_xuser_13_reg		(uc2rb_desc_5_xuser_13_reg[31:0]),
       .uc2rb_desc_5_xuser_14_reg		(uc2rb_desc_5_xuser_14_reg[31:0]),
       .uc2rb_desc_5_xuser_15_reg		(uc2rb_desc_5_xuser_15_reg[31:0]),
       .uc2rb_desc_6_xuser_0_reg			(uc2rb_desc_6_xuser_0_reg[31:0]),
       .uc2rb_desc_6_xuser_1_reg			(uc2rb_desc_6_xuser_1_reg[31:0]),
       .uc2rb_desc_6_xuser_2_reg			(uc2rb_desc_6_xuser_2_reg[31:0]),
       .uc2rb_desc_6_xuser_3_reg			(uc2rb_desc_6_xuser_3_reg[31:0]),
       .uc2rb_desc_6_xuser_4_reg			(uc2rb_desc_6_xuser_4_reg[31:0]),
       .uc2rb_desc_6_xuser_5_reg			(uc2rb_desc_6_xuser_5_reg[31:0]),
       .uc2rb_desc_6_xuser_6_reg			(uc2rb_desc_6_xuser_6_reg[31:0]),
       .uc2rb_desc_6_xuser_7_reg			(uc2rb_desc_6_xuser_7_reg[31:0]),
       .uc2rb_desc_6_xuser_8_reg			(uc2rb_desc_6_xuser_8_reg[31:0]),
       .uc2rb_desc_6_xuser_9_reg			(uc2rb_desc_6_xuser_9_reg[31:0]),
       .uc2rb_desc_6_xuser_10_reg		(uc2rb_desc_6_xuser_10_reg[31:0]),
       .uc2rb_desc_6_xuser_11_reg		(uc2rb_desc_6_xuser_11_reg[31:0]),
       .uc2rb_desc_6_xuser_12_reg		(uc2rb_desc_6_xuser_12_reg[31:0]),
       .uc2rb_desc_6_xuser_13_reg		(uc2rb_desc_6_xuser_13_reg[31:0]),
       .uc2rb_desc_6_xuser_14_reg		(uc2rb_desc_6_xuser_14_reg[31:0]),
       .uc2rb_desc_6_xuser_15_reg		(uc2rb_desc_6_xuser_15_reg[31:0]),
       .uc2rb_desc_7_xuser_0_reg			(uc2rb_desc_7_xuser_0_reg[31:0]),
       .uc2rb_desc_7_xuser_1_reg			(uc2rb_desc_7_xuser_1_reg[31:0]),
       .uc2rb_desc_7_xuser_2_reg			(uc2rb_desc_7_xuser_2_reg[31:0]),
       .uc2rb_desc_7_xuser_3_reg			(uc2rb_desc_7_xuser_3_reg[31:0]),
       .uc2rb_desc_7_xuser_4_reg			(uc2rb_desc_7_xuser_4_reg[31:0]),
       .uc2rb_desc_7_xuser_5_reg			(uc2rb_desc_7_xuser_5_reg[31:0]),
       .uc2rb_desc_7_xuser_6_reg			(uc2rb_desc_7_xuser_6_reg[31:0]),
       .uc2rb_desc_7_xuser_7_reg			(uc2rb_desc_7_xuser_7_reg[31:0]),
       .uc2rb_desc_7_xuser_8_reg			(uc2rb_desc_7_xuser_8_reg[31:0]),
       .uc2rb_desc_7_xuser_9_reg			(uc2rb_desc_7_xuser_9_reg[31:0]),
       .uc2rb_desc_7_xuser_10_reg		(uc2rb_desc_7_xuser_10_reg[31:0]),
       .uc2rb_desc_7_xuser_11_reg		(uc2rb_desc_7_xuser_11_reg[31:0]),
       .uc2rb_desc_7_xuser_12_reg		(uc2rb_desc_7_xuser_12_reg[31:0]),
       .uc2rb_desc_7_xuser_13_reg		(uc2rb_desc_7_xuser_13_reg[31:0]),
       .uc2rb_desc_7_xuser_14_reg		(uc2rb_desc_7_xuser_14_reg[31:0]),
       .uc2rb_desc_7_xuser_15_reg		(uc2rb_desc_7_xuser_15_reg[31:0]),
       .uc2rb_desc_8_xuser_0_reg			(uc2rb_desc_8_xuser_0_reg[31:0]),
       .uc2rb_desc_8_xuser_1_reg			(uc2rb_desc_8_xuser_1_reg[31:0]),
       .uc2rb_desc_8_xuser_2_reg			(uc2rb_desc_8_xuser_2_reg[31:0]),
       .uc2rb_desc_8_xuser_3_reg			(uc2rb_desc_8_xuser_3_reg[31:0]),
       .uc2rb_desc_8_xuser_4_reg			(uc2rb_desc_8_xuser_4_reg[31:0]),
       .uc2rb_desc_8_xuser_5_reg			(uc2rb_desc_8_xuser_5_reg[31:0]),
       .uc2rb_desc_8_xuser_6_reg			(uc2rb_desc_8_xuser_6_reg[31:0]),
       .uc2rb_desc_8_xuser_7_reg			(uc2rb_desc_8_xuser_7_reg[31:0]),
       .uc2rb_desc_8_xuser_8_reg			(uc2rb_desc_8_xuser_8_reg[31:0]),
       .uc2rb_desc_8_xuser_9_reg			(uc2rb_desc_8_xuser_9_reg[31:0]),
       .uc2rb_desc_8_xuser_10_reg		(uc2rb_desc_8_xuser_10_reg[31:0]),
       .uc2rb_desc_8_xuser_11_reg		(uc2rb_desc_8_xuser_11_reg[31:0]),
       .uc2rb_desc_8_xuser_12_reg		(uc2rb_desc_8_xuser_12_reg[31:0]),
       .uc2rb_desc_8_xuser_13_reg		(uc2rb_desc_8_xuser_13_reg[31:0]),
       .uc2rb_desc_8_xuser_14_reg		(uc2rb_desc_8_xuser_14_reg[31:0]),
       .uc2rb_desc_8_xuser_15_reg		(uc2rb_desc_8_xuser_15_reg[31:0]),
       .uc2rb_desc_9_xuser_0_reg			(uc2rb_desc_9_xuser_0_reg[31:0]),
       .uc2rb_desc_9_xuser_1_reg			(uc2rb_desc_9_xuser_1_reg[31:0]),
       .uc2rb_desc_9_xuser_2_reg			(uc2rb_desc_9_xuser_2_reg[31:0]),
       .uc2rb_desc_9_xuser_3_reg			(uc2rb_desc_9_xuser_3_reg[31:0]),
       .uc2rb_desc_9_xuser_4_reg			(uc2rb_desc_9_xuser_4_reg[31:0]),
       .uc2rb_desc_9_xuser_5_reg			(uc2rb_desc_9_xuser_5_reg[31:0]),
       .uc2rb_desc_9_xuser_6_reg			(uc2rb_desc_9_xuser_6_reg[31:0]),
       .uc2rb_desc_9_xuser_7_reg			(uc2rb_desc_9_xuser_7_reg[31:0]),
       .uc2rb_desc_9_xuser_8_reg			(uc2rb_desc_9_xuser_8_reg[31:0]),
       .uc2rb_desc_9_xuser_9_reg			(uc2rb_desc_9_xuser_9_reg[31:0]),
       .uc2rb_desc_9_xuser_10_reg		(uc2rb_desc_9_xuser_10_reg[31:0]),
       .uc2rb_desc_9_xuser_11_reg		(uc2rb_desc_9_xuser_11_reg[31:0]),
       .uc2rb_desc_9_xuser_12_reg		(uc2rb_desc_9_xuser_12_reg[31:0]),
       .uc2rb_desc_9_xuser_13_reg		(uc2rb_desc_9_xuser_13_reg[31:0]),
       .uc2rb_desc_9_xuser_14_reg		(uc2rb_desc_9_xuser_14_reg[31:0]),
       .uc2rb_desc_9_xuser_15_reg		(uc2rb_desc_9_xuser_15_reg[31:0]),
       .uc2rb_desc_10_xuser_0_reg		(uc2rb_desc_10_xuser_0_reg[31:0]),
       .uc2rb_desc_10_xuser_1_reg		(uc2rb_desc_10_xuser_1_reg[31:0]),
       .uc2rb_desc_10_xuser_2_reg		(uc2rb_desc_10_xuser_2_reg[31:0]),
       .uc2rb_desc_10_xuser_3_reg		(uc2rb_desc_10_xuser_3_reg[31:0]),
       .uc2rb_desc_10_xuser_4_reg		(uc2rb_desc_10_xuser_4_reg[31:0]),
       .uc2rb_desc_10_xuser_5_reg		(uc2rb_desc_10_xuser_5_reg[31:0]),
       .uc2rb_desc_10_xuser_6_reg		(uc2rb_desc_10_xuser_6_reg[31:0]),
       .uc2rb_desc_10_xuser_7_reg		(uc2rb_desc_10_xuser_7_reg[31:0]),
       .uc2rb_desc_10_xuser_8_reg		(uc2rb_desc_10_xuser_8_reg[31:0]),
       .uc2rb_desc_10_xuser_9_reg		(uc2rb_desc_10_xuser_9_reg[31:0]),
       .uc2rb_desc_10_xuser_10_reg		(uc2rb_desc_10_xuser_10_reg[31:0]),
       .uc2rb_desc_10_xuser_11_reg		(uc2rb_desc_10_xuser_11_reg[31:0]),
       .uc2rb_desc_10_xuser_12_reg		(uc2rb_desc_10_xuser_12_reg[31:0]),
       .uc2rb_desc_10_xuser_13_reg		(uc2rb_desc_10_xuser_13_reg[31:0]),
       .uc2rb_desc_10_xuser_14_reg		(uc2rb_desc_10_xuser_14_reg[31:0]),
       .uc2rb_desc_10_xuser_15_reg		(uc2rb_desc_10_xuser_15_reg[31:0]),
       .uc2rb_desc_11_xuser_0_reg		(uc2rb_desc_11_xuser_0_reg[31:0]),
       .uc2rb_desc_11_xuser_1_reg		(uc2rb_desc_11_xuser_1_reg[31:0]),
       .uc2rb_desc_11_xuser_2_reg		(uc2rb_desc_11_xuser_2_reg[31:0]),
       .uc2rb_desc_11_xuser_3_reg		(uc2rb_desc_11_xuser_3_reg[31:0]),
       .uc2rb_desc_11_xuser_4_reg		(uc2rb_desc_11_xuser_4_reg[31:0]),
       .uc2rb_desc_11_xuser_5_reg		(uc2rb_desc_11_xuser_5_reg[31:0]),
       .uc2rb_desc_11_xuser_6_reg		(uc2rb_desc_11_xuser_6_reg[31:0]),
       .uc2rb_desc_11_xuser_7_reg		(uc2rb_desc_11_xuser_7_reg[31:0]),
       .uc2rb_desc_11_xuser_8_reg		(uc2rb_desc_11_xuser_8_reg[31:0]),
       .uc2rb_desc_11_xuser_9_reg		(uc2rb_desc_11_xuser_9_reg[31:0]),
       .uc2rb_desc_11_xuser_10_reg		(uc2rb_desc_11_xuser_10_reg[31:0]),
       .uc2rb_desc_11_xuser_11_reg		(uc2rb_desc_11_xuser_11_reg[31:0]),
       .uc2rb_desc_11_xuser_12_reg		(uc2rb_desc_11_xuser_12_reg[31:0]),
       .uc2rb_desc_11_xuser_13_reg		(uc2rb_desc_11_xuser_13_reg[31:0]),
       .uc2rb_desc_11_xuser_14_reg		(uc2rb_desc_11_xuser_14_reg[31:0]),
       .uc2rb_desc_11_xuser_15_reg		(uc2rb_desc_11_xuser_15_reg[31:0]),
       .uc2rb_desc_12_xuser_0_reg		(uc2rb_desc_12_xuser_0_reg[31:0]),
       .uc2rb_desc_12_xuser_1_reg		(uc2rb_desc_12_xuser_1_reg[31:0]),
       .uc2rb_desc_12_xuser_2_reg		(uc2rb_desc_12_xuser_2_reg[31:0]),
       .uc2rb_desc_12_xuser_3_reg		(uc2rb_desc_12_xuser_3_reg[31:0]),
       .uc2rb_desc_12_xuser_4_reg		(uc2rb_desc_12_xuser_4_reg[31:0]),
       .uc2rb_desc_12_xuser_5_reg		(uc2rb_desc_12_xuser_5_reg[31:0]),
       .uc2rb_desc_12_xuser_6_reg		(uc2rb_desc_12_xuser_6_reg[31:0]),
       .uc2rb_desc_12_xuser_7_reg		(uc2rb_desc_12_xuser_7_reg[31:0]),
       .uc2rb_desc_12_xuser_8_reg		(uc2rb_desc_12_xuser_8_reg[31:0]),
       .uc2rb_desc_12_xuser_9_reg		(uc2rb_desc_12_xuser_9_reg[31:0]),
       .uc2rb_desc_12_xuser_10_reg		(uc2rb_desc_12_xuser_10_reg[31:0]),
       .uc2rb_desc_12_xuser_11_reg		(uc2rb_desc_12_xuser_11_reg[31:0]),
       .uc2rb_desc_12_xuser_12_reg		(uc2rb_desc_12_xuser_12_reg[31:0]),
       .uc2rb_desc_12_xuser_13_reg		(uc2rb_desc_12_xuser_13_reg[31:0]),
       .uc2rb_desc_12_xuser_14_reg		(uc2rb_desc_12_xuser_14_reg[31:0]),
       .uc2rb_desc_12_xuser_15_reg		(uc2rb_desc_12_xuser_15_reg[31:0]),
       .uc2rb_desc_13_xuser_0_reg		(uc2rb_desc_13_xuser_0_reg[31:0]),
       .uc2rb_desc_13_xuser_1_reg		(uc2rb_desc_13_xuser_1_reg[31:0]),
       .uc2rb_desc_13_xuser_2_reg		(uc2rb_desc_13_xuser_2_reg[31:0]),
       .uc2rb_desc_13_xuser_3_reg		(uc2rb_desc_13_xuser_3_reg[31:0]),
       .uc2rb_desc_13_xuser_4_reg		(uc2rb_desc_13_xuser_4_reg[31:0]),
       .uc2rb_desc_13_xuser_5_reg		(uc2rb_desc_13_xuser_5_reg[31:0]),
       .uc2rb_desc_13_xuser_6_reg		(uc2rb_desc_13_xuser_6_reg[31:0]),
       .uc2rb_desc_13_xuser_7_reg		(uc2rb_desc_13_xuser_7_reg[31:0]),
       .uc2rb_desc_13_xuser_8_reg		(uc2rb_desc_13_xuser_8_reg[31:0]),
       .uc2rb_desc_13_xuser_9_reg		(uc2rb_desc_13_xuser_9_reg[31:0]),
       .uc2rb_desc_13_xuser_10_reg		(uc2rb_desc_13_xuser_10_reg[31:0]),
       .uc2rb_desc_13_xuser_11_reg		(uc2rb_desc_13_xuser_11_reg[31:0]),
       .uc2rb_desc_13_xuser_12_reg		(uc2rb_desc_13_xuser_12_reg[31:0]),
       .uc2rb_desc_13_xuser_13_reg		(uc2rb_desc_13_xuser_13_reg[31:0]),
       .uc2rb_desc_13_xuser_14_reg		(uc2rb_desc_13_xuser_14_reg[31:0]),
       .uc2rb_desc_13_xuser_15_reg		(uc2rb_desc_13_xuser_15_reg[31:0]),
       .uc2rb_desc_14_xuser_0_reg		(uc2rb_desc_14_xuser_0_reg[31:0]),
       .uc2rb_desc_14_xuser_1_reg		(uc2rb_desc_14_xuser_1_reg[31:0]),
       .uc2rb_desc_14_xuser_2_reg		(uc2rb_desc_14_xuser_2_reg[31:0]),
       .uc2rb_desc_14_xuser_3_reg		(uc2rb_desc_14_xuser_3_reg[31:0]),
       .uc2rb_desc_14_xuser_4_reg		(uc2rb_desc_14_xuser_4_reg[31:0]),
       .uc2rb_desc_14_xuser_5_reg		(uc2rb_desc_14_xuser_5_reg[31:0]),
       .uc2rb_desc_14_xuser_6_reg		(uc2rb_desc_14_xuser_6_reg[31:0]),
       .uc2rb_desc_14_xuser_7_reg		(uc2rb_desc_14_xuser_7_reg[31:0]),
       .uc2rb_desc_14_xuser_8_reg		(uc2rb_desc_14_xuser_8_reg[31:0]),
       .uc2rb_desc_14_xuser_9_reg		(uc2rb_desc_14_xuser_9_reg[31:0]),
       .uc2rb_desc_14_xuser_10_reg		(uc2rb_desc_14_xuser_10_reg[31:0]),
       .uc2rb_desc_14_xuser_11_reg		(uc2rb_desc_14_xuser_11_reg[31:0]),
       .uc2rb_desc_14_xuser_12_reg		(uc2rb_desc_14_xuser_12_reg[31:0]),
       .uc2rb_desc_14_xuser_13_reg		(uc2rb_desc_14_xuser_13_reg[31:0]),
       .uc2rb_desc_14_xuser_14_reg		(uc2rb_desc_14_xuser_14_reg[31:0]),
       .uc2rb_desc_14_xuser_15_reg		(uc2rb_desc_14_xuser_15_reg[31:0]),
       .uc2rb_desc_15_xuser_0_reg		(uc2rb_desc_15_xuser_0_reg[31:0]),
       .uc2rb_desc_15_xuser_1_reg		(uc2rb_desc_15_xuser_1_reg[31:0]),
       .uc2rb_desc_15_xuser_2_reg		(uc2rb_desc_15_xuser_2_reg[31:0]),
       .uc2rb_desc_15_xuser_3_reg		(uc2rb_desc_15_xuser_3_reg[31:0]),
       .uc2rb_desc_15_xuser_4_reg		(uc2rb_desc_15_xuser_4_reg[31:0]),
       .uc2rb_desc_15_xuser_5_reg		(uc2rb_desc_15_xuser_5_reg[31:0]),
       .uc2rb_desc_15_xuser_6_reg		(uc2rb_desc_15_xuser_6_reg[31:0]),
       .uc2rb_desc_15_xuser_7_reg		(uc2rb_desc_15_xuser_7_reg[31:0]),
       .uc2rb_desc_15_xuser_8_reg		(uc2rb_desc_15_xuser_8_reg[31:0]),
       .uc2rb_desc_15_xuser_9_reg		(uc2rb_desc_15_xuser_9_reg[31:0]),
       .uc2rb_desc_15_xuser_10_reg		(uc2rb_desc_15_xuser_10_reg[31:0]),
       .uc2rb_desc_15_xuser_11_reg		(uc2rb_desc_15_xuser_11_reg[31:0]),
       .uc2rb_desc_15_xuser_12_reg		(uc2rb_desc_15_xuser_12_reg[31:0]),
       .uc2rb_desc_15_xuser_13_reg		(uc2rb_desc_15_xuser_13_reg[31:0]),
       .uc2rb_desc_15_xuser_14_reg		(uc2rb_desc_15_xuser_14_reg[31:0]),
       .uc2rb_desc_15_xuser_15_reg		(uc2rb_desc_15_xuser_15_reg[31:0]),
       .uc2rb_intr_error_status_reg_we	(uc2rb_intr_error_status_reg_we[31:0]),
       .uc2rb_ownership_reg_we			(uc2rb_ownership_reg_we[31:0]),
       .uc2rb_intr_comp_status_reg_we	(uc2rb_intr_comp_status_reg_we[31:0]),
       .uc2rb_status_resp_reg_we			(uc2rb_status_resp_reg_we[31:0]),
       .uc2rb_status_busy_reg_we			(uc2rb_status_busy_reg_we[31:0]),
       .uc2rb_desc_0_xuser_0_reg_we		(uc2rb_desc_0_xuser_0_reg_we[31:0]),
       .uc2rb_desc_0_xuser_1_reg_we		(uc2rb_desc_0_xuser_1_reg_we[31:0]),
       .uc2rb_desc_0_xuser_2_reg_we		(uc2rb_desc_0_xuser_2_reg_we[31:0]),
       .uc2rb_desc_0_xuser_3_reg_we		(uc2rb_desc_0_xuser_3_reg_we[31:0]),
       .uc2rb_desc_0_xuser_4_reg_we		(uc2rb_desc_0_xuser_4_reg_we[31:0]),
       .uc2rb_desc_0_xuser_5_reg_we		(uc2rb_desc_0_xuser_5_reg_we[31:0]),
       .uc2rb_desc_0_xuser_6_reg_we		(uc2rb_desc_0_xuser_6_reg_we[31:0]),
       .uc2rb_desc_0_xuser_7_reg_we		(uc2rb_desc_0_xuser_7_reg_we[31:0]),
       .uc2rb_desc_0_xuser_8_reg_we		(uc2rb_desc_0_xuser_8_reg_we[31:0]),
       .uc2rb_desc_0_xuser_9_reg_we		(uc2rb_desc_0_xuser_9_reg_we[31:0]),
       .uc2rb_desc_0_xuser_10_reg_we		(uc2rb_desc_0_xuser_10_reg_we[31:0]),
       .uc2rb_desc_0_xuser_11_reg_we		(uc2rb_desc_0_xuser_11_reg_we[31:0]),
       .uc2rb_desc_0_xuser_12_reg_we		(uc2rb_desc_0_xuser_12_reg_we[31:0]),
       .uc2rb_desc_0_xuser_13_reg_we		(uc2rb_desc_0_xuser_13_reg_we[31:0]),
       .uc2rb_desc_0_xuser_14_reg_we		(uc2rb_desc_0_xuser_14_reg_we[31:0]),
       .uc2rb_desc_0_xuser_15_reg_we		(uc2rb_desc_0_xuser_15_reg_we[31:0]),
       .uc2rb_desc_1_xuser_0_reg_we		(uc2rb_desc_1_xuser_0_reg_we[31:0]),
       .uc2rb_desc_1_xuser_1_reg_we		(uc2rb_desc_1_xuser_1_reg_we[31:0]),
       .uc2rb_desc_1_xuser_2_reg_we		(uc2rb_desc_1_xuser_2_reg_we[31:0]),
       .uc2rb_desc_1_xuser_3_reg_we		(uc2rb_desc_1_xuser_3_reg_we[31:0]),
       .uc2rb_desc_1_xuser_4_reg_we		(uc2rb_desc_1_xuser_4_reg_we[31:0]),
       .uc2rb_desc_1_xuser_5_reg_we		(uc2rb_desc_1_xuser_5_reg_we[31:0]),
       .uc2rb_desc_1_xuser_6_reg_we		(uc2rb_desc_1_xuser_6_reg_we[31:0]),
       .uc2rb_desc_1_xuser_7_reg_we		(uc2rb_desc_1_xuser_7_reg_we[31:0]),
       .uc2rb_desc_1_xuser_8_reg_we		(uc2rb_desc_1_xuser_8_reg_we[31:0]),
       .uc2rb_desc_1_xuser_9_reg_we		(uc2rb_desc_1_xuser_9_reg_we[31:0]),
       .uc2rb_desc_1_xuser_10_reg_we		(uc2rb_desc_1_xuser_10_reg_we[31:0]),
       .uc2rb_desc_1_xuser_11_reg_we		(uc2rb_desc_1_xuser_11_reg_we[31:0]),
       .uc2rb_desc_1_xuser_12_reg_we		(uc2rb_desc_1_xuser_12_reg_we[31:0]),
       .uc2rb_desc_1_xuser_13_reg_we		(uc2rb_desc_1_xuser_13_reg_we[31:0]),
       .uc2rb_desc_1_xuser_14_reg_we		(uc2rb_desc_1_xuser_14_reg_we[31:0]),
       .uc2rb_desc_1_xuser_15_reg_we		(uc2rb_desc_1_xuser_15_reg_we[31:0]),
       .uc2rb_desc_2_xuser_0_reg_we		(uc2rb_desc_2_xuser_0_reg_we[31:0]),
       .uc2rb_desc_2_xuser_1_reg_we		(uc2rb_desc_2_xuser_1_reg_we[31:0]),
       .uc2rb_desc_2_xuser_2_reg_we		(uc2rb_desc_2_xuser_2_reg_we[31:0]),
       .uc2rb_desc_2_xuser_3_reg_we		(uc2rb_desc_2_xuser_3_reg_we[31:0]),
       .uc2rb_desc_2_xuser_4_reg_we		(uc2rb_desc_2_xuser_4_reg_we[31:0]),
       .uc2rb_desc_2_xuser_5_reg_we		(uc2rb_desc_2_xuser_5_reg_we[31:0]),
       .uc2rb_desc_2_xuser_6_reg_we		(uc2rb_desc_2_xuser_6_reg_we[31:0]),
       .uc2rb_desc_2_xuser_7_reg_we		(uc2rb_desc_2_xuser_7_reg_we[31:0]),
       .uc2rb_desc_2_xuser_8_reg_we		(uc2rb_desc_2_xuser_8_reg_we[31:0]),
       .uc2rb_desc_2_xuser_9_reg_we		(uc2rb_desc_2_xuser_9_reg_we[31:0]),
       .uc2rb_desc_2_xuser_10_reg_we		(uc2rb_desc_2_xuser_10_reg_we[31:0]),
       .uc2rb_desc_2_xuser_11_reg_we		(uc2rb_desc_2_xuser_11_reg_we[31:0]),
       .uc2rb_desc_2_xuser_12_reg_we		(uc2rb_desc_2_xuser_12_reg_we[31:0]),
       .uc2rb_desc_2_xuser_13_reg_we		(uc2rb_desc_2_xuser_13_reg_we[31:0]),
       .uc2rb_desc_2_xuser_14_reg_we		(uc2rb_desc_2_xuser_14_reg_we[31:0]),
       .uc2rb_desc_2_xuser_15_reg_we		(uc2rb_desc_2_xuser_15_reg_we[31:0]),
       .uc2rb_desc_3_xuser_0_reg_we		(uc2rb_desc_3_xuser_0_reg_we[31:0]),
       .uc2rb_desc_3_xuser_1_reg_we		(uc2rb_desc_3_xuser_1_reg_we[31:0]),
       .uc2rb_desc_3_xuser_2_reg_we		(uc2rb_desc_3_xuser_2_reg_we[31:0]),
       .uc2rb_desc_3_xuser_3_reg_we		(uc2rb_desc_3_xuser_3_reg_we[31:0]),
       .uc2rb_desc_3_xuser_4_reg_we		(uc2rb_desc_3_xuser_4_reg_we[31:0]),
       .uc2rb_desc_3_xuser_5_reg_we		(uc2rb_desc_3_xuser_5_reg_we[31:0]),
       .uc2rb_desc_3_xuser_6_reg_we		(uc2rb_desc_3_xuser_6_reg_we[31:0]),
       .uc2rb_desc_3_xuser_7_reg_we		(uc2rb_desc_3_xuser_7_reg_we[31:0]),
       .uc2rb_desc_3_xuser_8_reg_we		(uc2rb_desc_3_xuser_8_reg_we[31:0]),
       .uc2rb_desc_3_xuser_9_reg_we		(uc2rb_desc_3_xuser_9_reg_we[31:0]),
       .uc2rb_desc_3_xuser_10_reg_we		(uc2rb_desc_3_xuser_10_reg_we[31:0]),
       .uc2rb_desc_3_xuser_11_reg_we		(uc2rb_desc_3_xuser_11_reg_we[31:0]),
       .uc2rb_desc_3_xuser_12_reg_we		(uc2rb_desc_3_xuser_12_reg_we[31:0]),
       .uc2rb_desc_3_xuser_13_reg_we		(uc2rb_desc_3_xuser_13_reg_we[31:0]),
       .uc2rb_desc_3_xuser_14_reg_we		(uc2rb_desc_3_xuser_14_reg_we[31:0]),
       .uc2rb_desc_3_xuser_15_reg_we		(uc2rb_desc_3_xuser_15_reg_we[31:0]),
       .uc2rb_desc_4_xuser_0_reg_we		(uc2rb_desc_4_xuser_0_reg_we[31:0]),
       .uc2rb_desc_4_xuser_1_reg_we		(uc2rb_desc_4_xuser_1_reg_we[31:0]),
       .uc2rb_desc_4_xuser_2_reg_we		(uc2rb_desc_4_xuser_2_reg_we[31:0]),
       .uc2rb_desc_4_xuser_3_reg_we		(uc2rb_desc_4_xuser_3_reg_we[31:0]),
       .uc2rb_desc_4_xuser_4_reg_we		(uc2rb_desc_4_xuser_4_reg_we[31:0]),
       .uc2rb_desc_4_xuser_5_reg_we		(uc2rb_desc_4_xuser_5_reg_we[31:0]),
       .uc2rb_desc_4_xuser_6_reg_we		(uc2rb_desc_4_xuser_6_reg_we[31:0]),
       .uc2rb_desc_4_xuser_7_reg_we		(uc2rb_desc_4_xuser_7_reg_we[31:0]),
       .uc2rb_desc_4_xuser_8_reg_we		(uc2rb_desc_4_xuser_8_reg_we[31:0]),
       .uc2rb_desc_4_xuser_9_reg_we		(uc2rb_desc_4_xuser_9_reg_we[31:0]),
       .uc2rb_desc_4_xuser_10_reg_we		(uc2rb_desc_4_xuser_10_reg_we[31:0]),
       .uc2rb_desc_4_xuser_11_reg_we		(uc2rb_desc_4_xuser_11_reg_we[31:0]),
       .uc2rb_desc_4_xuser_12_reg_we		(uc2rb_desc_4_xuser_12_reg_we[31:0]),
       .uc2rb_desc_4_xuser_13_reg_we		(uc2rb_desc_4_xuser_13_reg_we[31:0]),
       .uc2rb_desc_4_xuser_14_reg_we		(uc2rb_desc_4_xuser_14_reg_we[31:0]),
       .uc2rb_desc_4_xuser_15_reg_we		(uc2rb_desc_4_xuser_15_reg_we[31:0]),
       .uc2rb_desc_5_xuser_0_reg_we		(uc2rb_desc_5_xuser_0_reg_we[31:0]),
       .uc2rb_desc_5_xuser_1_reg_we		(uc2rb_desc_5_xuser_1_reg_we[31:0]),
       .uc2rb_desc_5_xuser_2_reg_we		(uc2rb_desc_5_xuser_2_reg_we[31:0]),
       .uc2rb_desc_5_xuser_3_reg_we		(uc2rb_desc_5_xuser_3_reg_we[31:0]),
       .uc2rb_desc_5_xuser_4_reg_we		(uc2rb_desc_5_xuser_4_reg_we[31:0]),
       .uc2rb_desc_5_xuser_5_reg_we		(uc2rb_desc_5_xuser_5_reg_we[31:0]),
       .uc2rb_desc_5_xuser_6_reg_we		(uc2rb_desc_5_xuser_6_reg_we[31:0]),
       .uc2rb_desc_5_xuser_7_reg_we		(uc2rb_desc_5_xuser_7_reg_we[31:0]),
       .uc2rb_desc_5_xuser_8_reg_we		(uc2rb_desc_5_xuser_8_reg_we[31:0]),
       .uc2rb_desc_5_xuser_9_reg_we		(uc2rb_desc_5_xuser_9_reg_we[31:0]),
       .uc2rb_desc_5_xuser_10_reg_we		(uc2rb_desc_5_xuser_10_reg_we[31:0]),
       .uc2rb_desc_5_xuser_11_reg_we		(uc2rb_desc_5_xuser_11_reg_we[31:0]),
       .uc2rb_desc_5_xuser_12_reg_we		(uc2rb_desc_5_xuser_12_reg_we[31:0]),
       .uc2rb_desc_5_xuser_13_reg_we		(uc2rb_desc_5_xuser_13_reg_we[31:0]),
       .uc2rb_desc_5_xuser_14_reg_we		(uc2rb_desc_5_xuser_14_reg_we[31:0]),
       .uc2rb_desc_5_xuser_15_reg_we		(uc2rb_desc_5_xuser_15_reg_we[31:0]),
       .uc2rb_desc_6_xuser_0_reg_we		(uc2rb_desc_6_xuser_0_reg_we[31:0]),
       .uc2rb_desc_6_xuser_1_reg_we		(uc2rb_desc_6_xuser_1_reg_we[31:0]),
       .uc2rb_desc_6_xuser_2_reg_we		(uc2rb_desc_6_xuser_2_reg_we[31:0]),
       .uc2rb_desc_6_xuser_3_reg_we		(uc2rb_desc_6_xuser_3_reg_we[31:0]),
       .uc2rb_desc_6_xuser_4_reg_we		(uc2rb_desc_6_xuser_4_reg_we[31:0]),
       .uc2rb_desc_6_xuser_5_reg_we		(uc2rb_desc_6_xuser_5_reg_we[31:0]),
       .uc2rb_desc_6_xuser_6_reg_we		(uc2rb_desc_6_xuser_6_reg_we[31:0]),
       .uc2rb_desc_6_xuser_7_reg_we		(uc2rb_desc_6_xuser_7_reg_we[31:0]),
       .uc2rb_desc_6_xuser_8_reg_we		(uc2rb_desc_6_xuser_8_reg_we[31:0]),
       .uc2rb_desc_6_xuser_9_reg_we		(uc2rb_desc_6_xuser_9_reg_we[31:0]),
       .uc2rb_desc_6_xuser_10_reg_we		(uc2rb_desc_6_xuser_10_reg_we[31:0]),
       .uc2rb_desc_6_xuser_11_reg_we		(uc2rb_desc_6_xuser_11_reg_we[31:0]),
       .uc2rb_desc_6_xuser_12_reg_we		(uc2rb_desc_6_xuser_12_reg_we[31:0]),
       .uc2rb_desc_6_xuser_13_reg_we		(uc2rb_desc_6_xuser_13_reg_we[31:0]),
       .uc2rb_desc_6_xuser_14_reg_we		(uc2rb_desc_6_xuser_14_reg_we[31:0]),
       .uc2rb_desc_6_xuser_15_reg_we		(uc2rb_desc_6_xuser_15_reg_we[31:0]),
       .uc2rb_desc_7_xuser_0_reg_we		(uc2rb_desc_7_xuser_0_reg_we[31:0]),
       .uc2rb_desc_7_xuser_1_reg_we		(uc2rb_desc_7_xuser_1_reg_we[31:0]),
       .uc2rb_desc_7_xuser_2_reg_we		(uc2rb_desc_7_xuser_2_reg_we[31:0]),
       .uc2rb_desc_7_xuser_3_reg_we		(uc2rb_desc_7_xuser_3_reg_we[31:0]),
       .uc2rb_desc_7_xuser_4_reg_we		(uc2rb_desc_7_xuser_4_reg_we[31:0]),
       .uc2rb_desc_7_xuser_5_reg_we		(uc2rb_desc_7_xuser_5_reg_we[31:0]),
       .uc2rb_desc_7_xuser_6_reg_we		(uc2rb_desc_7_xuser_6_reg_we[31:0]),
       .uc2rb_desc_7_xuser_7_reg_we		(uc2rb_desc_7_xuser_7_reg_we[31:0]),
       .uc2rb_desc_7_xuser_8_reg_we		(uc2rb_desc_7_xuser_8_reg_we[31:0]),
       .uc2rb_desc_7_xuser_9_reg_we		(uc2rb_desc_7_xuser_9_reg_we[31:0]),
       .uc2rb_desc_7_xuser_10_reg_we		(uc2rb_desc_7_xuser_10_reg_we[31:0]),
       .uc2rb_desc_7_xuser_11_reg_we		(uc2rb_desc_7_xuser_11_reg_we[31:0]),
       .uc2rb_desc_7_xuser_12_reg_we		(uc2rb_desc_7_xuser_12_reg_we[31:0]),
       .uc2rb_desc_7_xuser_13_reg_we		(uc2rb_desc_7_xuser_13_reg_we[31:0]),
       .uc2rb_desc_7_xuser_14_reg_we		(uc2rb_desc_7_xuser_14_reg_we[31:0]),
       .uc2rb_desc_7_xuser_15_reg_we		(uc2rb_desc_7_xuser_15_reg_we[31:0]),
       .uc2rb_desc_8_xuser_0_reg_we		(uc2rb_desc_8_xuser_0_reg_we[31:0]),
       .uc2rb_desc_8_xuser_1_reg_we		(uc2rb_desc_8_xuser_1_reg_we[31:0]),
       .uc2rb_desc_8_xuser_2_reg_we		(uc2rb_desc_8_xuser_2_reg_we[31:0]),
       .uc2rb_desc_8_xuser_3_reg_we		(uc2rb_desc_8_xuser_3_reg_we[31:0]),
       .uc2rb_desc_8_xuser_4_reg_we		(uc2rb_desc_8_xuser_4_reg_we[31:0]),
       .uc2rb_desc_8_xuser_5_reg_we		(uc2rb_desc_8_xuser_5_reg_we[31:0]),
       .uc2rb_desc_8_xuser_6_reg_we		(uc2rb_desc_8_xuser_6_reg_we[31:0]),
       .uc2rb_desc_8_xuser_7_reg_we		(uc2rb_desc_8_xuser_7_reg_we[31:0]),
       .uc2rb_desc_8_xuser_8_reg_we		(uc2rb_desc_8_xuser_8_reg_we[31:0]),
       .uc2rb_desc_8_xuser_9_reg_we		(uc2rb_desc_8_xuser_9_reg_we[31:0]),
       .uc2rb_desc_8_xuser_10_reg_we		(uc2rb_desc_8_xuser_10_reg_we[31:0]),
       .uc2rb_desc_8_xuser_11_reg_we		(uc2rb_desc_8_xuser_11_reg_we[31:0]),
       .uc2rb_desc_8_xuser_12_reg_we		(uc2rb_desc_8_xuser_12_reg_we[31:0]),
       .uc2rb_desc_8_xuser_13_reg_we		(uc2rb_desc_8_xuser_13_reg_we[31:0]),
       .uc2rb_desc_8_xuser_14_reg_we		(uc2rb_desc_8_xuser_14_reg_we[31:0]),
       .uc2rb_desc_8_xuser_15_reg_we		(uc2rb_desc_8_xuser_15_reg_we[31:0]),
       .uc2rb_desc_9_xuser_0_reg_we		(uc2rb_desc_9_xuser_0_reg_we[31:0]),
       .uc2rb_desc_9_xuser_1_reg_we		(uc2rb_desc_9_xuser_1_reg_we[31:0]),
       .uc2rb_desc_9_xuser_2_reg_we		(uc2rb_desc_9_xuser_2_reg_we[31:0]),
       .uc2rb_desc_9_xuser_3_reg_we		(uc2rb_desc_9_xuser_3_reg_we[31:0]),
       .uc2rb_desc_9_xuser_4_reg_we		(uc2rb_desc_9_xuser_4_reg_we[31:0]),
       .uc2rb_desc_9_xuser_5_reg_we		(uc2rb_desc_9_xuser_5_reg_we[31:0]),
       .uc2rb_desc_9_xuser_6_reg_we		(uc2rb_desc_9_xuser_6_reg_we[31:0]),
       .uc2rb_desc_9_xuser_7_reg_we		(uc2rb_desc_9_xuser_7_reg_we[31:0]),
       .uc2rb_desc_9_xuser_8_reg_we		(uc2rb_desc_9_xuser_8_reg_we[31:0]),
       .uc2rb_desc_9_xuser_9_reg_we		(uc2rb_desc_9_xuser_9_reg_we[31:0]),
       .uc2rb_desc_9_xuser_10_reg_we		(uc2rb_desc_9_xuser_10_reg_we[31:0]),
       .uc2rb_desc_9_xuser_11_reg_we		(uc2rb_desc_9_xuser_11_reg_we[31:0]),
       .uc2rb_desc_9_xuser_12_reg_we		(uc2rb_desc_9_xuser_12_reg_we[31:0]),
       .uc2rb_desc_9_xuser_13_reg_we		(uc2rb_desc_9_xuser_13_reg_we[31:0]),
       .uc2rb_desc_9_xuser_14_reg_we		(uc2rb_desc_9_xuser_14_reg_we[31:0]),
       .uc2rb_desc_9_xuser_15_reg_we		(uc2rb_desc_9_xuser_15_reg_we[31:0]),
       .uc2rb_desc_10_xuser_0_reg_we		(uc2rb_desc_10_xuser_0_reg_we[31:0]),
       .uc2rb_desc_10_xuser_1_reg_we		(uc2rb_desc_10_xuser_1_reg_we[31:0]),
       .uc2rb_desc_10_xuser_2_reg_we		(uc2rb_desc_10_xuser_2_reg_we[31:0]),
       .uc2rb_desc_10_xuser_3_reg_we		(uc2rb_desc_10_xuser_3_reg_we[31:0]),
       .uc2rb_desc_10_xuser_4_reg_we		(uc2rb_desc_10_xuser_4_reg_we[31:0]),
       .uc2rb_desc_10_xuser_5_reg_we		(uc2rb_desc_10_xuser_5_reg_we[31:0]),
       .uc2rb_desc_10_xuser_6_reg_we		(uc2rb_desc_10_xuser_6_reg_we[31:0]),
       .uc2rb_desc_10_xuser_7_reg_we		(uc2rb_desc_10_xuser_7_reg_we[31:0]),
       .uc2rb_desc_10_xuser_8_reg_we		(uc2rb_desc_10_xuser_8_reg_we[31:0]),
       .uc2rb_desc_10_xuser_9_reg_we		(uc2rb_desc_10_xuser_9_reg_we[31:0]),
       .uc2rb_desc_10_xuser_10_reg_we	(uc2rb_desc_10_xuser_10_reg_we[31:0]),
       .uc2rb_desc_10_xuser_11_reg_we	(uc2rb_desc_10_xuser_11_reg_we[31:0]),
       .uc2rb_desc_10_xuser_12_reg_we	(uc2rb_desc_10_xuser_12_reg_we[31:0]),
       .uc2rb_desc_10_xuser_13_reg_we	(uc2rb_desc_10_xuser_13_reg_we[31:0]),
       .uc2rb_desc_10_xuser_14_reg_we	(uc2rb_desc_10_xuser_14_reg_we[31:0]),
       .uc2rb_desc_10_xuser_15_reg_we	(uc2rb_desc_10_xuser_15_reg_we[31:0]),
       .uc2rb_desc_11_xuser_0_reg_we		(uc2rb_desc_11_xuser_0_reg_we[31:0]),
       .uc2rb_desc_11_xuser_1_reg_we		(uc2rb_desc_11_xuser_1_reg_we[31:0]),
       .uc2rb_desc_11_xuser_2_reg_we		(uc2rb_desc_11_xuser_2_reg_we[31:0]),
       .uc2rb_desc_11_xuser_3_reg_we		(uc2rb_desc_11_xuser_3_reg_we[31:0]),
       .uc2rb_desc_11_xuser_4_reg_we		(uc2rb_desc_11_xuser_4_reg_we[31:0]),
       .uc2rb_desc_11_xuser_5_reg_we		(uc2rb_desc_11_xuser_5_reg_we[31:0]),
       .uc2rb_desc_11_xuser_6_reg_we		(uc2rb_desc_11_xuser_6_reg_we[31:0]),
       .uc2rb_desc_11_xuser_7_reg_we		(uc2rb_desc_11_xuser_7_reg_we[31:0]),
       .uc2rb_desc_11_xuser_8_reg_we		(uc2rb_desc_11_xuser_8_reg_we[31:0]),
       .uc2rb_desc_11_xuser_9_reg_we		(uc2rb_desc_11_xuser_9_reg_we[31:0]),
       .uc2rb_desc_11_xuser_10_reg_we	(uc2rb_desc_11_xuser_10_reg_we[31:0]),
       .uc2rb_desc_11_xuser_11_reg_we	(uc2rb_desc_11_xuser_11_reg_we[31:0]),
       .uc2rb_desc_11_xuser_12_reg_we	(uc2rb_desc_11_xuser_12_reg_we[31:0]),
       .uc2rb_desc_11_xuser_13_reg_we	(uc2rb_desc_11_xuser_13_reg_we[31:0]),
       .uc2rb_desc_11_xuser_14_reg_we	(uc2rb_desc_11_xuser_14_reg_we[31:0]),
       .uc2rb_desc_11_xuser_15_reg_we	(uc2rb_desc_11_xuser_15_reg_we[31:0]),
       .uc2rb_desc_12_xuser_0_reg_we		(uc2rb_desc_12_xuser_0_reg_we[31:0]),
       .uc2rb_desc_12_xuser_1_reg_we		(uc2rb_desc_12_xuser_1_reg_we[31:0]),
       .uc2rb_desc_12_xuser_2_reg_we		(uc2rb_desc_12_xuser_2_reg_we[31:0]),
       .uc2rb_desc_12_xuser_3_reg_we		(uc2rb_desc_12_xuser_3_reg_we[31:0]),
       .uc2rb_desc_12_xuser_4_reg_we		(uc2rb_desc_12_xuser_4_reg_we[31:0]),
       .uc2rb_desc_12_xuser_5_reg_we		(uc2rb_desc_12_xuser_5_reg_we[31:0]),
       .uc2rb_desc_12_xuser_6_reg_we		(uc2rb_desc_12_xuser_6_reg_we[31:0]),
       .uc2rb_desc_12_xuser_7_reg_we		(uc2rb_desc_12_xuser_7_reg_we[31:0]),
       .uc2rb_desc_12_xuser_8_reg_we		(uc2rb_desc_12_xuser_8_reg_we[31:0]),
       .uc2rb_desc_12_xuser_9_reg_we		(uc2rb_desc_12_xuser_9_reg_we[31:0]),
       .uc2rb_desc_12_xuser_10_reg_we	(uc2rb_desc_12_xuser_10_reg_we[31:0]),
       .uc2rb_desc_12_xuser_11_reg_we	(uc2rb_desc_12_xuser_11_reg_we[31:0]),
       .uc2rb_desc_12_xuser_12_reg_we	(uc2rb_desc_12_xuser_12_reg_we[31:0]),
       .uc2rb_desc_12_xuser_13_reg_we	(uc2rb_desc_12_xuser_13_reg_we[31:0]),
       .uc2rb_desc_12_xuser_14_reg_we	(uc2rb_desc_12_xuser_14_reg_we[31:0]),
       .uc2rb_desc_12_xuser_15_reg_we	(uc2rb_desc_12_xuser_15_reg_we[31:0]),
       .uc2rb_desc_13_xuser_0_reg_we		(uc2rb_desc_13_xuser_0_reg_we[31:0]),
       .uc2rb_desc_13_xuser_1_reg_we		(uc2rb_desc_13_xuser_1_reg_we[31:0]),
       .uc2rb_desc_13_xuser_2_reg_we		(uc2rb_desc_13_xuser_2_reg_we[31:0]),
       .uc2rb_desc_13_xuser_3_reg_we		(uc2rb_desc_13_xuser_3_reg_we[31:0]),
       .uc2rb_desc_13_xuser_4_reg_we		(uc2rb_desc_13_xuser_4_reg_we[31:0]),
       .uc2rb_desc_13_xuser_5_reg_we		(uc2rb_desc_13_xuser_5_reg_we[31:0]),
       .uc2rb_desc_13_xuser_6_reg_we		(uc2rb_desc_13_xuser_6_reg_we[31:0]),
       .uc2rb_desc_13_xuser_7_reg_we		(uc2rb_desc_13_xuser_7_reg_we[31:0]),
       .uc2rb_desc_13_xuser_8_reg_we		(uc2rb_desc_13_xuser_8_reg_we[31:0]),
       .uc2rb_desc_13_xuser_9_reg_we		(uc2rb_desc_13_xuser_9_reg_we[31:0]),
       .uc2rb_desc_13_xuser_10_reg_we	(uc2rb_desc_13_xuser_10_reg_we[31:0]),
       .uc2rb_desc_13_xuser_11_reg_we	(uc2rb_desc_13_xuser_11_reg_we[31:0]),
       .uc2rb_desc_13_xuser_12_reg_we	(uc2rb_desc_13_xuser_12_reg_we[31:0]),
       .uc2rb_desc_13_xuser_13_reg_we	(uc2rb_desc_13_xuser_13_reg_we[31:0]),
       .uc2rb_desc_13_xuser_14_reg_we	(uc2rb_desc_13_xuser_14_reg_we[31:0]),
       .uc2rb_desc_13_xuser_15_reg_we	(uc2rb_desc_13_xuser_15_reg_we[31:0]),
       .uc2rb_desc_14_xuser_0_reg_we		(uc2rb_desc_14_xuser_0_reg_we[31:0]),
       .uc2rb_desc_14_xuser_1_reg_we		(uc2rb_desc_14_xuser_1_reg_we[31:0]),
       .uc2rb_desc_14_xuser_2_reg_we		(uc2rb_desc_14_xuser_2_reg_we[31:0]),
       .uc2rb_desc_14_xuser_3_reg_we		(uc2rb_desc_14_xuser_3_reg_we[31:0]),
       .uc2rb_desc_14_xuser_4_reg_we		(uc2rb_desc_14_xuser_4_reg_we[31:0]),
       .uc2rb_desc_14_xuser_5_reg_we		(uc2rb_desc_14_xuser_5_reg_we[31:0]),
       .uc2rb_desc_14_xuser_6_reg_we		(uc2rb_desc_14_xuser_6_reg_we[31:0]),
       .uc2rb_desc_14_xuser_7_reg_we		(uc2rb_desc_14_xuser_7_reg_we[31:0]),
       .uc2rb_desc_14_xuser_8_reg_we		(uc2rb_desc_14_xuser_8_reg_we[31:0]),
       .uc2rb_desc_14_xuser_9_reg_we		(uc2rb_desc_14_xuser_9_reg_we[31:0]),
       .uc2rb_desc_14_xuser_10_reg_we	(uc2rb_desc_14_xuser_10_reg_we[31:0]),
       .uc2rb_desc_14_xuser_11_reg_we	(uc2rb_desc_14_xuser_11_reg_we[31:0]),
       .uc2rb_desc_14_xuser_12_reg_we	(uc2rb_desc_14_xuser_12_reg_we[31:0]),
       .uc2rb_desc_14_xuser_13_reg_we	(uc2rb_desc_14_xuser_13_reg_we[31:0]),
       .uc2rb_desc_14_xuser_14_reg_we	(uc2rb_desc_14_xuser_14_reg_we[31:0]),
       .uc2rb_desc_14_xuser_15_reg_we	(uc2rb_desc_14_xuser_15_reg_we[31:0]),
       .uc2rb_desc_15_xuser_0_reg_we		(uc2rb_desc_15_xuser_0_reg_we[31:0]),
       .uc2rb_desc_15_xuser_1_reg_we		(uc2rb_desc_15_xuser_1_reg_we[31:0]),
       .uc2rb_desc_15_xuser_2_reg_we		(uc2rb_desc_15_xuser_2_reg_we[31:0]),
       .uc2rb_desc_15_xuser_3_reg_we		(uc2rb_desc_15_xuser_3_reg_we[31:0]),
       .uc2rb_desc_15_xuser_4_reg_we		(uc2rb_desc_15_xuser_4_reg_we[31:0]),
       .uc2rb_desc_15_xuser_5_reg_we		(uc2rb_desc_15_xuser_5_reg_we[31:0]),
       .uc2rb_desc_15_xuser_6_reg_we		(uc2rb_desc_15_xuser_6_reg_we[31:0]),
       .uc2rb_desc_15_xuser_7_reg_we		(uc2rb_desc_15_xuser_7_reg_we[31:0]),
       .uc2rb_desc_15_xuser_8_reg_we		(uc2rb_desc_15_xuser_8_reg_we[31:0]),
       .uc2rb_desc_15_xuser_9_reg_we		(uc2rb_desc_15_xuser_9_reg_we[31:0]),
       .uc2rb_desc_15_xuser_10_reg_we	(uc2rb_desc_15_xuser_10_reg_we[31:0]),
       .uc2rb_desc_15_xuser_11_reg_we	(uc2rb_desc_15_xuser_11_reg_we[31:0]),
       .uc2rb_desc_15_xuser_12_reg_we	(uc2rb_desc_15_xuser_12_reg_we[31:0]),
       .uc2rb_desc_15_xuser_13_reg_we	(uc2rb_desc_15_xuser_13_reg_we[31:0]),
       .uc2rb_desc_15_xuser_14_reg_we	(uc2rb_desc_15_xuser_14_reg_we[31:0]),
       .uc2rb_desc_15_xuser_15_reg_we	(uc2rb_desc_15_xuser_15_reg_we[31:0]),
       .m_axi_usr_awid					(m_axi_usr_awid[M_AXI_USR_ID_WIDTH-1:0]),
       .m_axi_usr_awaddr					(m_axi_usr_awaddr[M_AXI_USR_ADDR_WIDTH-1:0]),
       .m_axi_usr_awlen					(m_axi_usr_awlen[M_AXI_USR_LEN_WIDTH-1:0]),
       .m_axi_usr_awsize					(m_axi_usr_awsize[2:0]),
       .m_axi_usr_awburst				(m_axi_usr_awburst[1:0]),
       .m_axi_usr_awlock					(m_axi_usr_awlock),
       .m_axi_usr_awcache				(m_axi_usr_awcache[3:0]),
       .m_axi_usr_awprot					(m_axi_usr_awprot[2:0]),
       .m_axi_usr_awqos					(m_axi_usr_awqos[3:0]),
       .m_axi_usr_awregion				(m_axi_usr_awregion[3:0]),
       .m_axi_usr_awuser					(m_axi_usr_awuser ),
       .m_axi_usr_awvalid				(m_axi_usr_awvalid),
       .m_axi_usr_wdata					(m_axi_usr_wdata[M_AXI_USR_DATA_WIDTH-1:0]),
       .m_axi_usr_wstrb					(m_axi_usr_wstrb[(M_AXI_USR_DATA_WIDTH/8)-1:0]),
       .m_axi_usr_wlast					(m_axi_usr_wlast),
       .m_axi_usr_wuser					(m_axi_usr_wuser ),
       .m_axi_usr_wvalid					(m_axi_usr_wvalid),
       .m_axi_usr_bready					(m_axi_usr_bready),
       .m_axi_usr_arid					(m_axi_usr_arid[M_AXI_USR_ID_WIDTH-1:0]),
       .m_axi_usr_araddr					(m_axi_usr_araddr[M_AXI_USR_ADDR_WIDTH-1:0]),
       .m_axi_usr_arlen					(m_axi_usr_arlen[M_AXI_USR_LEN_WIDTH-1:0]),
       .m_axi_usr_arsize					(m_axi_usr_arsize[2:0]),
       .m_axi_usr_arburst				(m_axi_usr_arburst[1:0]),
       .m_axi_usr_arlock					(m_axi_usr_arlock),
       .m_axi_usr_arcache				(m_axi_usr_arcache[3:0]),
       .m_axi_usr_arprot					(m_axi_usr_arprot[2:0]),
       .m_axi_usr_arqos					(m_axi_usr_arqos[3:0]),
       .m_axi_usr_arregion				(m_axi_usr_arregion[3:0]),
       .m_axi_usr_aruser					(m_axi_usr_aruser ),
       .m_axi_usr_arvalid				(m_axi_usr_arvalid),
       .m_axi_usr_rready					(m_axi_usr_rready),
       .m_axi_usr_wid					(m_axi_usr_wid[M_AXI_USR_ID_WIDTH-1:0]),
       // Inputs
       .axi_aclk							(axi_aclk),
       .axi_aresetn						(axi_aresetn),
       .rb2uc_rd_data					(rb2uc_rd_data[M_AXI_USR_DATA_WIDTH-1:0]),
       .rb2uc_rd_wstrb					(rb2uc_rd_wstrb[(M_AXI_USR_DATA_WIDTH/8-1):0]),
       .hm2uc_done						(hm2uc_done[15:0]),
       .version_reg						(version_reg[31:0]),
       .bridge_type_reg					(bridge_type_reg[31:0]),
       .mode_select_reg					(mode_select_reg[31:0]),
       .reset_reg						(reset_reg[31:0]),
       .intr_h2c_0_reg					(intr_h2c_0_reg[31:0]),
       .intr_h2c_1_reg					(intr_h2c_1_reg[31:0]),
       .intr_c2h_0_status_reg			(intr_c2h_0_status_reg[31:0]),
       .intr_c2h_1_status_reg			(intr_c2h_1_status_reg[31:0]),
       .c2h_gpio_0_status_reg			(c2h_gpio_0_status_reg[31:0]),
       .c2h_gpio_1_status_reg			(c2h_gpio_1_status_reg[31:0]),
       .c2h_gpio_2_status_reg			(c2h_gpio_2_status_reg[31:0]),
       .c2h_gpio_3_status_reg			(c2h_gpio_3_status_reg[31:0]),
       .c2h_gpio_4_status_reg			(c2h_gpio_4_status_reg[31:0]),
       .c2h_gpio_5_status_reg			(c2h_gpio_5_status_reg[31:0]),
       .c2h_gpio_6_status_reg			(c2h_gpio_6_status_reg[31:0]),
       .c2h_gpio_7_status_reg			(c2h_gpio_7_status_reg[31:0]),
       .c2h_gpio_8_status_reg			(c2h_gpio_8_status_reg[31:0]),
       .c2h_gpio_9_status_reg			(c2h_gpio_9_status_reg[31:0]),
       .c2h_gpio_10_status_reg			(c2h_gpio_10_status_reg[31:0]),
       .c2h_gpio_11_status_reg			(c2h_gpio_11_status_reg[31:0]),
       .c2h_gpio_12_status_reg			(c2h_gpio_12_status_reg[31:0]),
       .c2h_gpio_13_status_reg			(c2h_gpio_13_status_reg[31:0]),
       .c2h_gpio_14_status_reg			(c2h_gpio_14_status_reg[31:0]),
       .c2h_gpio_15_status_reg			(c2h_gpio_15_status_reg[31:0]),
       .axi_bridge_config_reg			(axi_bridge_config_reg[31:0]),
       .axi_max_desc_reg					(axi_max_desc_reg[31:0]),
       .intr_status_reg					(intr_status_reg[31:0]),
       .intr_error_status_reg			(intr_error_status_reg[31:0]),
       .intr_error_clear_reg				(intr_error_clear_reg[31:0]),
       .intr_error_enable_reg			(intr_error_enable_reg[31:0]),
       .ownership_reg					(ownership_reg[31:0]),
       .ownership_flip_reg				(ownership_flip_reg[31:0]),
       .status_resp_reg					(status_resp_reg[31:0]),
       .intr_comp_status_reg				(intr_comp_status_reg[31:0]),
       .intr_comp_clear_reg				(intr_comp_clear_reg[31:0]),
       .intr_comp_enable_reg				(intr_comp_enable_reg[31:0]),
       .desc_0_txn_type_reg				(desc_0_txn_type_reg[31:0]),
       .desc_0_size_reg					(desc_0_size_reg[31:0]),
       .desc_0_data_offset_reg			(desc_0_data_offset_reg[31:0]),
       .desc_0_data_host_addr_0_reg		(desc_0_data_host_addr_0_reg[31:0]),
       .desc_0_data_host_addr_1_reg		(desc_0_data_host_addr_1_reg[31:0]),
       .desc_0_data_host_addr_2_reg		(desc_0_data_host_addr_2_reg[31:0]),
       .desc_0_data_host_addr_3_reg		(desc_0_data_host_addr_3_reg[31:0]),
       .desc_0_wstrb_host_addr_0_reg		(desc_0_wstrb_host_addr_0_reg[31:0]),
       .desc_0_wstrb_host_addr_1_reg		(desc_0_wstrb_host_addr_1_reg[31:0]),
       .desc_0_wstrb_host_addr_2_reg		(desc_0_wstrb_host_addr_2_reg[31:0]),
       .desc_0_wstrb_host_addr_3_reg		(desc_0_wstrb_host_addr_3_reg[31:0]),
       .desc_0_axsize_reg				(desc_0_axsize_reg[31:0]),
       .desc_0_attr_reg					(desc_0_attr_reg[31:0]),
       .desc_0_axaddr_0_reg				(desc_0_axaddr_0_reg[31:0]),
       .desc_0_axaddr_1_reg				(desc_0_axaddr_1_reg[31:0]),
       .desc_0_axaddr_2_reg				(desc_0_axaddr_2_reg[31:0]),
       .desc_0_axaddr_3_reg				(desc_0_axaddr_3_reg[31:0]),
       .desc_0_axid_0_reg				(desc_0_axid_0_reg[31:0]),
       .desc_0_axid_1_reg				(desc_0_axid_1_reg[31:0]),
       .desc_0_axid_2_reg				(desc_0_axid_2_reg[31:0]),
       .desc_0_axid_3_reg				(desc_0_axid_3_reg[31:0]),
       .desc_0_axuser_0_reg				(desc_0_axuser_0_reg[31:0]),
       .desc_0_axuser_1_reg				(desc_0_axuser_1_reg[31:0]),
       .desc_0_axuser_2_reg				(desc_0_axuser_2_reg[31:0]),
       .desc_0_axuser_3_reg				(desc_0_axuser_3_reg[31:0]),
       .desc_0_axuser_4_reg				(desc_0_axuser_4_reg[31:0]),
       .desc_0_axuser_5_reg				(desc_0_axuser_5_reg[31:0]),
       .desc_0_axuser_6_reg				(desc_0_axuser_6_reg[31:0]),
       .desc_0_axuser_7_reg				(desc_0_axuser_7_reg[31:0]),
       .desc_0_axuser_8_reg				(desc_0_axuser_8_reg[31:0]),
       .desc_0_axuser_9_reg				(desc_0_axuser_9_reg[31:0]),
       .desc_0_axuser_10_reg				(desc_0_axuser_10_reg[31:0]),
       .desc_0_axuser_11_reg				(desc_0_axuser_11_reg[31:0]),
       .desc_0_axuser_12_reg				(desc_0_axuser_12_reg[31:0]),
       .desc_0_axuser_13_reg				(desc_0_axuser_13_reg[31:0]),
       .desc_0_axuser_14_reg				(desc_0_axuser_14_reg[31:0]),
       .desc_0_axuser_15_reg				(desc_0_axuser_15_reg[31:0]),
       .desc_0_xuser_0_reg				(desc_0_xuser_0_reg[31:0]),
       .desc_0_xuser_1_reg				(desc_0_xuser_1_reg[31:0]),
       .desc_0_xuser_2_reg				(desc_0_xuser_2_reg[31:0]),
       .desc_0_xuser_3_reg				(desc_0_xuser_3_reg[31:0]),
       .desc_0_xuser_4_reg				(desc_0_xuser_4_reg[31:0]),
       .desc_0_xuser_5_reg				(desc_0_xuser_5_reg[31:0]),
       .desc_0_xuser_6_reg				(desc_0_xuser_6_reg[31:0]),
       .desc_0_xuser_7_reg				(desc_0_xuser_7_reg[31:0]),
       .desc_0_xuser_8_reg				(desc_0_xuser_8_reg[31:0]),
       .desc_0_xuser_9_reg				(desc_0_xuser_9_reg[31:0]),
       .desc_0_xuser_10_reg				(desc_0_xuser_10_reg[31:0]),
       .desc_0_xuser_11_reg				(desc_0_xuser_11_reg[31:0]),
       .desc_0_xuser_12_reg				(desc_0_xuser_12_reg[31:0]),
       .desc_0_xuser_13_reg				(desc_0_xuser_13_reg[31:0]),
       .desc_0_xuser_14_reg				(desc_0_xuser_14_reg[31:0]),
       .desc_0_xuser_15_reg				(desc_0_xuser_15_reg[31:0]),
       .desc_0_wuser_0_reg				(desc_0_wuser_0_reg[31:0]),
       .desc_0_wuser_1_reg				(desc_0_wuser_1_reg[31:0]),
       .desc_0_wuser_2_reg				(desc_0_wuser_2_reg[31:0]),
       .desc_0_wuser_3_reg				(desc_0_wuser_3_reg[31:0]),
       .desc_0_wuser_4_reg				(desc_0_wuser_4_reg[31:0]),
       .desc_0_wuser_5_reg				(desc_0_wuser_5_reg[31:0]),
       .desc_0_wuser_6_reg				(desc_0_wuser_6_reg[31:0]),
       .desc_0_wuser_7_reg				(desc_0_wuser_7_reg[31:0]),
       .desc_0_wuser_8_reg				(desc_0_wuser_8_reg[31:0]),
       .desc_0_wuser_9_reg				(desc_0_wuser_9_reg[31:0]),
       .desc_0_wuser_10_reg				(desc_0_wuser_10_reg[31:0]),
       .desc_0_wuser_11_reg				(desc_0_wuser_11_reg[31:0]),
       .desc_0_wuser_12_reg				(desc_0_wuser_12_reg[31:0]),
       .desc_0_wuser_13_reg				(desc_0_wuser_13_reg[31:0]),
       .desc_0_wuser_14_reg				(desc_0_wuser_14_reg[31:0]),
       .desc_0_wuser_15_reg				(desc_0_wuser_15_reg[31:0]),
       .desc_1_txn_type_reg				(desc_1_txn_type_reg[31:0]),
       .desc_1_size_reg					(desc_1_size_reg[31:0]),
       .desc_1_data_offset_reg			(desc_1_data_offset_reg[31:0]),
       .desc_1_data_host_addr_0_reg		(desc_1_data_host_addr_0_reg[31:0]),
       .desc_1_data_host_addr_1_reg		(desc_1_data_host_addr_1_reg[31:0]),
       .desc_1_data_host_addr_2_reg		(desc_1_data_host_addr_2_reg[31:0]),
       .desc_1_data_host_addr_3_reg		(desc_1_data_host_addr_3_reg[31:0]),
       .desc_1_wstrb_host_addr_0_reg		(desc_1_wstrb_host_addr_0_reg[31:0]),
       .desc_1_wstrb_host_addr_1_reg		(desc_1_wstrb_host_addr_1_reg[31:0]),
       .desc_1_wstrb_host_addr_2_reg		(desc_1_wstrb_host_addr_2_reg[31:0]),
       .desc_1_wstrb_host_addr_3_reg		(desc_1_wstrb_host_addr_3_reg[31:0]),
       .desc_1_axsize_reg				(desc_1_axsize_reg[31:0]),
       .desc_1_attr_reg					(desc_1_attr_reg[31:0]),
       .desc_1_axaddr_0_reg				(desc_1_axaddr_0_reg[31:0]),
       .desc_1_axaddr_1_reg				(desc_1_axaddr_1_reg[31:0]),
       .desc_1_axaddr_2_reg				(desc_1_axaddr_2_reg[31:0]),
       .desc_1_axaddr_3_reg				(desc_1_axaddr_3_reg[31:0]),
       .desc_1_axid_0_reg				(desc_1_axid_0_reg[31:0]),
       .desc_1_axid_1_reg				(desc_1_axid_1_reg[31:0]),
       .desc_1_axid_2_reg				(desc_1_axid_2_reg[31:0]),
       .desc_1_axid_3_reg				(desc_1_axid_3_reg[31:0]),
       .desc_1_axuser_0_reg				(desc_1_axuser_0_reg[31:0]),
       .desc_1_axuser_1_reg				(desc_1_axuser_1_reg[31:0]),
       .desc_1_axuser_2_reg				(desc_1_axuser_2_reg[31:0]),
       .desc_1_axuser_3_reg				(desc_1_axuser_3_reg[31:0]),
       .desc_1_axuser_4_reg				(desc_1_axuser_4_reg[31:0]),
       .desc_1_axuser_5_reg				(desc_1_axuser_5_reg[31:0]),
       .desc_1_axuser_6_reg				(desc_1_axuser_6_reg[31:0]),
       .desc_1_axuser_7_reg				(desc_1_axuser_7_reg[31:0]),
       .desc_1_axuser_8_reg				(desc_1_axuser_8_reg[31:0]),
       .desc_1_axuser_9_reg				(desc_1_axuser_9_reg[31:0]),
       .desc_1_axuser_10_reg				(desc_1_axuser_10_reg[31:0]),
       .desc_1_axuser_11_reg				(desc_1_axuser_11_reg[31:0]),
       .desc_1_axuser_12_reg				(desc_1_axuser_12_reg[31:0]),
       .desc_1_axuser_13_reg				(desc_1_axuser_13_reg[31:0]),
       .desc_1_axuser_14_reg				(desc_1_axuser_14_reg[31:0]),
       .desc_1_axuser_15_reg				(desc_1_axuser_15_reg[31:0]),
       .desc_1_xuser_0_reg				(desc_1_xuser_0_reg[31:0]),
       .desc_1_xuser_1_reg				(desc_1_xuser_1_reg[31:0]),
       .desc_1_xuser_2_reg				(desc_1_xuser_2_reg[31:0]),
       .desc_1_xuser_3_reg				(desc_1_xuser_3_reg[31:0]),
       .desc_1_xuser_4_reg				(desc_1_xuser_4_reg[31:0]),
       .desc_1_xuser_5_reg				(desc_1_xuser_5_reg[31:0]),
       .desc_1_xuser_6_reg				(desc_1_xuser_6_reg[31:0]),
       .desc_1_xuser_7_reg				(desc_1_xuser_7_reg[31:0]),
       .desc_1_xuser_8_reg				(desc_1_xuser_8_reg[31:0]),
       .desc_1_xuser_9_reg				(desc_1_xuser_9_reg[31:0]),
       .desc_1_xuser_10_reg				(desc_1_xuser_10_reg[31:0]),
       .desc_1_xuser_11_reg				(desc_1_xuser_11_reg[31:0]),
       .desc_1_xuser_12_reg				(desc_1_xuser_12_reg[31:0]),
       .desc_1_xuser_13_reg				(desc_1_xuser_13_reg[31:0]),
       .desc_1_xuser_14_reg				(desc_1_xuser_14_reg[31:0]),
       .desc_1_xuser_15_reg				(desc_1_xuser_15_reg[31:0]),
       .desc_1_wuser_0_reg				(desc_1_wuser_0_reg[31:0]),
       .desc_1_wuser_1_reg				(desc_1_wuser_1_reg[31:0]),
       .desc_1_wuser_2_reg				(desc_1_wuser_2_reg[31:0]),
       .desc_1_wuser_3_reg				(desc_1_wuser_3_reg[31:0]),
       .desc_1_wuser_4_reg				(desc_1_wuser_4_reg[31:0]),
       .desc_1_wuser_5_reg				(desc_1_wuser_5_reg[31:0]),
       .desc_1_wuser_6_reg				(desc_1_wuser_6_reg[31:0]),
       .desc_1_wuser_7_reg				(desc_1_wuser_7_reg[31:0]),
       .desc_1_wuser_8_reg				(desc_1_wuser_8_reg[31:0]),
       .desc_1_wuser_9_reg				(desc_1_wuser_9_reg[31:0]),
       .desc_1_wuser_10_reg				(desc_1_wuser_10_reg[31:0]),
       .desc_1_wuser_11_reg				(desc_1_wuser_11_reg[31:0]),
       .desc_1_wuser_12_reg				(desc_1_wuser_12_reg[31:0]),
       .desc_1_wuser_13_reg				(desc_1_wuser_13_reg[31:0]),
       .desc_1_wuser_14_reg				(desc_1_wuser_14_reg[31:0]),
       .desc_1_wuser_15_reg				(desc_1_wuser_15_reg[31:0]),
       .desc_2_txn_type_reg				(desc_2_txn_type_reg[31:0]),
       .desc_2_size_reg					(desc_2_size_reg[31:0]),
       .desc_2_data_offset_reg			(desc_2_data_offset_reg[31:0]),
       .desc_2_data_host_addr_0_reg		(desc_2_data_host_addr_0_reg[31:0]),
       .desc_2_data_host_addr_1_reg		(desc_2_data_host_addr_1_reg[31:0]),
       .desc_2_data_host_addr_2_reg		(desc_2_data_host_addr_2_reg[31:0]),
       .desc_2_data_host_addr_3_reg		(desc_2_data_host_addr_3_reg[31:0]),
       .desc_2_wstrb_host_addr_0_reg		(desc_2_wstrb_host_addr_0_reg[31:0]),
       .desc_2_wstrb_host_addr_1_reg		(desc_2_wstrb_host_addr_1_reg[31:0]),
       .desc_2_wstrb_host_addr_2_reg		(desc_2_wstrb_host_addr_2_reg[31:0]),
       .desc_2_wstrb_host_addr_3_reg		(desc_2_wstrb_host_addr_3_reg[31:0]),
       .desc_2_axsize_reg				(desc_2_axsize_reg[31:0]),
       .desc_2_attr_reg					(desc_2_attr_reg[31:0]),
       .desc_2_axaddr_0_reg				(desc_2_axaddr_0_reg[31:0]),
       .desc_2_axaddr_1_reg				(desc_2_axaddr_1_reg[31:0]),
       .desc_2_axaddr_2_reg				(desc_2_axaddr_2_reg[31:0]),
       .desc_2_axaddr_3_reg				(desc_2_axaddr_3_reg[31:0]),
       .desc_2_axid_0_reg				(desc_2_axid_0_reg[31:0]),
       .desc_2_axid_1_reg				(desc_2_axid_1_reg[31:0]),
       .desc_2_axid_2_reg				(desc_2_axid_2_reg[31:0]),
       .desc_2_axid_3_reg				(desc_2_axid_3_reg[31:0]),
       .desc_2_axuser_0_reg				(desc_2_axuser_0_reg[31:0]),
       .desc_2_axuser_1_reg				(desc_2_axuser_1_reg[31:0]),
       .desc_2_axuser_2_reg				(desc_2_axuser_2_reg[31:0]),
       .desc_2_axuser_3_reg				(desc_2_axuser_3_reg[31:0]),
       .desc_2_axuser_4_reg				(desc_2_axuser_4_reg[31:0]),
       .desc_2_axuser_5_reg				(desc_2_axuser_5_reg[31:0]),
       .desc_2_axuser_6_reg				(desc_2_axuser_6_reg[31:0]),
       .desc_2_axuser_7_reg				(desc_2_axuser_7_reg[31:0]),
       .desc_2_axuser_8_reg				(desc_2_axuser_8_reg[31:0]),
       .desc_2_axuser_9_reg				(desc_2_axuser_9_reg[31:0]),
       .desc_2_axuser_10_reg				(desc_2_axuser_10_reg[31:0]),
       .desc_2_axuser_11_reg				(desc_2_axuser_11_reg[31:0]),
       .desc_2_axuser_12_reg				(desc_2_axuser_12_reg[31:0]),
       .desc_2_axuser_13_reg				(desc_2_axuser_13_reg[31:0]),
       .desc_2_axuser_14_reg				(desc_2_axuser_14_reg[31:0]),
       .desc_2_axuser_15_reg				(desc_2_axuser_15_reg[31:0]),
       .desc_2_xuser_0_reg				(desc_2_xuser_0_reg[31:0]),
       .desc_2_xuser_1_reg				(desc_2_xuser_1_reg[31:0]),
       .desc_2_xuser_2_reg				(desc_2_xuser_2_reg[31:0]),
       .desc_2_xuser_3_reg				(desc_2_xuser_3_reg[31:0]),
       .desc_2_xuser_4_reg				(desc_2_xuser_4_reg[31:0]),
       .desc_2_xuser_5_reg				(desc_2_xuser_5_reg[31:0]),
       .desc_2_xuser_6_reg				(desc_2_xuser_6_reg[31:0]),
       .desc_2_xuser_7_reg				(desc_2_xuser_7_reg[31:0]),
       .desc_2_xuser_8_reg				(desc_2_xuser_8_reg[31:0]),
       .desc_2_xuser_9_reg				(desc_2_xuser_9_reg[31:0]),
       .desc_2_xuser_10_reg				(desc_2_xuser_10_reg[31:0]),
       .desc_2_xuser_11_reg				(desc_2_xuser_11_reg[31:0]),
       .desc_2_xuser_12_reg				(desc_2_xuser_12_reg[31:0]),
       .desc_2_xuser_13_reg				(desc_2_xuser_13_reg[31:0]),
       .desc_2_xuser_14_reg				(desc_2_xuser_14_reg[31:0]),
       .desc_2_xuser_15_reg				(desc_2_xuser_15_reg[31:0]),
       .desc_2_wuser_0_reg				(desc_2_wuser_0_reg[31:0]),
       .desc_2_wuser_1_reg				(desc_2_wuser_1_reg[31:0]),
       .desc_2_wuser_2_reg				(desc_2_wuser_2_reg[31:0]),
       .desc_2_wuser_3_reg				(desc_2_wuser_3_reg[31:0]),
       .desc_2_wuser_4_reg				(desc_2_wuser_4_reg[31:0]),
       .desc_2_wuser_5_reg				(desc_2_wuser_5_reg[31:0]),
       .desc_2_wuser_6_reg				(desc_2_wuser_6_reg[31:0]),
       .desc_2_wuser_7_reg				(desc_2_wuser_7_reg[31:0]),
       .desc_2_wuser_8_reg				(desc_2_wuser_8_reg[31:0]),
       .desc_2_wuser_9_reg				(desc_2_wuser_9_reg[31:0]),
       .desc_2_wuser_10_reg				(desc_2_wuser_10_reg[31:0]),
       .desc_2_wuser_11_reg				(desc_2_wuser_11_reg[31:0]),
       .desc_2_wuser_12_reg				(desc_2_wuser_12_reg[31:0]),
       .desc_2_wuser_13_reg				(desc_2_wuser_13_reg[31:0]),
       .desc_2_wuser_14_reg				(desc_2_wuser_14_reg[31:0]),
       .desc_2_wuser_15_reg				(desc_2_wuser_15_reg[31:0]),
       .desc_3_txn_type_reg				(desc_3_txn_type_reg[31:0]),
       .desc_3_size_reg					(desc_3_size_reg[31:0]),
       .desc_3_data_offset_reg			(desc_3_data_offset_reg[31:0]),
       .desc_3_data_host_addr_0_reg		(desc_3_data_host_addr_0_reg[31:0]),
       .desc_3_data_host_addr_1_reg		(desc_3_data_host_addr_1_reg[31:0]),
       .desc_3_data_host_addr_2_reg		(desc_3_data_host_addr_2_reg[31:0]),
       .desc_3_data_host_addr_3_reg		(desc_3_data_host_addr_3_reg[31:0]),
       .desc_3_wstrb_host_addr_0_reg		(desc_3_wstrb_host_addr_0_reg[31:0]),
       .desc_3_wstrb_host_addr_1_reg		(desc_3_wstrb_host_addr_1_reg[31:0]),
       .desc_3_wstrb_host_addr_2_reg		(desc_3_wstrb_host_addr_2_reg[31:0]),
       .desc_3_wstrb_host_addr_3_reg		(desc_3_wstrb_host_addr_3_reg[31:0]),
       .desc_3_axsize_reg				(desc_3_axsize_reg[31:0]),
       .desc_3_attr_reg					(desc_3_attr_reg[31:0]),
       .desc_3_axaddr_0_reg				(desc_3_axaddr_0_reg[31:0]),
       .desc_3_axaddr_1_reg				(desc_3_axaddr_1_reg[31:0]),
       .desc_3_axaddr_2_reg				(desc_3_axaddr_2_reg[31:0]),
       .desc_3_axaddr_3_reg				(desc_3_axaddr_3_reg[31:0]),
       .desc_3_axid_0_reg				(desc_3_axid_0_reg[31:0]),
       .desc_3_axid_1_reg				(desc_3_axid_1_reg[31:0]),
       .desc_3_axid_2_reg				(desc_3_axid_2_reg[31:0]),
       .desc_3_axid_3_reg				(desc_3_axid_3_reg[31:0]),
       .desc_3_axuser_0_reg				(desc_3_axuser_0_reg[31:0]),
       .desc_3_axuser_1_reg				(desc_3_axuser_1_reg[31:0]),
       .desc_3_axuser_2_reg				(desc_3_axuser_2_reg[31:0]),
       .desc_3_axuser_3_reg				(desc_3_axuser_3_reg[31:0]),
       .desc_3_axuser_4_reg				(desc_3_axuser_4_reg[31:0]),
       .desc_3_axuser_5_reg				(desc_3_axuser_5_reg[31:0]),
       .desc_3_axuser_6_reg				(desc_3_axuser_6_reg[31:0]),
       .desc_3_axuser_7_reg				(desc_3_axuser_7_reg[31:0]),
       .desc_3_axuser_8_reg				(desc_3_axuser_8_reg[31:0]),
       .desc_3_axuser_9_reg				(desc_3_axuser_9_reg[31:0]),
       .desc_3_axuser_10_reg				(desc_3_axuser_10_reg[31:0]),
       .desc_3_axuser_11_reg				(desc_3_axuser_11_reg[31:0]),
       .desc_3_axuser_12_reg				(desc_3_axuser_12_reg[31:0]),
       .desc_3_axuser_13_reg				(desc_3_axuser_13_reg[31:0]),
       .desc_3_axuser_14_reg				(desc_3_axuser_14_reg[31:0]),
       .desc_3_axuser_15_reg				(desc_3_axuser_15_reg[31:0]),
       .desc_3_xuser_0_reg				(desc_3_xuser_0_reg[31:0]),
       .desc_3_xuser_1_reg				(desc_3_xuser_1_reg[31:0]),
       .desc_3_xuser_2_reg				(desc_3_xuser_2_reg[31:0]),
       .desc_3_xuser_3_reg				(desc_3_xuser_3_reg[31:0]),
       .desc_3_xuser_4_reg				(desc_3_xuser_4_reg[31:0]),
       .desc_3_xuser_5_reg				(desc_3_xuser_5_reg[31:0]),
       .desc_3_xuser_6_reg				(desc_3_xuser_6_reg[31:0]),
       .desc_3_xuser_7_reg				(desc_3_xuser_7_reg[31:0]),
       .desc_3_xuser_8_reg				(desc_3_xuser_8_reg[31:0]),
       .desc_3_xuser_9_reg				(desc_3_xuser_9_reg[31:0]),
       .desc_3_xuser_10_reg				(desc_3_xuser_10_reg[31:0]),
       .desc_3_xuser_11_reg				(desc_3_xuser_11_reg[31:0]),
       .desc_3_xuser_12_reg				(desc_3_xuser_12_reg[31:0]),
       .desc_3_xuser_13_reg				(desc_3_xuser_13_reg[31:0]),
       .desc_3_xuser_14_reg				(desc_3_xuser_14_reg[31:0]),
       .desc_3_xuser_15_reg				(desc_3_xuser_15_reg[31:0]),
       .desc_3_wuser_0_reg				(desc_3_wuser_0_reg[31:0]),
       .desc_3_wuser_1_reg				(desc_3_wuser_1_reg[31:0]),
       .desc_3_wuser_2_reg				(desc_3_wuser_2_reg[31:0]),
       .desc_3_wuser_3_reg				(desc_3_wuser_3_reg[31:0]),
       .desc_3_wuser_4_reg				(desc_3_wuser_4_reg[31:0]),
       .desc_3_wuser_5_reg				(desc_3_wuser_5_reg[31:0]),
       .desc_3_wuser_6_reg				(desc_3_wuser_6_reg[31:0]),
       .desc_3_wuser_7_reg				(desc_3_wuser_7_reg[31:0]),
       .desc_3_wuser_8_reg				(desc_3_wuser_8_reg[31:0]),
       .desc_3_wuser_9_reg				(desc_3_wuser_9_reg[31:0]),
       .desc_3_wuser_10_reg				(desc_3_wuser_10_reg[31:0]),
       .desc_3_wuser_11_reg				(desc_3_wuser_11_reg[31:0]),
       .desc_3_wuser_12_reg				(desc_3_wuser_12_reg[31:0]),
       .desc_3_wuser_13_reg				(desc_3_wuser_13_reg[31:0]),
       .desc_3_wuser_14_reg				(desc_3_wuser_14_reg[31:0]),
       .desc_3_wuser_15_reg				(desc_3_wuser_15_reg[31:0]),
       .desc_4_txn_type_reg				(desc_4_txn_type_reg[31:0]),
       .desc_4_size_reg					(desc_4_size_reg[31:0]),
       .desc_4_data_offset_reg			(desc_4_data_offset_reg[31:0]),
       .desc_4_data_host_addr_0_reg		(desc_4_data_host_addr_0_reg[31:0]),
       .desc_4_data_host_addr_1_reg		(desc_4_data_host_addr_1_reg[31:0]),
       .desc_4_data_host_addr_2_reg		(desc_4_data_host_addr_2_reg[31:0]),
       .desc_4_data_host_addr_3_reg		(desc_4_data_host_addr_3_reg[31:0]),
       .desc_4_wstrb_host_addr_0_reg		(desc_4_wstrb_host_addr_0_reg[31:0]),
       .desc_4_wstrb_host_addr_1_reg		(desc_4_wstrb_host_addr_1_reg[31:0]),
       .desc_4_wstrb_host_addr_2_reg		(desc_4_wstrb_host_addr_2_reg[31:0]),
       .desc_4_wstrb_host_addr_3_reg		(desc_4_wstrb_host_addr_3_reg[31:0]),
       .desc_4_axsize_reg				(desc_4_axsize_reg[31:0]),
       .desc_4_attr_reg					(desc_4_attr_reg[31:0]),
       .desc_4_axaddr_0_reg				(desc_4_axaddr_0_reg[31:0]),
       .desc_4_axaddr_1_reg				(desc_4_axaddr_1_reg[31:0]),
       .desc_4_axaddr_2_reg				(desc_4_axaddr_2_reg[31:0]),
       .desc_4_axaddr_3_reg				(desc_4_axaddr_3_reg[31:0]),
       .desc_4_axid_0_reg				(desc_4_axid_0_reg[31:0]),
       .desc_4_axid_1_reg				(desc_4_axid_1_reg[31:0]),
       .desc_4_axid_2_reg				(desc_4_axid_2_reg[31:0]),
       .desc_4_axid_3_reg				(desc_4_axid_3_reg[31:0]),
       .desc_4_axuser_0_reg				(desc_4_axuser_0_reg[31:0]),
       .desc_4_axuser_1_reg				(desc_4_axuser_1_reg[31:0]),
       .desc_4_axuser_2_reg				(desc_4_axuser_2_reg[31:0]),
       .desc_4_axuser_3_reg				(desc_4_axuser_3_reg[31:0]),
       .desc_4_axuser_4_reg				(desc_4_axuser_4_reg[31:0]),
       .desc_4_axuser_5_reg				(desc_4_axuser_5_reg[31:0]),
       .desc_4_axuser_6_reg				(desc_4_axuser_6_reg[31:0]),
       .desc_4_axuser_7_reg				(desc_4_axuser_7_reg[31:0]),
       .desc_4_axuser_8_reg				(desc_4_axuser_8_reg[31:0]),
       .desc_4_axuser_9_reg				(desc_4_axuser_9_reg[31:0]),
       .desc_4_axuser_10_reg				(desc_4_axuser_10_reg[31:0]),
       .desc_4_axuser_11_reg				(desc_4_axuser_11_reg[31:0]),
       .desc_4_axuser_12_reg				(desc_4_axuser_12_reg[31:0]),
       .desc_4_axuser_13_reg				(desc_4_axuser_13_reg[31:0]),
       .desc_4_axuser_14_reg				(desc_4_axuser_14_reg[31:0]),
       .desc_4_axuser_15_reg				(desc_4_axuser_15_reg[31:0]),
       .desc_4_xuser_0_reg				(desc_4_xuser_0_reg[31:0]),
       .desc_4_xuser_1_reg				(desc_4_xuser_1_reg[31:0]),
       .desc_4_xuser_2_reg				(desc_4_xuser_2_reg[31:0]),
       .desc_4_xuser_3_reg				(desc_4_xuser_3_reg[31:0]),
       .desc_4_xuser_4_reg				(desc_4_xuser_4_reg[31:0]),
       .desc_4_xuser_5_reg				(desc_4_xuser_5_reg[31:0]),
       .desc_4_xuser_6_reg				(desc_4_xuser_6_reg[31:0]),
       .desc_4_xuser_7_reg				(desc_4_xuser_7_reg[31:0]),
       .desc_4_xuser_8_reg				(desc_4_xuser_8_reg[31:0]),
       .desc_4_xuser_9_reg				(desc_4_xuser_9_reg[31:0]),
       .desc_4_xuser_10_reg				(desc_4_xuser_10_reg[31:0]),
       .desc_4_xuser_11_reg				(desc_4_xuser_11_reg[31:0]),
       .desc_4_xuser_12_reg				(desc_4_xuser_12_reg[31:0]),
       .desc_4_xuser_13_reg				(desc_4_xuser_13_reg[31:0]),
       .desc_4_xuser_14_reg				(desc_4_xuser_14_reg[31:0]),
       .desc_4_xuser_15_reg				(desc_4_xuser_15_reg[31:0]),
       .desc_4_wuser_0_reg				(desc_4_wuser_0_reg[31:0]),
       .desc_4_wuser_1_reg				(desc_4_wuser_1_reg[31:0]),
       .desc_4_wuser_2_reg				(desc_4_wuser_2_reg[31:0]),
       .desc_4_wuser_3_reg				(desc_4_wuser_3_reg[31:0]),
       .desc_4_wuser_4_reg				(desc_4_wuser_4_reg[31:0]),
       .desc_4_wuser_5_reg				(desc_4_wuser_5_reg[31:0]),
       .desc_4_wuser_6_reg				(desc_4_wuser_6_reg[31:0]),
       .desc_4_wuser_7_reg				(desc_4_wuser_7_reg[31:0]),
       .desc_4_wuser_8_reg				(desc_4_wuser_8_reg[31:0]),
       .desc_4_wuser_9_reg				(desc_4_wuser_9_reg[31:0]),
       .desc_4_wuser_10_reg				(desc_4_wuser_10_reg[31:0]),
       .desc_4_wuser_11_reg				(desc_4_wuser_11_reg[31:0]),
       .desc_4_wuser_12_reg				(desc_4_wuser_12_reg[31:0]),
       .desc_4_wuser_13_reg				(desc_4_wuser_13_reg[31:0]),
       .desc_4_wuser_14_reg				(desc_4_wuser_14_reg[31:0]),
       .desc_4_wuser_15_reg				(desc_4_wuser_15_reg[31:0]),
       .desc_5_txn_type_reg				(desc_5_txn_type_reg[31:0]),
       .desc_5_size_reg					(desc_5_size_reg[31:0]),
       .desc_5_data_offset_reg			(desc_5_data_offset_reg[31:0]),
       .desc_5_data_host_addr_0_reg		(desc_5_data_host_addr_0_reg[31:0]),
       .desc_5_data_host_addr_1_reg		(desc_5_data_host_addr_1_reg[31:0]),
       .desc_5_data_host_addr_2_reg		(desc_5_data_host_addr_2_reg[31:0]),
       .desc_5_data_host_addr_3_reg		(desc_5_data_host_addr_3_reg[31:0]),
       .desc_5_wstrb_host_addr_0_reg		(desc_5_wstrb_host_addr_0_reg[31:0]),
       .desc_5_wstrb_host_addr_1_reg		(desc_5_wstrb_host_addr_1_reg[31:0]),
       .desc_5_wstrb_host_addr_2_reg		(desc_5_wstrb_host_addr_2_reg[31:0]),
       .desc_5_wstrb_host_addr_3_reg		(desc_5_wstrb_host_addr_3_reg[31:0]),
       .desc_5_axsize_reg				(desc_5_axsize_reg[31:0]),
       .desc_5_attr_reg					(desc_5_attr_reg[31:0]),
       .desc_5_axaddr_0_reg				(desc_5_axaddr_0_reg[31:0]),
       .desc_5_axaddr_1_reg				(desc_5_axaddr_1_reg[31:0]),
       .desc_5_axaddr_2_reg				(desc_5_axaddr_2_reg[31:0]),
       .desc_5_axaddr_3_reg				(desc_5_axaddr_3_reg[31:0]),
       .desc_5_axid_0_reg				(desc_5_axid_0_reg[31:0]),
       .desc_5_axid_1_reg				(desc_5_axid_1_reg[31:0]),
       .desc_5_axid_2_reg				(desc_5_axid_2_reg[31:0]),
       .desc_5_axid_3_reg				(desc_5_axid_3_reg[31:0]),
       .desc_5_axuser_0_reg				(desc_5_axuser_0_reg[31:0]),
       .desc_5_axuser_1_reg				(desc_5_axuser_1_reg[31:0]),
       .desc_5_axuser_2_reg				(desc_5_axuser_2_reg[31:0]),
       .desc_5_axuser_3_reg				(desc_5_axuser_3_reg[31:0]),
       .desc_5_axuser_4_reg				(desc_5_axuser_4_reg[31:0]),
       .desc_5_axuser_5_reg				(desc_5_axuser_5_reg[31:0]),
       .desc_5_axuser_6_reg				(desc_5_axuser_6_reg[31:0]),
       .desc_5_axuser_7_reg				(desc_5_axuser_7_reg[31:0]),
       .desc_5_axuser_8_reg				(desc_5_axuser_8_reg[31:0]),
       .desc_5_axuser_9_reg				(desc_5_axuser_9_reg[31:0]),
       .desc_5_axuser_10_reg				(desc_5_axuser_10_reg[31:0]),
       .desc_5_axuser_11_reg				(desc_5_axuser_11_reg[31:0]),
       .desc_5_axuser_12_reg				(desc_5_axuser_12_reg[31:0]),
       .desc_5_axuser_13_reg				(desc_5_axuser_13_reg[31:0]),
       .desc_5_axuser_14_reg				(desc_5_axuser_14_reg[31:0]),
       .desc_5_axuser_15_reg				(desc_5_axuser_15_reg[31:0]),
       .desc_5_xuser_0_reg				(desc_5_xuser_0_reg[31:0]),
       .desc_5_xuser_1_reg				(desc_5_xuser_1_reg[31:0]),
       .desc_5_xuser_2_reg				(desc_5_xuser_2_reg[31:0]),
       .desc_5_xuser_3_reg				(desc_5_xuser_3_reg[31:0]),
       .desc_5_xuser_4_reg				(desc_5_xuser_4_reg[31:0]),
       .desc_5_xuser_5_reg				(desc_5_xuser_5_reg[31:0]),
       .desc_5_xuser_6_reg				(desc_5_xuser_6_reg[31:0]),
       .desc_5_xuser_7_reg				(desc_5_xuser_7_reg[31:0]),
       .desc_5_xuser_8_reg				(desc_5_xuser_8_reg[31:0]),
       .desc_5_xuser_9_reg				(desc_5_xuser_9_reg[31:0]),
       .desc_5_xuser_10_reg				(desc_5_xuser_10_reg[31:0]),
       .desc_5_xuser_11_reg				(desc_5_xuser_11_reg[31:0]),
       .desc_5_xuser_12_reg				(desc_5_xuser_12_reg[31:0]),
       .desc_5_xuser_13_reg				(desc_5_xuser_13_reg[31:0]),
       .desc_5_xuser_14_reg				(desc_5_xuser_14_reg[31:0]),
       .desc_5_xuser_15_reg				(desc_5_xuser_15_reg[31:0]),
       .desc_5_wuser_0_reg				(desc_5_wuser_0_reg[31:0]),
       .desc_5_wuser_1_reg				(desc_5_wuser_1_reg[31:0]),
       .desc_5_wuser_2_reg				(desc_5_wuser_2_reg[31:0]),
       .desc_5_wuser_3_reg				(desc_5_wuser_3_reg[31:0]),
       .desc_5_wuser_4_reg				(desc_5_wuser_4_reg[31:0]),
       .desc_5_wuser_5_reg				(desc_5_wuser_5_reg[31:0]),
       .desc_5_wuser_6_reg				(desc_5_wuser_6_reg[31:0]),
       .desc_5_wuser_7_reg				(desc_5_wuser_7_reg[31:0]),
       .desc_5_wuser_8_reg				(desc_5_wuser_8_reg[31:0]),
       .desc_5_wuser_9_reg				(desc_5_wuser_9_reg[31:0]),
       .desc_5_wuser_10_reg				(desc_5_wuser_10_reg[31:0]),
       .desc_5_wuser_11_reg				(desc_5_wuser_11_reg[31:0]),
       .desc_5_wuser_12_reg				(desc_5_wuser_12_reg[31:0]),
       .desc_5_wuser_13_reg				(desc_5_wuser_13_reg[31:0]),
       .desc_5_wuser_14_reg				(desc_5_wuser_14_reg[31:0]),
       .desc_5_wuser_15_reg				(desc_5_wuser_15_reg[31:0]),
       .desc_6_txn_type_reg				(desc_6_txn_type_reg[31:0]),
       .desc_6_size_reg					(desc_6_size_reg[31:0]),
       .desc_6_data_offset_reg			(desc_6_data_offset_reg[31:0]),
       .desc_6_data_host_addr_0_reg		(desc_6_data_host_addr_0_reg[31:0]),
       .desc_6_data_host_addr_1_reg		(desc_6_data_host_addr_1_reg[31:0]),
       .desc_6_data_host_addr_2_reg		(desc_6_data_host_addr_2_reg[31:0]),
       .desc_6_data_host_addr_3_reg		(desc_6_data_host_addr_3_reg[31:0]),
       .desc_6_wstrb_host_addr_0_reg		(desc_6_wstrb_host_addr_0_reg[31:0]),
       .desc_6_wstrb_host_addr_1_reg		(desc_6_wstrb_host_addr_1_reg[31:0]),
       .desc_6_wstrb_host_addr_2_reg		(desc_6_wstrb_host_addr_2_reg[31:0]),
       .desc_6_wstrb_host_addr_3_reg		(desc_6_wstrb_host_addr_3_reg[31:0]),
       .desc_6_axsize_reg				(desc_6_axsize_reg[31:0]),
       .desc_6_attr_reg					(desc_6_attr_reg[31:0]),
       .desc_6_axaddr_0_reg				(desc_6_axaddr_0_reg[31:0]),
       .desc_6_axaddr_1_reg				(desc_6_axaddr_1_reg[31:0]),
       .desc_6_axaddr_2_reg				(desc_6_axaddr_2_reg[31:0]),
       .desc_6_axaddr_3_reg				(desc_6_axaddr_3_reg[31:0]),
       .desc_6_axid_0_reg				(desc_6_axid_0_reg[31:0]),
       .desc_6_axid_1_reg				(desc_6_axid_1_reg[31:0]),
       .desc_6_axid_2_reg				(desc_6_axid_2_reg[31:0]),
       .desc_6_axid_3_reg				(desc_6_axid_3_reg[31:0]),
       .desc_6_axuser_0_reg				(desc_6_axuser_0_reg[31:0]),
       .desc_6_axuser_1_reg				(desc_6_axuser_1_reg[31:0]),
       .desc_6_axuser_2_reg				(desc_6_axuser_2_reg[31:0]),
       .desc_6_axuser_3_reg				(desc_6_axuser_3_reg[31:0]),
       .desc_6_axuser_4_reg				(desc_6_axuser_4_reg[31:0]),
       .desc_6_axuser_5_reg				(desc_6_axuser_5_reg[31:0]),
       .desc_6_axuser_6_reg				(desc_6_axuser_6_reg[31:0]),
       .desc_6_axuser_7_reg				(desc_6_axuser_7_reg[31:0]),
       .desc_6_axuser_8_reg				(desc_6_axuser_8_reg[31:0]),
       .desc_6_axuser_9_reg				(desc_6_axuser_9_reg[31:0]),
       .desc_6_axuser_10_reg				(desc_6_axuser_10_reg[31:0]),
       .desc_6_axuser_11_reg				(desc_6_axuser_11_reg[31:0]),
       .desc_6_axuser_12_reg				(desc_6_axuser_12_reg[31:0]),
       .desc_6_axuser_13_reg				(desc_6_axuser_13_reg[31:0]),
       .desc_6_axuser_14_reg				(desc_6_axuser_14_reg[31:0]),
       .desc_6_axuser_15_reg				(desc_6_axuser_15_reg[31:0]),
       .desc_6_xuser_0_reg				(desc_6_xuser_0_reg[31:0]),
       .desc_6_xuser_1_reg				(desc_6_xuser_1_reg[31:0]),
       .desc_6_xuser_2_reg				(desc_6_xuser_2_reg[31:0]),
       .desc_6_xuser_3_reg				(desc_6_xuser_3_reg[31:0]),
       .desc_6_xuser_4_reg				(desc_6_xuser_4_reg[31:0]),
       .desc_6_xuser_5_reg				(desc_6_xuser_5_reg[31:0]),
       .desc_6_xuser_6_reg				(desc_6_xuser_6_reg[31:0]),
       .desc_6_xuser_7_reg				(desc_6_xuser_7_reg[31:0]),
       .desc_6_xuser_8_reg				(desc_6_xuser_8_reg[31:0]),
       .desc_6_xuser_9_reg				(desc_6_xuser_9_reg[31:0]),
       .desc_6_xuser_10_reg				(desc_6_xuser_10_reg[31:0]),
       .desc_6_xuser_11_reg				(desc_6_xuser_11_reg[31:0]),
       .desc_6_xuser_12_reg				(desc_6_xuser_12_reg[31:0]),
       .desc_6_xuser_13_reg				(desc_6_xuser_13_reg[31:0]),
       .desc_6_xuser_14_reg				(desc_6_xuser_14_reg[31:0]),
       .desc_6_xuser_15_reg				(desc_6_xuser_15_reg[31:0]),
       .desc_6_wuser_0_reg				(desc_6_wuser_0_reg[31:0]),
       .desc_6_wuser_1_reg				(desc_6_wuser_1_reg[31:0]),
       .desc_6_wuser_2_reg				(desc_6_wuser_2_reg[31:0]),
       .desc_6_wuser_3_reg				(desc_6_wuser_3_reg[31:0]),
       .desc_6_wuser_4_reg				(desc_6_wuser_4_reg[31:0]),
       .desc_6_wuser_5_reg				(desc_6_wuser_5_reg[31:0]),
       .desc_6_wuser_6_reg				(desc_6_wuser_6_reg[31:0]),
       .desc_6_wuser_7_reg				(desc_6_wuser_7_reg[31:0]),
       .desc_6_wuser_8_reg				(desc_6_wuser_8_reg[31:0]),
       .desc_6_wuser_9_reg				(desc_6_wuser_9_reg[31:0]),
       .desc_6_wuser_10_reg				(desc_6_wuser_10_reg[31:0]),
       .desc_6_wuser_11_reg				(desc_6_wuser_11_reg[31:0]),
       .desc_6_wuser_12_reg				(desc_6_wuser_12_reg[31:0]),
       .desc_6_wuser_13_reg				(desc_6_wuser_13_reg[31:0]),
       .desc_6_wuser_14_reg				(desc_6_wuser_14_reg[31:0]),
       .desc_6_wuser_15_reg				(desc_6_wuser_15_reg[31:0]),
       .desc_7_txn_type_reg				(desc_7_txn_type_reg[31:0]),
       .desc_7_size_reg					(desc_7_size_reg[31:0]),
       .desc_7_data_offset_reg			(desc_7_data_offset_reg[31:0]),
       .desc_7_data_host_addr_0_reg		(desc_7_data_host_addr_0_reg[31:0]),
       .desc_7_data_host_addr_1_reg		(desc_7_data_host_addr_1_reg[31:0]),
       .desc_7_data_host_addr_2_reg		(desc_7_data_host_addr_2_reg[31:0]),
       .desc_7_data_host_addr_3_reg		(desc_7_data_host_addr_3_reg[31:0]),
       .desc_7_wstrb_host_addr_0_reg		(desc_7_wstrb_host_addr_0_reg[31:0]),
       .desc_7_wstrb_host_addr_1_reg		(desc_7_wstrb_host_addr_1_reg[31:0]),
       .desc_7_wstrb_host_addr_2_reg		(desc_7_wstrb_host_addr_2_reg[31:0]),
       .desc_7_wstrb_host_addr_3_reg		(desc_7_wstrb_host_addr_3_reg[31:0]),
       .desc_7_axsize_reg				(desc_7_axsize_reg[31:0]),
       .desc_7_attr_reg					(desc_7_attr_reg[31:0]),
       .desc_7_axaddr_0_reg				(desc_7_axaddr_0_reg[31:0]),
       .desc_7_axaddr_1_reg				(desc_7_axaddr_1_reg[31:0]),
       .desc_7_axaddr_2_reg				(desc_7_axaddr_2_reg[31:0]),
       .desc_7_axaddr_3_reg				(desc_7_axaddr_3_reg[31:0]),
       .desc_7_axid_0_reg				(desc_7_axid_0_reg[31:0]),
       .desc_7_axid_1_reg				(desc_7_axid_1_reg[31:0]),
       .desc_7_axid_2_reg				(desc_7_axid_2_reg[31:0]),
       .desc_7_axid_3_reg				(desc_7_axid_3_reg[31:0]),
       .desc_7_axuser_0_reg				(desc_7_axuser_0_reg[31:0]),
       .desc_7_axuser_1_reg				(desc_7_axuser_1_reg[31:0]),
       .desc_7_axuser_2_reg				(desc_7_axuser_2_reg[31:0]),
       .desc_7_axuser_3_reg				(desc_7_axuser_3_reg[31:0]),
       .desc_7_axuser_4_reg				(desc_7_axuser_4_reg[31:0]),
       .desc_7_axuser_5_reg				(desc_7_axuser_5_reg[31:0]),
       .desc_7_axuser_6_reg				(desc_7_axuser_6_reg[31:0]),
       .desc_7_axuser_7_reg				(desc_7_axuser_7_reg[31:0]),
       .desc_7_axuser_8_reg				(desc_7_axuser_8_reg[31:0]),
       .desc_7_axuser_9_reg				(desc_7_axuser_9_reg[31:0]),
       .desc_7_axuser_10_reg				(desc_7_axuser_10_reg[31:0]),
       .desc_7_axuser_11_reg				(desc_7_axuser_11_reg[31:0]),
       .desc_7_axuser_12_reg				(desc_7_axuser_12_reg[31:0]),
       .desc_7_axuser_13_reg				(desc_7_axuser_13_reg[31:0]),
       .desc_7_axuser_14_reg				(desc_7_axuser_14_reg[31:0]),
       .desc_7_axuser_15_reg				(desc_7_axuser_15_reg[31:0]),
       .desc_7_xuser_0_reg				(desc_7_xuser_0_reg[31:0]),
       .desc_7_xuser_1_reg				(desc_7_xuser_1_reg[31:0]),
       .desc_7_xuser_2_reg				(desc_7_xuser_2_reg[31:0]),
       .desc_7_xuser_3_reg				(desc_7_xuser_3_reg[31:0]),
       .desc_7_xuser_4_reg				(desc_7_xuser_4_reg[31:0]),
       .desc_7_xuser_5_reg				(desc_7_xuser_5_reg[31:0]),
       .desc_7_xuser_6_reg				(desc_7_xuser_6_reg[31:0]),
       .desc_7_xuser_7_reg				(desc_7_xuser_7_reg[31:0]),
       .desc_7_xuser_8_reg				(desc_7_xuser_8_reg[31:0]),
       .desc_7_xuser_9_reg				(desc_7_xuser_9_reg[31:0]),
       .desc_7_xuser_10_reg				(desc_7_xuser_10_reg[31:0]),
       .desc_7_xuser_11_reg				(desc_7_xuser_11_reg[31:0]),
       .desc_7_xuser_12_reg				(desc_7_xuser_12_reg[31:0]),
       .desc_7_xuser_13_reg				(desc_7_xuser_13_reg[31:0]),
       .desc_7_xuser_14_reg				(desc_7_xuser_14_reg[31:0]),
       .desc_7_xuser_15_reg				(desc_7_xuser_15_reg[31:0]),
       .desc_7_wuser_0_reg				(desc_7_wuser_0_reg[31:0]),
       .desc_7_wuser_1_reg				(desc_7_wuser_1_reg[31:0]),
       .desc_7_wuser_2_reg				(desc_7_wuser_2_reg[31:0]),
       .desc_7_wuser_3_reg				(desc_7_wuser_3_reg[31:0]),
       .desc_7_wuser_4_reg				(desc_7_wuser_4_reg[31:0]),
       .desc_7_wuser_5_reg				(desc_7_wuser_5_reg[31:0]),
       .desc_7_wuser_6_reg				(desc_7_wuser_6_reg[31:0]),
       .desc_7_wuser_7_reg				(desc_7_wuser_7_reg[31:0]),
       .desc_7_wuser_8_reg				(desc_7_wuser_8_reg[31:0]),
       .desc_7_wuser_9_reg				(desc_7_wuser_9_reg[31:0]),
       .desc_7_wuser_10_reg				(desc_7_wuser_10_reg[31:0]),
       .desc_7_wuser_11_reg				(desc_7_wuser_11_reg[31:0]),
       .desc_7_wuser_12_reg				(desc_7_wuser_12_reg[31:0]),
       .desc_7_wuser_13_reg				(desc_7_wuser_13_reg[31:0]),
       .desc_7_wuser_14_reg				(desc_7_wuser_14_reg[31:0]),
       .desc_7_wuser_15_reg				(desc_7_wuser_15_reg[31:0]),
       .desc_8_txn_type_reg				(desc_8_txn_type_reg[31:0]),
       .desc_8_size_reg					(desc_8_size_reg[31:0]),
       .desc_8_data_offset_reg			(desc_8_data_offset_reg[31:0]),
       .desc_8_data_host_addr_0_reg		(desc_8_data_host_addr_0_reg[31:0]),
       .desc_8_data_host_addr_1_reg		(desc_8_data_host_addr_1_reg[31:0]),
       .desc_8_data_host_addr_2_reg		(desc_8_data_host_addr_2_reg[31:0]),
       .desc_8_data_host_addr_3_reg		(desc_8_data_host_addr_3_reg[31:0]),
       .desc_8_wstrb_host_addr_0_reg		(desc_8_wstrb_host_addr_0_reg[31:0]),
       .desc_8_wstrb_host_addr_1_reg		(desc_8_wstrb_host_addr_1_reg[31:0]),
       .desc_8_wstrb_host_addr_2_reg		(desc_8_wstrb_host_addr_2_reg[31:0]),
       .desc_8_wstrb_host_addr_3_reg		(desc_8_wstrb_host_addr_3_reg[31:0]),
       .desc_8_axsize_reg				(desc_8_axsize_reg[31:0]),
       .desc_8_attr_reg					(desc_8_attr_reg[31:0]),
       .desc_8_axaddr_0_reg				(desc_8_axaddr_0_reg[31:0]),
       .desc_8_axaddr_1_reg				(desc_8_axaddr_1_reg[31:0]),
       .desc_8_axaddr_2_reg				(desc_8_axaddr_2_reg[31:0]),
       .desc_8_axaddr_3_reg				(desc_8_axaddr_3_reg[31:0]),
       .desc_8_axid_0_reg				(desc_8_axid_0_reg[31:0]),
       .desc_8_axid_1_reg				(desc_8_axid_1_reg[31:0]),
       .desc_8_axid_2_reg				(desc_8_axid_2_reg[31:0]),
       .desc_8_axid_3_reg				(desc_8_axid_3_reg[31:0]),
       .desc_8_axuser_0_reg				(desc_8_axuser_0_reg[31:0]),
       .desc_8_axuser_1_reg				(desc_8_axuser_1_reg[31:0]),
       .desc_8_axuser_2_reg				(desc_8_axuser_2_reg[31:0]),
       .desc_8_axuser_3_reg				(desc_8_axuser_3_reg[31:0]),
       .desc_8_axuser_4_reg				(desc_8_axuser_4_reg[31:0]),
       .desc_8_axuser_5_reg				(desc_8_axuser_5_reg[31:0]),
       .desc_8_axuser_6_reg				(desc_8_axuser_6_reg[31:0]),
       .desc_8_axuser_7_reg				(desc_8_axuser_7_reg[31:0]),
       .desc_8_axuser_8_reg				(desc_8_axuser_8_reg[31:0]),
       .desc_8_axuser_9_reg				(desc_8_axuser_9_reg[31:0]),
       .desc_8_axuser_10_reg				(desc_8_axuser_10_reg[31:0]),
       .desc_8_axuser_11_reg				(desc_8_axuser_11_reg[31:0]),
       .desc_8_axuser_12_reg				(desc_8_axuser_12_reg[31:0]),
       .desc_8_axuser_13_reg				(desc_8_axuser_13_reg[31:0]),
       .desc_8_axuser_14_reg				(desc_8_axuser_14_reg[31:0]),
       .desc_8_axuser_15_reg				(desc_8_axuser_15_reg[31:0]),
       .desc_8_xuser_0_reg				(desc_8_xuser_0_reg[31:0]),
       .desc_8_xuser_1_reg				(desc_8_xuser_1_reg[31:0]),
       .desc_8_xuser_2_reg				(desc_8_xuser_2_reg[31:0]),
       .desc_8_xuser_3_reg				(desc_8_xuser_3_reg[31:0]),
       .desc_8_xuser_4_reg				(desc_8_xuser_4_reg[31:0]),
       .desc_8_xuser_5_reg				(desc_8_xuser_5_reg[31:0]),
       .desc_8_xuser_6_reg				(desc_8_xuser_6_reg[31:0]),
       .desc_8_xuser_7_reg				(desc_8_xuser_7_reg[31:0]),
       .desc_8_xuser_8_reg				(desc_8_xuser_8_reg[31:0]),
       .desc_8_xuser_9_reg				(desc_8_xuser_9_reg[31:0]),
       .desc_8_xuser_10_reg				(desc_8_xuser_10_reg[31:0]),
       .desc_8_xuser_11_reg				(desc_8_xuser_11_reg[31:0]),
       .desc_8_xuser_12_reg				(desc_8_xuser_12_reg[31:0]),
       .desc_8_xuser_13_reg				(desc_8_xuser_13_reg[31:0]),
       .desc_8_xuser_14_reg				(desc_8_xuser_14_reg[31:0]),
       .desc_8_xuser_15_reg				(desc_8_xuser_15_reg[31:0]),
       .desc_8_wuser_0_reg				(desc_8_wuser_0_reg[31:0]),
       .desc_8_wuser_1_reg				(desc_8_wuser_1_reg[31:0]),
       .desc_8_wuser_2_reg				(desc_8_wuser_2_reg[31:0]),
       .desc_8_wuser_3_reg				(desc_8_wuser_3_reg[31:0]),
       .desc_8_wuser_4_reg				(desc_8_wuser_4_reg[31:0]),
       .desc_8_wuser_5_reg				(desc_8_wuser_5_reg[31:0]),
       .desc_8_wuser_6_reg				(desc_8_wuser_6_reg[31:0]),
       .desc_8_wuser_7_reg				(desc_8_wuser_7_reg[31:0]),
       .desc_8_wuser_8_reg				(desc_8_wuser_8_reg[31:0]),
       .desc_8_wuser_9_reg				(desc_8_wuser_9_reg[31:0]),
       .desc_8_wuser_10_reg				(desc_8_wuser_10_reg[31:0]),
       .desc_8_wuser_11_reg				(desc_8_wuser_11_reg[31:0]),
       .desc_8_wuser_12_reg				(desc_8_wuser_12_reg[31:0]),
       .desc_8_wuser_13_reg				(desc_8_wuser_13_reg[31:0]),
       .desc_8_wuser_14_reg				(desc_8_wuser_14_reg[31:0]),
       .desc_8_wuser_15_reg				(desc_8_wuser_15_reg[31:0]),
       .desc_9_txn_type_reg				(desc_9_txn_type_reg[31:0]),
       .desc_9_size_reg					(desc_9_size_reg[31:0]),
       .desc_9_data_offset_reg			(desc_9_data_offset_reg[31:0]),
       .desc_9_data_host_addr_0_reg		(desc_9_data_host_addr_0_reg[31:0]),
       .desc_9_data_host_addr_1_reg		(desc_9_data_host_addr_1_reg[31:0]),
       .desc_9_data_host_addr_2_reg		(desc_9_data_host_addr_2_reg[31:0]),
       .desc_9_data_host_addr_3_reg		(desc_9_data_host_addr_3_reg[31:0]),
       .desc_9_wstrb_host_addr_0_reg		(desc_9_wstrb_host_addr_0_reg[31:0]),
       .desc_9_wstrb_host_addr_1_reg		(desc_9_wstrb_host_addr_1_reg[31:0]),
       .desc_9_wstrb_host_addr_2_reg		(desc_9_wstrb_host_addr_2_reg[31:0]),
       .desc_9_wstrb_host_addr_3_reg		(desc_9_wstrb_host_addr_3_reg[31:0]),
       .desc_9_axsize_reg				(desc_9_axsize_reg[31:0]),
       .desc_9_attr_reg					(desc_9_attr_reg[31:0]),
       .desc_9_axaddr_0_reg				(desc_9_axaddr_0_reg[31:0]),
       .desc_9_axaddr_1_reg				(desc_9_axaddr_1_reg[31:0]),
       .desc_9_axaddr_2_reg				(desc_9_axaddr_2_reg[31:0]),
       .desc_9_axaddr_3_reg				(desc_9_axaddr_3_reg[31:0]),
       .desc_9_axid_0_reg				(desc_9_axid_0_reg[31:0]),
       .desc_9_axid_1_reg				(desc_9_axid_1_reg[31:0]),
       .desc_9_axid_2_reg				(desc_9_axid_2_reg[31:0]),
       .desc_9_axid_3_reg				(desc_9_axid_3_reg[31:0]),
       .desc_9_axuser_0_reg				(desc_9_axuser_0_reg[31:0]),
       .desc_9_axuser_1_reg				(desc_9_axuser_1_reg[31:0]),
       .desc_9_axuser_2_reg				(desc_9_axuser_2_reg[31:0]),
       .desc_9_axuser_3_reg				(desc_9_axuser_3_reg[31:0]),
       .desc_9_axuser_4_reg				(desc_9_axuser_4_reg[31:0]),
       .desc_9_axuser_5_reg				(desc_9_axuser_5_reg[31:0]),
       .desc_9_axuser_6_reg				(desc_9_axuser_6_reg[31:0]),
       .desc_9_axuser_7_reg				(desc_9_axuser_7_reg[31:0]),
       .desc_9_axuser_8_reg				(desc_9_axuser_8_reg[31:0]),
       .desc_9_axuser_9_reg				(desc_9_axuser_9_reg[31:0]),
       .desc_9_axuser_10_reg				(desc_9_axuser_10_reg[31:0]),
       .desc_9_axuser_11_reg				(desc_9_axuser_11_reg[31:0]),
       .desc_9_axuser_12_reg				(desc_9_axuser_12_reg[31:0]),
       .desc_9_axuser_13_reg				(desc_9_axuser_13_reg[31:0]),
       .desc_9_axuser_14_reg				(desc_9_axuser_14_reg[31:0]),
       .desc_9_axuser_15_reg				(desc_9_axuser_15_reg[31:0]),
       .desc_9_xuser_0_reg				(desc_9_xuser_0_reg[31:0]),
       .desc_9_xuser_1_reg				(desc_9_xuser_1_reg[31:0]),
       .desc_9_xuser_2_reg				(desc_9_xuser_2_reg[31:0]),
       .desc_9_xuser_3_reg				(desc_9_xuser_3_reg[31:0]),
       .desc_9_xuser_4_reg				(desc_9_xuser_4_reg[31:0]),
       .desc_9_xuser_5_reg				(desc_9_xuser_5_reg[31:0]),
       .desc_9_xuser_6_reg				(desc_9_xuser_6_reg[31:0]),
       .desc_9_xuser_7_reg				(desc_9_xuser_7_reg[31:0]),
       .desc_9_xuser_8_reg				(desc_9_xuser_8_reg[31:0]),
       .desc_9_xuser_9_reg				(desc_9_xuser_9_reg[31:0]),
       .desc_9_xuser_10_reg				(desc_9_xuser_10_reg[31:0]),
       .desc_9_xuser_11_reg				(desc_9_xuser_11_reg[31:0]),
       .desc_9_xuser_12_reg				(desc_9_xuser_12_reg[31:0]),
       .desc_9_xuser_13_reg				(desc_9_xuser_13_reg[31:0]),
       .desc_9_xuser_14_reg				(desc_9_xuser_14_reg[31:0]),
       .desc_9_xuser_15_reg				(desc_9_xuser_15_reg[31:0]),
       .desc_9_wuser_0_reg				(desc_9_wuser_0_reg[31:0]),
       .desc_9_wuser_1_reg				(desc_9_wuser_1_reg[31:0]),
       .desc_9_wuser_2_reg				(desc_9_wuser_2_reg[31:0]),
       .desc_9_wuser_3_reg				(desc_9_wuser_3_reg[31:0]),
       .desc_9_wuser_4_reg				(desc_9_wuser_4_reg[31:0]),
       .desc_9_wuser_5_reg				(desc_9_wuser_5_reg[31:0]),
       .desc_9_wuser_6_reg				(desc_9_wuser_6_reg[31:0]),
       .desc_9_wuser_7_reg				(desc_9_wuser_7_reg[31:0]),
       .desc_9_wuser_8_reg				(desc_9_wuser_8_reg[31:0]),
       .desc_9_wuser_9_reg				(desc_9_wuser_9_reg[31:0]),
       .desc_9_wuser_10_reg				(desc_9_wuser_10_reg[31:0]),
       .desc_9_wuser_11_reg				(desc_9_wuser_11_reg[31:0]),
       .desc_9_wuser_12_reg				(desc_9_wuser_12_reg[31:0]),
       .desc_9_wuser_13_reg				(desc_9_wuser_13_reg[31:0]),
       .desc_9_wuser_14_reg				(desc_9_wuser_14_reg[31:0]),
       .desc_9_wuser_15_reg				(desc_9_wuser_15_reg[31:0]),
       .desc_10_txn_type_reg				(desc_10_txn_type_reg[31:0]),
       .desc_10_size_reg					(desc_10_size_reg[31:0]),
       .desc_10_data_offset_reg			(desc_10_data_offset_reg[31:0]),
       .desc_10_data_host_addr_0_reg		(desc_10_data_host_addr_0_reg[31:0]),
       .desc_10_data_host_addr_1_reg		(desc_10_data_host_addr_1_reg[31:0]),
       .desc_10_data_host_addr_2_reg		(desc_10_data_host_addr_2_reg[31:0]),
       .desc_10_data_host_addr_3_reg		(desc_10_data_host_addr_3_reg[31:0]),
       .desc_10_wstrb_host_addr_0_reg	(desc_10_wstrb_host_addr_0_reg[31:0]),
       .desc_10_wstrb_host_addr_1_reg	(desc_10_wstrb_host_addr_1_reg[31:0]),
       .desc_10_wstrb_host_addr_2_reg	(desc_10_wstrb_host_addr_2_reg[31:0]),
       .desc_10_wstrb_host_addr_3_reg	(desc_10_wstrb_host_addr_3_reg[31:0]),
       .desc_10_axsize_reg				(desc_10_axsize_reg[31:0]),
       .desc_10_attr_reg					(desc_10_attr_reg[31:0]),
       .desc_10_axaddr_0_reg				(desc_10_axaddr_0_reg[31:0]),
       .desc_10_axaddr_1_reg				(desc_10_axaddr_1_reg[31:0]),
       .desc_10_axaddr_2_reg				(desc_10_axaddr_2_reg[31:0]),
       .desc_10_axaddr_3_reg				(desc_10_axaddr_3_reg[31:0]),
       .desc_10_axid_0_reg				(desc_10_axid_0_reg[31:0]),
       .desc_10_axid_1_reg				(desc_10_axid_1_reg[31:0]),
       .desc_10_axid_2_reg				(desc_10_axid_2_reg[31:0]),
       .desc_10_axid_3_reg				(desc_10_axid_3_reg[31:0]),
       .desc_10_axuser_0_reg				(desc_10_axuser_0_reg[31:0]),
       .desc_10_axuser_1_reg				(desc_10_axuser_1_reg[31:0]),
       .desc_10_axuser_2_reg				(desc_10_axuser_2_reg[31:0]),
       .desc_10_axuser_3_reg				(desc_10_axuser_3_reg[31:0]),
       .desc_10_axuser_4_reg				(desc_10_axuser_4_reg[31:0]),
       .desc_10_axuser_5_reg				(desc_10_axuser_5_reg[31:0]),
       .desc_10_axuser_6_reg				(desc_10_axuser_6_reg[31:0]),
       .desc_10_axuser_7_reg				(desc_10_axuser_7_reg[31:0]),
       .desc_10_axuser_8_reg				(desc_10_axuser_8_reg[31:0]),
       .desc_10_axuser_9_reg				(desc_10_axuser_9_reg[31:0]),
       .desc_10_axuser_10_reg			(desc_10_axuser_10_reg[31:0]),
       .desc_10_axuser_11_reg			(desc_10_axuser_11_reg[31:0]),
       .desc_10_axuser_12_reg			(desc_10_axuser_12_reg[31:0]),
       .desc_10_axuser_13_reg			(desc_10_axuser_13_reg[31:0]),
       .desc_10_axuser_14_reg			(desc_10_axuser_14_reg[31:0]),
       .desc_10_axuser_15_reg			(desc_10_axuser_15_reg[31:0]),
       .desc_10_xuser_0_reg				(desc_10_xuser_0_reg[31:0]),
       .desc_10_xuser_1_reg				(desc_10_xuser_1_reg[31:0]),
       .desc_10_xuser_2_reg				(desc_10_xuser_2_reg[31:0]),
       .desc_10_xuser_3_reg				(desc_10_xuser_3_reg[31:0]),
       .desc_10_xuser_4_reg				(desc_10_xuser_4_reg[31:0]),
       .desc_10_xuser_5_reg				(desc_10_xuser_5_reg[31:0]),
       .desc_10_xuser_6_reg				(desc_10_xuser_6_reg[31:0]),
       .desc_10_xuser_7_reg				(desc_10_xuser_7_reg[31:0]),
       .desc_10_xuser_8_reg				(desc_10_xuser_8_reg[31:0]),
       .desc_10_xuser_9_reg				(desc_10_xuser_9_reg[31:0]),
       .desc_10_xuser_10_reg				(desc_10_xuser_10_reg[31:0]),
       .desc_10_xuser_11_reg				(desc_10_xuser_11_reg[31:0]),
       .desc_10_xuser_12_reg				(desc_10_xuser_12_reg[31:0]),
       .desc_10_xuser_13_reg				(desc_10_xuser_13_reg[31:0]),
       .desc_10_xuser_14_reg				(desc_10_xuser_14_reg[31:0]),
       .desc_10_xuser_15_reg				(desc_10_xuser_15_reg[31:0]),
       .desc_10_wuser_0_reg				(desc_10_wuser_0_reg[31:0]),
       .desc_10_wuser_1_reg				(desc_10_wuser_1_reg[31:0]),
       .desc_10_wuser_2_reg				(desc_10_wuser_2_reg[31:0]),
       .desc_10_wuser_3_reg				(desc_10_wuser_3_reg[31:0]),
       .desc_10_wuser_4_reg				(desc_10_wuser_4_reg[31:0]),
       .desc_10_wuser_5_reg				(desc_10_wuser_5_reg[31:0]),
       .desc_10_wuser_6_reg				(desc_10_wuser_6_reg[31:0]),
       .desc_10_wuser_7_reg				(desc_10_wuser_7_reg[31:0]),
       .desc_10_wuser_8_reg				(desc_10_wuser_8_reg[31:0]),
       .desc_10_wuser_9_reg				(desc_10_wuser_9_reg[31:0]),
       .desc_10_wuser_10_reg				(desc_10_wuser_10_reg[31:0]),
       .desc_10_wuser_11_reg				(desc_10_wuser_11_reg[31:0]),
       .desc_10_wuser_12_reg				(desc_10_wuser_12_reg[31:0]),
       .desc_10_wuser_13_reg				(desc_10_wuser_13_reg[31:0]),
       .desc_10_wuser_14_reg				(desc_10_wuser_14_reg[31:0]),
       .desc_10_wuser_15_reg				(desc_10_wuser_15_reg[31:0]),
       .desc_11_txn_type_reg				(desc_11_txn_type_reg[31:0]),
       .desc_11_size_reg					(desc_11_size_reg[31:0]),
       .desc_11_data_offset_reg			(desc_11_data_offset_reg[31:0]),
       .desc_11_data_host_addr_0_reg		(desc_11_data_host_addr_0_reg[31:0]),
       .desc_11_data_host_addr_1_reg		(desc_11_data_host_addr_1_reg[31:0]),
       .desc_11_data_host_addr_2_reg		(desc_11_data_host_addr_2_reg[31:0]),
       .desc_11_data_host_addr_3_reg		(desc_11_data_host_addr_3_reg[31:0]),
       .desc_11_wstrb_host_addr_0_reg	(desc_11_wstrb_host_addr_0_reg[31:0]),
       .desc_11_wstrb_host_addr_1_reg	(desc_11_wstrb_host_addr_1_reg[31:0]),
       .desc_11_wstrb_host_addr_2_reg	(desc_11_wstrb_host_addr_2_reg[31:0]),
       .desc_11_wstrb_host_addr_3_reg	(desc_11_wstrb_host_addr_3_reg[31:0]),
       .desc_11_axsize_reg				(desc_11_axsize_reg[31:0]),
       .desc_11_attr_reg					(desc_11_attr_reg[31:0]),
       .desc_11_axaddr_0_reg				(desc_11_axaddr_0_reg[31:0]),
       .desc_11_axaddr_1_reg				(desc_11_axaddr_1_reg[31:0]),
       .desc_11_axaddr_2_reg				(desc_11_axaddr_2_reg[31:0]),
       .desc_11_axaddr_3_reg				(desc_11_axaddr_3_reg[31:0]),
       .desc_11_axid_0_reg				(desc_11_axid_0_reg[31:0]),
       .desc_11_axid_1_reg				(desc_11_axid_1_reg[31:0]),
       .desc_11_axid_2_reg				(desc_11_axid_2_reg[31:0]),
       .desc_11_axid_3_reg				(desc_11_axid_3_reg[31:0]),
       .desc_11_axuser_0_reg				(desc_11_axuser_0_reg[31:0]),
       .desc_11_axuser_1_reg				(desc_11_axuser_1_reg[31:0]),
       .desc_11_axuser_2_reg				(desc_11_axuser_2_reg[31:0]),
       .desc_11_axuser_3_reg				(desc_11_axuser_3_reg[31:0]),
       .desc_11_axuser_4_reg				(desc_11_axuser_4_reg[31:0]),
       .desc_11_axuser_5_reg				(desc_11_axuser_5_reg[31:0]),
       .desc_11_axuser_6_reg				(desc_11_axuser_6_reg[31:0]),
       .desc_11_axuser_7_reg				(desc_11_axuser_7_reg[31:0]),
       .desc_11_axuser_8_reg				(desc_11_axuser_8_reg[31:0]),
       .desc_11_axuser_9_reg				(desc_11_axuser_9_reg[31:0]),
       .desc_11_axuser_10_reg			(desc_11_axuser_10_reg[31:0]),
       .desc_11_axuser_11_reg			(desc_11_axuser_11_reg[31:0]),
       .desc_11_axuser_12_reg			(desc_11_axuser_12_reg[31:0]),
       .desc_11_axuser_13_reg			(desc_11_axuser_13_reg[31:0]),
       .desc_11_axuser_14_reg			(desc_11_axuser_14_reg[31:0]),
       .desc_11_axuser_15_reg			(desc_11_axuser_15_reg[31:0]),
       .desc_11_xuser_0_reg				(desc_11_xuser_0_reg[31:0]),
       .desc_11_xuser_1_reg				(desc_11_xuser_1_reg[31:0]),
       .desc_11_xuser_2_reg				(desc_11_xuser_2_reg[31:0]),
       .desc_11_xuser_3_reg				(desc_11_xuser_3_reg[31:0]),
       .desc_11_xuser_4_reg				(desc_11_xuser_4_reg[31:0]),
       .desc_11_xuser_5_reg				(desc_11_xuser_5_reg[31:0]),
       .desc_11_xuser_6_reg				(desc_11_xuser_6_reg[31:0]),
       .desc_11_xuser_7_reg				(desc_11_xuser_7_reg[31:0]),
       .desc_11_xuser_8_reg				(desc_11_xuser_8_reg[31:0]),
       .desc_11_xuser_9_reg				(desc_11_xuser_9_reg[31:0]),
       .desc_11_xuser_10_reg				(desc_11_xuser_10_reg[31:0]),
       .desc_11_xuser_11_reg				(desc_11_xuser_11_reg[31:0]),
       .desc_11_xuser_12_reg				(desc_11_xuser_12_reg[31:0]),
       .desc_11_xuser_13_reg				(desc_11_xuser_13_reg[31:0]),
       .desc_11_xuser_14_reg				(desc_11_xuser_14_reg[31:0]),
       .desc_11_xuser_15_reg				(desc_11_xuser_15_reg[31:0]),
       .desc_11_wuser_0_reg				(desc_11_wuser_0_reg[31:0]),
       .desc_11_wuser_1_reg				(desc_11_wuser_1_reg[31:0]),
       .desc_11_wuser_2_reg				(desc_11_wuser_2_reg[31:0]),
       .desc_11_wuser_3_reg				(desc_11_wuser_3_reg[31:0]),
       .desc_11_wuser_4_reg				(desc_11_wuser_4_reg[31:0]),
       .desc_11_wuser_5_reg				(desc_11_wuser_5_reg[31:0]),
       .desc_11_wuser_6_reg				(desc_11_wuser_6_reg[31:0]),
       .desc_11_wuser_7_reg				(desc_11_wuser_7_reg[31:0]),
       .desc_11_wuser_8_reg				(desc_11_wuser_8_reg[31:0]),
       .desc_11_wuser_9_reg				(desc_11_wuser_9_reg[31:0]),
       .desc_11_wuser_10_reg				(desc_11_wuser_10_reg[31:0]),
       .desc_11_wuser_11_reg				(desc_11_wuser_11_reg[31:0]),
       .desc_11_wuser_12_reg				(desc_11_wuser_12_reg[31:0]),
       .desc_11_wuser_13_reg				(desc_11_wuser_13_reg[31:0]),
       .desc_11_wuser_14_reg				(desc_11_wuser_14_reg[31:0]),
       .desc_11_wuser_15_reg				(desc_11_wuser_15_reg[31:0]),
       .desc_12_txn_type_reg				(desc_12_txn_type_reg[31:0]),
       .desc_12_size_reg					(desc_12_size_reg[31:0]),
       .desc_12_data_offset_reg			(desc_12_data_offset_reg[31:0]),
       .desc_12_data_host_addr_0_reg		(desc_12_data_host_addr_0_reg[31:0]),
       .desc_12_data_host_addr_1_reg		(desc_12_data_host_addr_1_reg[31:0]),
       .desc_12_data_host_addr_2_reg		(desc_12_data_host_addr_2_reg[31:0]),
       .desc_12_data_host_addr_3_reg		(desc_12_data_host_addr_3_reg[31:0]),
       .desc_12_wstrb_host_addr_0_reg	(desc_12_wstrb_host_addr_0_reg[31:0]),
       .desc_12_wstrb_host_addr_1_reg	(desc_12_wstrb_host_addr_1_reg[31:0]),
       .desc_12_wstrb_host_addr_2_reg	(desc_12_wstrb_host_addr_2_reg[31:0]),
       .desc_12_wstrb_host_addr_3_reg	(desc_12_wstrb_host_addr_3_reg[31:0]),
       .desc_12_axsize_reg				(desc_12_axsize_reg[31:0]),
       .desc_12_attr_reg					(desc_12_attr_reg[31:0]),
       .desc_12_axaddr_0_reg				(desc_12_axaddr_0_reg[31:0]),
       .desc_12_axaddr_1_reg				(desc_12_axaddr_1_reg[31:0]),
       .desc_12_axaddr_2_reg				(desc_12_axaddr_2_reg[31:0]),
       .desc_12_axaddr_3_reg				(desc_12_axaddr_3_reg[31:0]),
       .desc_12_axid_0_reg				(desc_12_axid_0_reg[31:0]),
       .desc_12_axid_1_reg				(desc_12_axid_1_reg[31:0]),
       .desc_12_axid_2_reg				(desc_12_axid_2_reg[31:0]),
       .desc_12_axid_3_reg				(desc_12_axid_3_reg[31:0]),
       .desc_12_axuser_0_reg				(desc_12_axuser_0_reg[31:0]),
       .desc_12_axuser_1_reg				(desc_12_axuser_1_reg[31:0]),
       .desc_12_axuser_2_reg				(desc_12_axuser_2_reg[31:0]),
       .desc_12_axuser_3_reg				(desc_12_axuser_3_reg[31:0]),
       .desc_12_axuser_4_reg				(desc_12_axuser_4_reg[31:0]),
       .desc_12_axuser_5_reg				(desc_12_axuser_5_reg[31:0]),
       .desc_12_axuser_6_reg				(desc_12_axuser_6_reg[31:0]),
       .desc_12_axuser_7_reg				(desc_12_axuser_7_reg[31:0]),
       .desc_12_axuser_8_reg				(desc_12_axuser_8_reg[31:0]),
       .desc_12_axuser_9_reg				(desc_12_axuser_9_reg[31:0]),
       .desc_12_axuser_10_reg			(desc_12_axuser_10_reg[31:0]),
       .desc_12_axuser_11_reg			(desc_12_axuser_11_reg[31:0]),
       .desc_12_axuser_12_reg			(desc_12_axuser_12_reg[31:0]),
       .desc_12_axuser_13_reg			(desc_12_axuser_13_reg[31:0]),
       .desc_12_axuser_14_reg			(desc_12_axuser_14_reg[31:0]),
       .desc_12_axuser_15_reg			(desc_12_axuser_15_reg[31:0]),
       .desc_12_xuser_0_reg				(desc_12_xuser_0_reg[31:0]),
       .desc_12_xuser_1_reg				(desc_12_xuser_1_reg[31:0]),
       .desc_12_xuser_2_reg				(desc_12_xuser_2_reg[31:0]),
       .desc_12_xuser_3_reg				(desc_12_xuser_3_reg[31:0]),
       .desc_12_xuser_4_reg				(desc_12_xuser_4_reg[31:0]),
       .desc_12_xuser_5_reg				(desc_12_xuser_5_reg[31:0]),
       .desc_12_xuser_6_reg				(desc_12_xuser_6_reg[31:0]),
       .desc_12_xuser_7_reg				(desc_12_xuser_7_reg[31:0]),
       .desc_12_xuser_8_reg				(desc_12_xuser_8_reg[31:0]),
       .desc_12_xuser_9_reg				(desc_12_xuser_9_reg[31:0]),
       .desc_12_xuser_10_reg				(desc_12_xuser_10_reg[31:0]),
       .desc_12_xuser_11_reg				(desc_12_xuser_11_reg[31:0]),
       .desc_12_xuser_12_reg				(desc_12_xuser_12_reg[31:0]),
       .desc_12_xuser_13_reg				(desc_12_xuser_13_reg[31:0]),
       .desc_12_xuser_14_reg				(desc_12_xuser_14_reg[31:0]),
       .desc_12_xuser_15_reg				(desc_12_xuser_15_reg[31:0]),
       .desc_12_wuser_0_reg				(desc_12_wuser_0_reg[31:0]),
       .desc_12_wuser_1_reg				(desc_12_wuser_1_reg[31:0]),
       .desc_12_wuser_2_reg				(desc_12_wuser_2_reg[31:0]),
       .desc_12_wuser_3_reg				(desc_12_wuser_3_reg[31:0]),
       .desc_12_wuser_4_reg				(desc_12_wuser_4_reg[31:0]),
       .desc_12_wuser_5_reg				(desc_12_wuser_5_reg[31:0]),
       .desc_12_wuser_6_reg				(desc_12_wuser_6_reg[31:0]),
       .desc_12_wuser_7_reg				(desc_12_wuser_7_reg[31:0]),
       .desc_12_wuser_8_reg				(desc_12_wuser_8_reg[31:0]),
       .desc_12_wuser_9_reg				(desc_12_wuser_9_reg[31:0]),
       .desc_12_wuser_10_reg				(desc_12_wuser_10_reg[31:0]),
       .desc_12_wuser_11_reg				(desc_12_wuser_11_reg[31:0]),
       .desc_12_wuser_12_reg				(desc_12_wuser_12_reg[31:0]),
       .desc_12_wuser_13_reg				(desc_12_wuser_13_reg[31:0]),
       .desc_12_wuser_14_reg				(desc_12_wuser_14_reg[31:0]),
       .desc_12_wuser_15_reg				(desc_12_wuser_15_reg[31:0]),
       .desc_13_txn_type_reg				(desc_13_txn_type_reg[31:0]),
       .desc_13_size_reg					(desc_13_size_reg[31:0]),
       .desc_13_data_offset_reg			(desc_13_data_offset_reg[31:0]),
       .desc_13_data_host_addr_0_reg		(desc_13_data_host_addr_0_reg[31:0]),
       .desc_13_data_host_addr_1_reg		(desc_13_data_host_addr_1_reg[31:0]),
       .desc_13_data_host_addr_2_reg		(desc_13_data_host_addr_2_reg[31:0]),
       .desc_13_data_host_addr_3_reg		(desc_13_data_host_addr_3_reg[31:0]),
       .desc_13_wstrb_host_addr_0_reg	(desc_13_wstrb_host_addr_0_reg[31:0]),
       .desc_13_wstrb_host_addr_1_reg	(desc_13_wstrb_host_addr_1_reg[31:0]),
       .desc_13_wstrb_host_addr_2_reg	(desc_13_wstrb_host_addr_2_reg[31:0]),
       .desc_13_wstrb_host_addr_3_reg	(desc_13_wstrb_host_addr_3_reg[31:0]),
       .desc_13_axsize_reg				(desc_13_axsize_reg[31:0]),
       .desc_13_attr_reg					(desc_13_attr_reg[31:0]),
       .desc_13_axaddr_0_reg				(desc_13_axaddr_0_reg[31:0]),
       .desc_13_axaddr_1_reg				(desc_13_axaddr_1_reg[31:0]),
       .desc_13_axaddr_2_reg				(desc_13_axaddr_2_reg[31:0]),
       .desc_13_axaddr_3_reg				(desc_13_axaddr_3_reg[31:0]),
       .desc_13_axid_0_reg				(desc_13_axid_0_reg[31:0]),
       .desc_13_axid_1_reg				(desc_13_axid_1_reg[31:0]),
       .desc_13_axid_2_reg				(desc_13_axid_2_reg[31:0]),
       .desc_13_axid_3_reg				(desc_13_axid_3_reg[31:0]),
       .desc_13_axuser_0_reg				(desc_13_axuser_0_reg[31:0]),
       .desc_13_axuser_1_reg				(desc_13_axuser_1_reg[31:0]),
       .desc_13_axuser_2_reg				(desc_13_axuser_2_reg[31:0]),
       .desc_13_axuser_3_reg				(desc_13_axuser_3_reg[31:0]),
       .desc_13_axuser_4_reg				(desc_13_axuser_4_reg[31:0]),
       .desc_13_axuser_5_reg				(desc_13_axuser_5_reg[31:0]),
       .desc_13_axuser_6_reg				(desc_13_axuser_6_reg[31:0]),
       .desc_13_axuser_7_reg				(desc_13_axuser_7_reg[31:0]),
       .desc_13_axuser_8_reg				(desc_13_axuser_8_reg[31:0]),
       .desc_13_axuser_9_reg				(desc_13_axuser_9_reg[31:0]),
       .desc_13_axuser_10_reg			(desc_13_axuser_10_reg[31:0]),
       .desc_13_axuser_11_reg			(desc_13_axuser_11_reg[31:0]),
       .desc_13_axuser_12_reg			(desc_13_axuser_12_reg[31:0]),
       .desc_13_axuser_13_reg			(desc_13_axuser_13_reg[31:0]),
       .desc_13_axuser_14_reg			(desc_13_axuser_14_reg[31:0]),
       .desc_13_axuser_15_reg			(desc_13_axuser_15_reg[31:0]),
       .desc_13_xuser_0_reg				(desc_13_xuser_0_reg[31:0]),
       .desc_13_xuser_1_reg				(desc_13_xuser_1_reg[31:0]),
       .desc_13_xuser_2_reg				(desc_13_xuser_2_reg[31:0]),
       .desc_13_xuser_3_reg				(desc_13_xuser_3_reg[31:0]),
       .desc_13_xuser_4_reg				(desc_13_xuser_4_reg[31:0]),
       .desc_13_xuser_5_reg				(desc_13_xuser_5_reg[31:0]),
       .desc_13_xuser_6_reg				(desc_13_xuser_6_reg[31:0]),
       .desc_13_xuser_7_reg				(desc_13_xuser_7_reg[31:0]),
       .desc_13_xuser_8_reg				(desc_13_xuser_8_reg[31:0]),
       .desc_13_xuser_9_reg				(desc_13_xuser_9_reg[31:0]),
       .desc_13_xuser_10_reg				(desc_13_xuser_10_reg[31:0]),
       .desc_13_xuser_11_reg				(desc_13_xuser_11_reg[31:0]),
       .desc_13_xuser_12_reg				(desc_13_xuser_12_reg[31:0]),
       .desc_13_xuser_13_reg				(desc_13_xuser_13_reg[31:0]),
       .desc_13_xuser_14_reg				(desc_13_xuser_14_reg[31:0]),
       .desc_13_xuser_15_reg				(desc_13_xuser_15_reg[31:0]),
       .desc_13_wuser_0_reg				(desc_13_wuser_0_reg[31:0]),
       .desc_13_wuser_1_reg				(desc_13_wuser_1_reg[31:0]),
       .desc_13_wuser_2_reg				(desc_13_wuser_2_reg[31:0]),
       .desc_13_wuser_3_reg				(desc_13_wuser_3_reg[31:0]),
       .desc_13_wuser_4_reg				(desc_13_wuser_4_reg[31:0]),
       .desc_13_wuser_5_reg				(desc_13_wuser_5_reg[31:0]),
       .desc_13_wuser_6_reg				(desc_13_wuser_6_reg[31:0]),
       .desc_13_wuser_7_reg				(desc_13_wuser_7_reg[31:0]),
       .desc_13_wuser_8_reg				(desc_13_wuser_8_reg[31:0]),
       .desc_13_wuser_9_reg				(desc_13_wuser_9_reg[31:0]),
       .desc_13_wuser_10_reg				(desc_13_wuser_10_reg[31:0]),
       .desc_13_wuser_11_reg				(desc_13_wuser_11_reg[31:0]),
       .desc_13_wuser_12_reg				(desc_13_wuser_12_reg[31:0]),
       .desc_13_wuser_13_reg				(desc_13_wuser_13_reg[31:0]),
       .desc_13_wuser_14_reg				(desc_13_wuser_14_reg[31:0]),
       .desc_13_wuser_15_reg				(desc_13_wuser_15_reg[31:0]),
       .desc_14_txn_type_reg				(desc_14_txn_type_reg[31:0]),
       .desc_14_size_reg					(desc_14_size_reg[31:0]),
       .desc_14_data_offset_reg			(desc_14_data_offset_reg[31:0]),
       .desc_14_data_host_addr_0_reg		(desc_14_data_host_addr_0_reg[31:0]),
       .desc_14_data_host_addr_1_reg		(desc_14_data_host_addr_1_reg[31:0]),
       .desc_14_data_host_addr_2_reg		(desc_14_data_host_addr_2_reg[31:0]),
       .desc_14_data_host_addr_3_reg		(desc_14_data_host_addr_3_reg[31:0]),
       .desc_14_wstrb_host_addr_0_reg	(desc_14_wstrb_host_addr_0_reg[31:0]),
       .desc_14_wstrb_host_addr_1_reg	(desc_14_wstrb_host_addr_1_reg[31:0]),
       .desc_14_wstrb_host_addr_2_reg	(desc_14_wstrb_host_addr_2_reg[31:0]),
       .desc_14_wstrb_host_addr_3_reg	(desc_14_wstrb_host_addr_3_reg[31:0]),
       .desc_14_axsize_reg				(desc_14_axsize_reg[31:0]),
       .desc_14_attr_reg					(desc_14_attr_reg[31:0]),
       .desc_14_axaddr_0_reg				(desc_14_axaddr_0_reg[31:0]),
       .desc_14_axaddr_1_reg				(desc_14_axaddr_1_reg[31:0]),
       .desc_14_axaddr_2_reg				(desc_14_axaddr_2_reg[31:0]),
       .desc_14_axaddr_3_reg				(desc_14_axaddr_3_reg[31:0]),
       .desc_14_axid_0_reg				(desc_14_axid_0_reg[31:0]),
       .desc_14_axid_1_reg				(desc_14_axid_1_reg[31:0]),
       .desc_14_axid_2_reg				(desc_14_axid_2_reg[31:0]),
       .desc_14_axid_3_reg				(desc_14_axid_3_reg[31:0]),
       .desc_14_axuser_0_reg				(desc_14_axuser_0_reg[31:0]),
       .desc_14_axuser_1_reg				(desc_14_axuser_1_reg[31:0]),
       .desc_14_axuser_2_reg				(desc_14_axuser_2_reg[31:0]),
       .desc_14_axuser_3_reg				(desc_14_axuser_3_reg[31:0]),
       .desc_14_axuser_4_reg				(desc_14_axuser_4_reg[31:0]),
       .desc_14_axuser_5_reg				(desc_14_axuser_5_reg[31:0]),
       .desc_14_axuser_6_reg				(desc_14_axuser_6_reg[31:0]),
       .desc_14_axuser_7_reg				(desc_14_axuser_7_reg[31:0]),
       .desc_14_axuser_8_reg				(desc_14_axuser_8_reg[31:0]),
       .desc_14_axuser_9_reg				(desc_14_axuser_9_reg[31:0]),
       .desc_14_axuser_10_reg			(desc_14_axuser_10_reg[31:0]),
       .desc_14_axuser_11_reg			(desc_14_axuser_11_reg[31:0]),
       .desc_14_axuser_12_reg			(desc_14_axuser_12_reg[31:0]),
       .desc_14_axuser_13_reg			(desc_14_axuser_13_reg[31:0]),
       .desc_14_axuser_14_reg			(desc_14_axuser_14_reg[31:0]),
       .desc_14_axuser_15_reg			(desc_14_axuser_15_reg[31:0]),
       .desc_14_xuser_0_reg				(desc_14_xuser_0_reg[31:0]),
       .desc_14_xuser_1_reg				(desc_14_xuser_1_reg[31:0]),
       .desc_14_xuser_2_reg				(desc_14_xuser_2_reg[31:0]),
       .desc_14_xuser_3_reg				(desc_14_xuser_3_reg[31:0]),
       .desc_14_xuser_4_reg				(desc_14_xuser_4_reg[31:0]),
       .desc_14_xuser_5_reg				(desc_14_xuser_5_reg[31:0]),
       .desc_14_xuser_6_reg				(desc_14_xuser_6_reg[31:0]),
       .desc_14_xuser_7_reg				(desc_14_xuser_7_reg[31:0]),
       .desc_14_xuser_8_reg				(desc_14_xuser_8_reg[31:0]),
       .desc_14_xuser_9_reg				(desc_14_xuser_9_reg[31:0]),
       .desc_14_xuser_10_reg				(desc_14_xuser_10_reg[31:0]),
       .desc_14_xuser_11_reg				(desc_14_xuser_11_reg[31:0]),
       .desc_14_xuser_12_reg				(desc_14_xuser_12_reg[31:0]),
       .desc_14_xuser_13_reg				(desc_14_xuser_13_reg[31:0]),
       .desc_14_xuser_14_reg				(desc_14_xuser_14_reg[31:0]),
       .desc_14_xuser_15_reg				(desc_14_xuser_15_reg[31:0]),
       .desc_14_wuser_0_reg				(desc_14_wuser_0_reg[31:0]),
       .desc_14_wuser_1_reg				(desc_14_wuser_1_reg[31:0]),
       .desc_14_wuser_2_reg				(desc_14_wuser_2_reg[31:0]),
       .desc_14_wuser_3_reg				(desc_14_wuser_3_reg[31:0]),
       .desc_14_wuser_4_reg				(desc_14_wuser_4_reg[31:0]),
       .desc_14_wuser_5_reg				(desc_14_wuser_5_reg[31:0]),
       .desc_14_wuser_6_reg				(desc_14_wuser_6_reg[31:0]),
       .desc_14_wuser_7_reg				(desc_14_wuser_7_reg[31:0]),
       .desc_14_wuser_8_reg				(desc_14_wuser_8_reg[31:0]),
       .desc_14_wuser_9_reg				(desc_14_wuser_9_reg[31:0]),
       .desc_14_wuser_10_reg				(desc_14_wuser_10_reg[31:0]),
       .desc_14_wuser_11_reg				(desc_14_wuser_11_reg[31:0]),
       .desc_14_wuser_12_reg				(desc_14_wuser_12_reg[31:0]),
       .desc_14_wuser_13_reg				(desc_14_wuser_13_reg[31:0]),
       .desc_14_wuser_14_reg				(desc_14_wuser_14_reg[31:0]),
       .desc_14_wuser_15_reg				(desc_14_wuser_15_reg[31:0]),
       .desc_15_txn_type_reg				(desc_15_txn_type_reg[31:0]),
       .desc_15_size_reg					(desc_15_size_reg[31:0]),
       .desc_15_data_offset_reg			(desc_15_data_offset_reg[31:0]),
       .desc_15_data_host_addr_0_reg		(desc_15_data_host_addr_0_reg[31:0]),
       .desc_15_data_host_addr_1_reg		(desc_15_data_host_addr_1_reg[31:0]),
       .desc_15_data_host_addr_2_reg		(desc_15_data_host_addr_2_reg[31:0]),
       .desc_15_data_host_addr_3_reg		(desc_15_data_host_addr_3_reg[31:0]),
       .desc_15_wstrb_host_addr_0_reg	(desc_15_wstrb_host_addr_0_reg[31:0]),
       .desc_15_wstrb_host_addr_1_reg	(desc_15_wstrb_host_addr_1_reg[31:0]),
       .desc_15_wstrb_host_addr_2_reg	(desc_15_wstrb_host_addr_2_reg[31:0]),
       .desc_15_wstrb_host_addr_3_reg	(desc_15_wstrb_host_addr_3_reg[31:0]),
       .desc_15_axsize_reg				(desc_15_axsize_reg[31:0]),
       .desc_15_attr_reg					(desc_15_attr_reg[31:0]),
       .desc_15_axaddr_0_reg				(desc_15_axaddr_0_reg[31:0]),
       .desc_15_axaddr_1_reg				(desc_15_axaddr_1_reg[31:0]),
       .desc_15_axaddr_2_reg				(desc_15_axaddr_2_reg[31:0]),
       .desc_15_axaddr_3_reg				(desc_15_axaddr_3_reg[31:0]),
       .desc_15_axid_0_reg				(desc_15_axid_0_reg[31:0]),
       .desc_15_axid_1_reg				(desc_15_axid_1_reg[31:0]),
       .desc_15_axid_2_reg				(desc_15_axid_2_reg[31:0]),
       .desc_15_axid_3_reg				(desc_15_axid_3_reg[31:0]),
       .desc_15_axuser_0_reg				(desc_15_axuser_0_reg[31:0]),
       .desc_15_axuser_1_reg				(desc_15_axuser_1_reg[31:0]),
       .desc_15_axuser_2_reg				(desc_15_axuser_2_reg[31:0]),
       .desc_15_axuser_3_reg				(desc_15_axuser_3_reg[31:0]),
       .desc_15_axuser_4_reg				(desc_15_axuser_4_reg[31:0]),
       .desc_15_axuser_5_reg				(desc_15_axuser_5_reg[31:0]),
       .desc_15_axuser_6_reg				(desc_15_axuser_6_reg[31:0]),
       .desc_15_axuser_7_reg				(desc_15_axuser_7_reg[31:0]),
       .desc_15_axuser_8_reg				(desc_15_axuser_8_reg[31:0]),
       .desc_15_axuser_9_reg				(desc_15_axuser_9_reg[31:0]),
       .desc_15_axuser_10_reg			(desc_15_axuser_10_reg[31:0]),
       .desc_15_axuser_11_reg			(desc_15_axuser_11_reg[31:0]),
       .desc_15_axuser_12_reg			(desc_15_axuser_12_reg[31:0]),
       .desc_15_axuser_13_reg			(desc_15_axuser_13_reg[31:0]),
       .desc_15_axuser_14_reg			(desc_15_axuser_14_reg[31:0]),
       .desc_15_axuser_15_reg			(desc_15_axuser_15_reg[31:0]),
       .desc_15_xuser_0_reg				(desc_15_xuser_0_reg[31:0]),
       .desc_15_xuser_1_reg				(desc_15_xuser_1_reg[31:0]),
       .desc_15_xuser_2_reg				(desc_15_xuser_2_reg[31:0]),
       .desc_15_xuser_3_reg				(desc_15_xuser_3_reg[31:0]),
       .desc_15_xuser_4_reg				(desc_15_xuser_4_reg[31:0]),
       .desc_15_xuser_5_reg				(desc_15_xuser_5_reg[31:0]),
       .desc_15_xuser_6_reg				(desc_15_xuser_6_reg[31:0]),
       .desc_15_xuser_7_reg				(desc_15_xuser_7_reg[31:0]),
       .desc_15_xuser_8_reg				(desc_15_xuser_8_reg[31:0]),
       .desc_15_xuser_9_reg				(desc_15_xuser_9_reg[31:0]),
       .desc_15_xuser_10_reg				(desc_15_xuser_10_reg[31:0]),
       .desc_15_xuser_11_reg				(desc_15_xuser_11_reg[31:0]),
       .desc_15_xuser_12_reg				(desc_15_xuser_12_reg[31:0]),
       .desc_15_xuser_13_reg				(desc_15_xuser_13_reg[31:0]),
       .desc_15_xuser_14_reg				(desc_15_xuser_14_reg[31:0]),
       .desc_15_xuser_15_reg				(desc_15_xuser_15_reg[31:0]),
       .desc_15_wuser_0_reg				(desc_15_wuser_0_reg[31:0]),
       .desc_15_wuser_1_reg				(desc_15_wuser_1_reg[31:0]),
       .desc_15_wuser_2_reg				(desc_15_wuser_2_reg[31:0]),
       .desc_15_wuser_3_reg				(desc_15_wuser_3_reg[31:0]),
       .desc_15_wuser_4_reg				(desc_15_wuser_4_reg[31:0]),
       .desc_15_wuser_5_reg				(desc_15_wuser_5_reg[31:0]),
       .desc_15_wuser_6_reg				(desc_15_wuser_6_reg[31:0]),
       .desc_15_wuser_7_reg				(desc_15_wuser_7_reg[31:0]),
       .desc_15_wuser_8_reg				(desc_15_wuser_8_reg[31:0]),
       .desc_15_wuser_9_reg				(desc_15_wuser_9_reg[31:0]),
       .desc_15_wuser_10_reg				(desc_15_wuser_10_reg[31:0]),
       .desc_15_wuser_11_reg				(desc_15_wuser_11_reg[31:0]),
       .desc_15_wuser_12_reg				(desc_15_wuser_12_reg[31:0]),
       .desc_15_wuser_13_reg				(desc_15_wuser_13_reg[31:0]),
       .desc_15_wuser_14_reg				(desc_15_wuser_14_reg[31:0]),
       .desc_15_wuser_15_reg				(desc_15_wuser_15_reg[31:0]),
       .m_axi_usr_awready				(m_axi_usr_awready),
       .m_axi_usr_wready					(m_axi_usr_wready),
       .m_axi_usr_bid					(m_axi_usr_bid[M_AXI_USR_ID_WIDTH-1:0]),
       .m_axi_usr_bresp					(m_axi_usr_bresp[1:0]),
       .m_axi_usr_buser					(m_axi_usr_buser ),
       .m_axi_usr_bvalid					(m_axi_usr_bvalid),
       .m_axi_usr_arready				(m_axi_usr_arready),
       .m_axi_usr_rid					(m_axi_usr_rid[M_AXI_USR_ID_WIDTH-1:0]),
       .m_axi_usr_rdata					(m_axi_usr_rdata[M_AXI_USR_DATA_WIDTH-1:0]),
       .m_axi_usr_rresp					(m_axi_usr_rresp[1:0]),
       .m_axi_usr_rlast					(m_axi_usr_rlast),
       .m_axi_usr_ruser					(m_axi_usr_ruser ),
       .m_axi_usr_rvalid					(m_axi_usr_rvalid));
   

endmodule // user_master_control




/* user_master_control.v ends here */
