/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *
 *
 */
,input [3:0] int_sn_desc_0_attr_acsnoop
 ,input [2:0] int_sn_desc_0_attr_acprot
 ,input [31:0] int_sn_desc_0_acaddr_0_addr
 ,input [31:0] int_sn_desc_0_acaddr_1_addr
 ,input [31:0] int_sn_desc_0_acaddr_2_addr
 ,input [31:0] int_sn_desc_0_acaddr_3_addr
 ,input [3:0] int_sn_desc_1_attr_acsnoop
 ,input [2:0] int_sn_desc_1_attr_acprot
 ,input [31:0] int_sn_desc_1_acaddr_0_addr
 ,input [31:0] int_sn_desc_1_acaddr_1_addr
 ,input [31:0] int_sn_desc_1_acaddr_2_addr
 ,input [31:0] int_sn_desc_1_acaddr_3_addr
 ,input [3:0] int_sn_desc_2_attr_acsnoop
 ,input [2:0] int_sn_desc_2_attr_acprot
 ,input [31:0] int_sn_desc_2_acaddr_0_addr
 ,input [31:0] int_sn_desc_2_acaddr_1_addr
 ,input [31:0] int_sn_desc_2_acaddr_2_addr
 ,input [31:0] int_sn_desc_2_acaddr_3_addr
 ,input [3:0] int_sn_desc_3_attr_acsnoop
 ,input [2:0] int_sn_desc_3_attr_acprot
 ,input [31:0] int_sn_desc_3_acaddr_0_addr
 ,input [31:0] int_sn_desc_3_acaddr_1_addr
 ,input [31:0] int_sn_desc_3_acaddr_2_addr
 ,input [31:0] int_sn_desc_3_acaddr_3_addr
 ,input [3:0] int_sn_desc_4_attr_acsnoop
 ,input [2:0] int_sn_desc_4_attr_acprot
 ,input [31:0] int_sn_desc_4_acaddr_0_addr
 ,input [31:0] int_sn_desc_4_acaddr_1_addr
 ,input [31:0] int_sn_desc_4_acaddr_2_addr
 ,input [31:0] int_sn_desc_4_acaddr_3_addr
 ,input [3:0] int_sn_desc_5_attr_acsnoop
 ,input [2:0] int_sn_desc_5_attr_acprot
 ,input [31:0] int_sn_desc_5_acaddr_0_addr
 ,input [31:0] int_sn_desc_5_acaddr_1_addr
 ,input [31:0] int_sn_desc_5_acaddr_2_addr
 ,input [31:0] int_sn_desc_5_acaddr_3_addr
 ,input [3:0] int_sn_desc_6_attr_acsnoop
 ,input [2:0] int_sn_desc_6_attr_acprot
 ,input [31:0] int_sn_desc_6_acaddr_0_addr
 ,input [31:0] int_sn_desc_6_acaddr_1_addr
 ,input [31:0] int_sn_desc_6_acaddr_2_addr
 ,input [31:0] int_sn_desc_6_acaddr_3_addr
 ,input [3:0] int_sn_desc_7_attr_acsnoop
 ,input [2:0] int_sn_desc_7_attr_acprot
 ,input [31:0] int_sn_desc_7_acaddr_0_addr
 ,input [31:0] int_sn_desc_7_acaddr_1_addr
 ,input [31:0] int_sn_desc_7_acaddr_2_addr
 ,input [31:0] int_sn_desc_7_acaddr_3_addr
