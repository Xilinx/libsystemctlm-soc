/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *   Wrapper around common rtl of AXI4, AXI4LITE and AXI3 rtl.
 *
 *
 */
`include "defines_common.vh"
module axi_slave_allprot    #(

                        parameter EN_INTFS_AXI4                  =  1, 
                        parameter EN_INTFS_AXI4LITE              =  0, 
                        parameter EN_INTFS_AXI3                  =  0, 
                        
                        parameter S_AXI_ADDR_WIDTH               = 64, 
                        parameter S_AXI_DATA_WIDTH               = 32, 
                        
                        parameter M_AXI_ADDR_WIDTH               = 64,    
                        parameter M_AXI_DATA_WIDTH               = 128, 
                        parameter M_AXI_ID_WIDTH                 = 16,  
                        parameter M_AXI_USER_WIDTH               = 32,    
                        
                        parameter S_AXI_USR_ADDR_WIDTH           = 64,    
                        parameter S_AXI_USR_DATA_WIDTH           = 128, 
                        parameter S_AXI_USR_ID_WIDTH             = 16,  
                        parameter S_AXI_USR_AWUSER_WIDTH         = 32,    
                        parameter S_AXI_USR_WUSER_WIDTH          = 32,    
                        parameter S_AXI_USR_BUSER_WIDTH          = 32,    
                        parameter S_AXI_USR_ARUSER_WIDTH         = 32,    
                        parameter S_AXI_USR_RUSER_WIDTH          = 32,    
                        
                        parameter RAM_SIZE                       = 16384, 
                        parameter MAX_DESC                       = 16,                   
                        parameter USR_RST_NUM                    = 4,
			parameter LAST_BRIDGE                    = 0,
			parameter EXTEND_WSTRB                   = 1,
                        parameter FORCE_RESP_ORDER               = 1
                        
                        )(
                          
                          //Clock and reset
                          input 								 axi_aclk, 
                          input 								 axi_aresetn, 
                          output [USR_RST_NUM-1:0] 				 usr_resetn,
                          //System Interrupt  
                          output 								 irq_out, 
                          input 								 irq_ack, 
                          //DUT Interrupt
                          output [127:0] 						 h2c_intr_out,
                          input [63:0] 							 c2h_intr_in,
                          //DUT GPIO
                          input [255:0] 						 c2h_gpio_in,
                          output [255:0] 						 h2c_gpio_out,
                          
                          // S_AXI - AXI4-Lite
                          input wire [S_AXI_ADDR_WIDTH-1:0] 	 s_axi_awaddr,
                          input wire [2:0] 						 s_axi_awprot,
                          input wire 							 s_axi_awvalid,
                          output wire 							 s_axi_awready,
                          input wire [S_AXI_DATA_WIDTH-1:0] 	 s_axi_wdata,
                          input wire [(S_AXI_DATA_WIDTH/8)-1:0]  s_axi_wstrb,
                          input wire 							 s_axi_wvalid,
                          output wire 							 s_axi_wready,
                          output wire [1:0] 					 s_axi_bresp,
                          output wire 							 s_axi_bvalid,
                          input wire 							 s_axi_bready,
                          input wire [S_AXI_ADDR_WIDTH-1:0] 	 s_axi_araddr,
                          input wire [2:0] 						 s_axi_arprot,
                          input wire 							 s_axi_arvalid,
                          output wire 							 s_axi_arready,
                          output wire [S_AXI_DATA_WIDTH-1:0] 	 s_axi_rdata,
                          output wire [1:0] 					 s_axi_rresp,
                          output wire 							 s_axi_rvalid,
                          input wire 							 s_axi_rready, 

                          // M_AXI - AXI4
                          output wire [M_AXI_ID_WIDTH-1 : 0] 	 m_axi_awid,
                          output wire [M_AXI_ADDR_WIDTH-1 : 0] 	 m_axi_awaddr,
                          output wire [7 : 0] 					 m_axi_awlen,
                          output wire [2 : 0] 					 m_axi_awsize,
                          output wire [1 : 0] 					 m_axi_awburst,
                          output wire 							 m_axi_awlock,
                          output wire [3 : 0] 					 m_axi_awcache,
                          output wire [2 : 0] 					 m_axi_awprot,
                          output wire [3 : 0] 					 m_axi_awqos,
                          output wire [3:0] 					 m_axi_awregion, 
                          output wire [M_AXI_USER_WIDTH-1 : 0] 	 m_axi_awuser,
                          output wire 							 m_axi_awvalid,
                          input wire 							 m_axi_awready,
                          output wire [M_AXI_DATA_WIDTH-1 : 0] 	 m_axi_wdata,
                          output wire [M_AXI_DATA_WIDTH/8-1 : 0] m_axi_wstrb,
                          output wire 							 m_axi_wlast,
                          output wire [M_AXI_USER_WIDTH-1 : 0] 	 m_axi_wuser,
                          output wire 							 m_axi_wvalid,
                          input wire 							 m_axi_wready,
                          input wire [M_AXI_ID_WIDTH-1 : 0] 	 m_axi_bid,
                          input wire [1 : 0] 					 m_axi_bresp,
                          input wire [M_AXI_USER_WIDTH-1 : 0] 	 m_axi_buser,
                          input wire 							 m_axi_bvalid,
                          output wire 							 m_axi_bready,
                          output wire [M_AXI_ID_WIDTH-1 : 0] 	 m_axi_arid,
                          output wire [M_AXI_ADDR_WIDTH-1 : 0] 	 m_axi_araddr,
                          output wire [7 : 0] 					 m_axi_arlen,
                          output wire [2 : 0] 					 m_axi_arsize,
                          output wire [1 : 0] 					 m_axi_arburst,
                          output wire 							 m_axi_arlock,
                          output wire [3 : 0] 					 m_axi_arcache,
                          output wire [2 : 0] 					 m_axi_arprot,
                          output wire [3 : 0] 					 m_axi_arqos,
                          output wire [3:0] 					 m_axi_arregion, 
                          output wire [M_AXI_USER_WIDTH-1 : 0] 	 m_axi_aruser,
                          output wire 							 m_axi_arvalid,
                          input wire 							 m_axi_arready,
                          input wire [M_AXI_ID_WIDTH-1 : 0] 	 m_axi_rid,
                          input wire [M_AXI_DATA_WIDTH-1 : 0] 	 m_axi_rdata,
                          input wire [1 : 0] 					 m_axi_rresp,
                          input wire 							 m_axi_rlast,
                          input wire [M_AXI_USER_WIDTH-1 : 0] 	 m_axi_ruser,
                          input wire 							 m_axi_rvalid,
                          output wire 							 m_axi_rready,

                          //S_AXI_USR
                          input [S_AXI_USR_ID_WIDTH-1:0] 		 s_axi_usr_awid, 
                          input [S_AXI_USR_ADDR_WIDTH-1:0] 		 s_axi_usr_awaddr, 
                          input [7:0] 							 s_axi_usr_awlen, 
                          input [2:0] 							 s_axi_usr_awsize, 
                          input [1:0] 							 s_axi_usr_awburst, 
                          input [1:0] 							 s_axi_usr_awlock, 
                          input [3:0] 							 s_axi_usr_awcache, 
                          input [2:0] 							 s_axi_usr_awprot, 
                          input [3:0] 							 s_axi_usr_awqos, 
                          input [3:0] 							 s_axi_usr_awregion, 
                          input [S_AXI_USR_AWUSER_WIDTH-1:0] 	 s_axi_usr_awuser, 
                          input 								 s_axi_usr_awvalid, 
                          output 								 s_axi_usr_awready, 
                          input [S_AXI_USR_DATA_WIDTH-1:0] 		 s_axi_usr_wdata, 
                          input [(S_AXI_USR_DATA_WIDTH/8)-1:0] 	 s_axi_usr_wstrb, 
                          input 								 s_axi_usr_wlast, 
                          input [S_AXI_USR_ID_WIDTH-1:0] 		 s_axi_usr_wid, 
                          input [S_AXI_USR_WUSER_WIDTH-1:0] 	 s_axi_usr_wuser, 
                          input 								 s_axi_usr_wvalid, 
                          output 								 s_axi_usr_wready, 
                          output [S_AXI_USR_ID_WIDTH-1:0] 		 s_axi_usr_bid, 
                          output [1:0] 							 s_axi_usr_bresp, 
                          output [S_AXI_USR_BUSER_WIDTH-1:0] 	 s_axi_usr_buser, 
                          output 								 s_axi_usr_bvalid, 
                          input 								 s_axi_usr_bready, 
                          input [S_AXI_USR_ID_WIDTH-1:0] 		 s_axi_usr_arid, 
                          input [S_AXI_USR_ADDR_WIDTH-1:0] 		 s_axi_usr_araddr, 
                          input [7:0] 							 s_axi_usr_arlen, 
                          input [2:0] 							 s_axi_usr_arsize, 
                          input [1:0] 							 s_axi_usr_arburst, 
                          input [1:0] 							 s_axi_usr_arlock, 
                          input [3:0] 							 s_axi_usr_arcache, 
                          input [2:0] 							 s_axi_usr_arprot, 
                          input [3:0] 							 s_axi_usr_arqos, 
                          input [3:0] 							 s_axi_usr_arregion, 
                          input [S_AXI_USR_ARUSER_WIDTH-1:0] 	 s_axi_usr_aruser, 
                          input 								 s_axi_usr_arvalid, 
                          output 								 s_axi_usr_arready, 
                          output [S_AXI_USR_ID_WIDTH-1:0] 		 s_axi_usr_rid, 
                          output [S_AXI_USR_DATA_WIDTH-1:0] 	 s_axi_usr_rdata, 
                          output [1:0] 							 s_axi_usr_rresp, 
                          output 								 s_axi_usr_rlast, 
                          output [S_AXI_USR_RUSER_WIDTH-1:0] 	 s_axi_usr_ruser, 
                          output 								 s_axi_usr_rvalid, 
                          input 								 s_axi_usr_rready 
  
                          );



wire                                                               rst_n;
wire [31:0]                                                        reset_reg;              
genvar                                                             gi;
 
   

assign rst_n = axi_aresetn & reset_reg[0];

generate 
for (gi=0; gi<=USR_RST_NUM-1; gi=gi+1) begin: gen_AW_fifo_valid
  assign usr_resetn[gi] = axi_aresetn & reset_reg[gi+1];
end
endgenerate




/*AUTOWIRE*/   
// Beginning of automatic wires (for undeclared instantiated-module outputs)
wire [31:0]             addr_in_0_reg;          
wire [31:0]             addr_in_1_reg;          
wire [31:0]             addr_in_2_reg;          
wire [31:0]             addr_in_3_reg;          
wire [31:0]             axi_bridge_config_reg;  
wire [31:0]             axi_max_desc_reg;       
wire [31:0]             bridge_type_reg;        
wire [31:0] 			c2h_gpio_0_reg;  
wire [31:0] 			c2h_gpio_10_reg; 
wire [31:0] 			c2h_gpio_11_reg; 
wire [31:0] 			c2h_gpio_12_reg; 
wire [31:0] 			c2h_gpio_13_reg; 
wire [31:0] 			c2h_gpio_14_reg; 
wire [31:0] 			c2h_gpio_15_reg; 
wire [31:0] 			c2h_gpio_1_reg;  
wire [31:0] 			c2h_gpio_2_reg;  
wire [31:0] 			c2h_gpio_3_reg;  
wire [31:0] 			c2h_gpio_4_reg;  
wire [31:0] 			c2h_gpio_5_reg;  
wire [31:0] 			c2h_gpio_6_reg;  
wire [31:0] 			c2h_gpio_7_reg;  
wire [31:0] 			c2h_gpio_8_reg;  
wire [31:0] 			c2h_gpio_9_reg;
wire [31:0] 			h2c_gpio_1_reg;  
wire [31:0] 			h2c_gpio_2_reg;  
wire [31:0] 			h2c_gpio_3_reg;  
wire [31:0] 			h2c_gpio_4_reg;  
wire [31:0] 			h2c_gpio_5_reg;  
wire [31:0] 			h2c_gpio_6_reg;  
wire [31:0] 			h2c_gpio_7_reg;  
wire [31:0] 			h2c_gpio_0_reg;  
wire [31:0]             desc_0_attr_reg;        
wire [31:0]             desc_0_axaddr_0_reg;    
wire [31:0]             desc_0_axaddr_1_reg;    
wire [31:0]             desc_0_axaddr_2_reg;    
wire [31:0]             desc_0_axaddr_3_reg;    
wire [31:0]             desc_0_axid_0_reg;      
wire [31:0]             desc_0_axid_1_reg;      
wire [31:0]             desc_0_axid_2_reg;      
wire [31:0]             desc_0_axid_3_reg;      
wire [31:0]             desc_0_axsize_reg;      
wire [31:0]             desc_0_axuser_0_reg;    
wire [31:0]             desc_0_axuser_10_reg;   
wire [31:0]             desc_0_axuser_11_reg;   
wire [31:0]             desc_0_axuser_12_reg;   
wire [31:0]             desc_0_axuser_13_reg;   
wire [31:0]             desc_0_axuser_14_reg;   
wire [31:0]             desc_0_axuser_15_reg;   
wire [31:0]             desc_0_axuser_1_reg;    
wire [31:0]             desc_0_axuser_2_reg;    
wire [31:0]             desc_0_axuser_3_reg;    
wire [31:0]             desc_0_axuser_4_reg;    
wire [31:0]             desc_0_axuser_5_reg;    
wire [31:0]             desc_0_axuser_6_reg;    
wire [31:0]             desc_0_axuser_7_reg;    
wire [31:0]             desc_0_axuser_8_reg;    
wire [31:0]             desc_0_axuser_9_reg;    
wire [31:0]             desc_0_data_host_addr_0_reg;
wire [31:0]             desc_0_data_host_addr_1_reg;
wire [31:0]             desc_0_data_host_addr_2_reg;
wire [31:0]             desc_0_data_host_addr_3_reg;
wire [31:0]             desc_0_data_offset_reg; 
wire [31:0]             desc_0_size_reg;        
wire [31:0]             desc_0_txn_type_reg;    
wire [31:0]             desc_0_wstrb_host_addr_0_reg;
wire [31:0]             desc_0_wstrb_host_addr_1_reg;
wire [31:0]             desc_0_wstrb_host_addr_2_reg;
wire [31:0]             desc_0_wstrb_host_addr_3_reg;
wire [31:0]             desc_0_wuser_0_reg;     
wire [31:0]             desc_0_wuser_10_reg;    
wire [31:0]             desc_0_wuser_11_reg;    
wire [31:0]             desc_0_wuser_12_reg;    
wire [31:0]             desc_0_wuser_13_reg;    
wire [31:0]             desc_0_wuser_14_reg;    
wire [31:0]             desc_0_wuser_15_reg;    
wire [31:0]             desc_0_wuser_1_reg;     
wire [31:0]             desc_0_wuser_2_reg;     
wire [31:0]             desc_0_wuser_3_reg;     
wire [31:0]             desc_0_wuser_4_reg;     
wire [31:0]             desc_0_wuser_5_reg;     
wire [31:0]             desc_0_wuser_6_reg;     
wire [31:0]             desc_0_wuser_7_reg;     
wire [31:0]             desc_0_wuser_8_reg;     
wire [31:0]             desc_0_wuser_9_reg;     
wire [31:0]             desc_0_xuser_0_reg;     
wire [31:0]             desc_0_xuser_10_reg;    
wire [31:0]             desc_0_xuser_11_reg;    
wire [31:0]             desc_0_xuser_12_reg;    
wire [31:0]             desc_0_xuser_13_reg;    
wire [31:0]             desc_0_xuser_14_reg;    
wire [31:0]             desc_0_xuser_15_reg;    
wire [31:0]             desc_0_xuser_1_reg;     
wire [31:0]             desc_0_xuser_2_reg;     
wire [31:0]             desc_0_xuser_3_reg;     
wire [31:0]             desc_0_xuser_4_reg;     
wire [31:0]             desc_0_xuser_5_reg;     
wire [31:0]             desc_0_xuser_6_reg;     
wire [31:0]             desc_0_xuser_7_reg;     
wire [31:0]             desc_0_xuser_8_reg;     
wire [31:0]             desc_0_xuser_9_reg;     
wire [31:0]             desc_10_attr_reg;       
wire [31:0]             desc_10_axaddr_0_reg;   
wire [31:0]             desc_10_axaddr_1_reg;   
wire [31:0]             desc_10_axaddr_2_reg;   
wire [31:0]             desc_10_axaddr_3_reg;   
wire [31:0]             desc_10_axid_0_reg;     
wire [31:0]             desc_10_axid_1_reg;     
wire [31:0]             desc_10_axid_2_reg;     
wire [31:0]             desc_10_axid_3_reg;     
wire [31:0]             desc_10_axsize_reg;     
wire [31:0]             desc_10_axuser_0_reg;   
wire [31:0]             desc_10_axuser_10_reg;  
wire [31:0]             desc_10_axuser_11_reg;  
wire [31:0]             desc_10_axuser_12_reg;  
wire [31:0]             desc_10_axuser_13_reg;  
wire [31:0]             desc_10_axuser_14_reg;  
wire [31:0]             desc_10_axuser_15_reg;  
wire [31:0]             desc_10_axuser_1_reg;   
wire [31:0]             desc_10_axuser_2_reg;   
wire [31:0]             desc_10_axuser_3_reg;   
wire [31:0]             desc_10_axuser_4_reg;   
wire [31:0]             desc_10_axuser_5_reg;   
wire [31:0]             desc_10_axuser_6_reg;   
wire [31:0]             desc_10_axuser_7_reg;   
wire [31:0]             desc_10_axuser_8_reg;   
wire [31:0]             desc_10_axuser_9_reg;   
wire [31:0]             desc_10_data_host_addr_0_reg;
wire [31:0]             desc_10_data_host_addr_1_reg;
wire [31:0]             desc_10_data_host_addr_2_reg;
wire [31:0]             desc_10_data_host_addr_3_reg;
wire [31:0]             desc_10_data_offset_reg;
wire [31:0]             desc_10_size_reg;       
wire [31:0]             desc_10_txn_type_reg;   
wire [31:0]             desc_10_wstrb_host_addr_0_reg;
wire [31:0]             desc_10_wstrb_host_addr_1_reg;
wire [31:0]             desc_10_wstrb_host_addr_2_reg;
wire [31:0]             desc_10_wstrb_host_addr_3_reg;
wire [31:0]             desc_10_wuser_0_reg;    
wire [31:0]             desc_10_wuser_10_reg;   
wire [31:0]             desc_10_wuser_11_reg;   
wire [31:0]             desc_10_wuser_12_reg;   
wire [31:0]             desc_10_wuser_13_reg;   
wire [31:0]             desc_10_wuser_14_reg;   
wire [31:0]             desc_10_wuser_15_reg;   
wire [31:0]             desc_10_wuser_1_reg;    
wire [31:0]             desc_10_wuser_2_reg;    
wire [31:0]             desc_10_wuser_3_reg;    
wire [31:0]             desc_10_wuser_4_reg;    
wire [31:0]             desc_10_wuser_5_reg;    
wire [31:0]             desc_10_wuser_6_reg;    
wire [31:0]             desc_10_wuser_7_reg;    
wire [31:0]             desc_10_wuser_8_reg;    
wire [31:0]             desc_10_wuser_9_reg;    
wire [31:0]             desc_10_xuser_0_reg;    
wire [31:0]             desc_10_xuser_10_reg;   
wire [31:0]             desc_10_xuser_11_reg;   
wire [31:0]             desc_10_xuser_12_reg;   
wire [31:0]             desc_10_xuser_13_reg;   
wire [31:0]             desc_10_xuser_14_reg;   
wire [31:0]             desc_10_xuser_15_reg;   
wire [31:0]             desc_10_xuser_1_reg;    
wire [31:0]             desc_10_xuser_2_reg;    
wire [31:0]             desc_10_xuser_3_reg;    
wire [31:0]             desc_10_xuser_4_reg;    
wire [31:0]             desc_10_xuser_5_reg;    
wire [31:0]             desc_10_xuser_6_reg;    
wire [31:0]             desc_10_xuser_7_reg;    
wire [31:0]             desc_10_xuser_8_reg;    
wire [31:0]             desc_10_xuser_9_reg;    
wire [31:0]             desc_11_attr_reg;       
wire [31:0]             desc_11_axaddr_0_reg;   
wire [31:0]             desc_11_axaddr_1_reg;   
wire [31:0]             desc_11_axaddr_2_reg;   
wire [31:0]             desc_11_axaddr_3_reg;   
wire [31:0]             desc_11_axid_0_reg;     
wire [31:0]             desc_11_axid_1_reg;     
wire [31:0]             desc_11_axid_2_reg;     
wire [31:0]             desc_11_axid_3_reg;     
wire [31:0]             desc_11_axsize_reg;     
wire [31:0]             desc_11_axuser_0_reg;   
wire [31:0]             desc_11_axuser_10_reg;  
wire [31:0]             desc_11_axuser_11_reg;  
wire [31:0]             desc_11_axuser_12_reg;  
wire [31:0]             desc_11_axuser_13_reg;  
wire [31:0]             desc_11_axuser_14_reg;  
wire [31:0]             desc_11_axuser_15_reg;  
wire [31:0]             desc_11_axuser_1_reg;   
wire [31:0]             desc_11_axuser_2_reg;   
wire [31:0]             desc_11_axuser_3_reg;   
wire [31:0]             desc_11_axuser_4_reg;   
wire [31:0]             desc_11_axuser_5_reg;   
wire [31:0]             desc_11_axuser_6_reg;   
wire [31:0]             desc_11_axuser_7_reg;   
wire [31:0]             desc_11_axuser_8_reg;   
wire [31:0]             desc_11_axuser_9_reg;   
wire [31:0]             desc_11_data_host_addr_0_reg;
wire [31:0]             desc_11_data_host_addr_1_reg;
wire [31:0]             desc_11_data_host_addr_2_reg;
wire [31:0]             desc_11_data_host_addr_3_reg;
wire [31:0]             desc_11_data_offset_reg;
wire [31:0]             desc_11_size_reg;       
wire [31:0]             desc_11_txn_type_reg;   
wire [31:0]             desc_11_wstrb_host_addr_0_reg;
wire [31:0]             desc_11_wstrb_host_addr_1_reg;
wire [31:0]             desc_11_wstrb_host_addr_2_reg;
wire [31:0]             desc_11_wstrb_host_addr_3_reg;
wire [31:0]             desc_11_wuser_0_reg;    
wire [31:0]             desc_11_wuser_10_reg;   
wire [31:0]             desc_11_wuser_11_reg;   
wire [31:0]             desc_11_wuser_12_reg;   
wire [31:0]             desc_11_wuser_13_reg;   
wire [31:0]             desc_11_wuser_14_reg;   
wire [31:0]             desc_11_wuser_15_reg;   
wire [31:0]             desc_11_wuser_1_reg;    
wire [31:0]             desc_11_wuser_2_reg;    
wire [31:0]             desc_11_wuser_3_reg;    
wire [31:0]             desc_11_wuser_4_reg;    
wire [31:0]             desc_11_wuser_5_reg;    
wire [31:0]             desc_11_wuser_6_reg;    
wire [31:0]             desc_11_wuser_7_reg;    
wire [31:0]             desc_11_wuser_8_reg;    
wire [31:0]             desc_11_wuser_9_reg;    
wire [31:0]             desc_11_xuser_0_reg;    
wire [31:0]             desc_11_xuser_10_reg;   
wire [31:0]             desc_11_xuser_11_reg;   
wire [31:0]             desc_11_xuser_12_reg;   
wire [31:0]             desc_11_xuser_13_reg;   
wire [31:0]             desc_11_xuser_14_reg;   
wire [31:0]             desc_11_xuser_15_reg;   
wire [31:0]             desc_11_xuser_1_reg;    
wire [31:0]             desc_11_xuser_2_reg;    
wire [31:0]             desc_11_xuser_3_reg;    
wire [31:0]             desc_11_xuser_4_reg;    
wire [31:0]             desc_11_xuser_5_reg;    
wire [31:0]             desc_11_xuser_6_reg;    
wire [31:0]             desc_11_xuser_7_reg;    
wire [31:0]             desc_11_xuser_8_reg;    
wire [31:0]             desc_11_xuser_9_reg;    
wire [31:0]             desc_12_attr_reg;       
wire [31:0]             desc_12_axaddr_0_reg;   
wire [31:0]             desc_12_axaddr_1_reg;   
wire [31:0]             desc_12_axaddr_2_reg;   
wire [31:0]             desc_12_axaddr_3_reg;   
wire [31:0]             desc_12_axid_0_reg;     
wire [31:0]             desc_12_axid_1_reg;     
wire [31:0]             desc_12_axid_2_reg;     
wire [31:0]             desc_12_axid_3_reg;     
wire [31:0]             desc_12_axsize_reg;     
wire [31:0]             desc_12_axuser_0_reg;   
wire [31:0]             desc_12_axuser_10_reg;  
wire [31:0]             desc_12_axuser_11_reg;  
wire [31:0]             desc_12_axuser_12_reg;  
wire [31:0]             desc_12_axuser_13_reg;  
wire [31:0]             desc_12_axuser_14_reg;  
wire [31:0]             desc_12_axuser_15_reg;  
wire [31:0]             desc_12_axuser_1_reg;   
wire [31:0]             desc_12_axuser_2_reg;   
wire [31:0]             desc_12_axuser_3_reg;   
wire [31:0]             desc_12_axuser_4_reg;   
wire [31:0]             desc_12_axuser_5_reg;   
wire [31:0]             desc_12_axuser_6_reg;   
wire [31:0]             desc_12_axuser_7_reg;   
wire [31:0]             desc_12_axuser_8_reg;   
wire [31:0]             desc_12_axuser_9_reg;   
wire [31:0]             desc_12_data_host_addr_0_reg;
wire [31:0]             desc_12_data_host_addr_1_reg;
wire [31:0]             desc_12_data_host_addr_2_reg;
wire [31:0]             desc_12_data_host_addr_3_reg;
wire [31:0]             desc_12_data_offset_reg;
wire [31:0]             desc_12_size_reg;       
wire [31:0]             desc_12_txn_type_reg;   
wire [31:0]             desc_12_wstrb_host_addr_0_reg;
wire [31:0]             desc_12_wstrb_host_addr_1_reg;
wire [31:0]             desc_12_wstrb_host_addr_2_reg;
wire [31:0]             desc_12_wstrb_host_addr_3_reg;
wire [31:0]             desc_12_wuser_0_reg;    
wire [31:0]             desc_12_wuser_10_reg;   
wire [31:0]             desc_12_wuser_11_reg;   
wire [31:0]             desc_12_wuser_12_reg;   
wire [31:0]             desc_12_wuser_13_reg;   
wire [31:0]             desc_12_wuser_14_reg;   
wire [31:0]             desc_12_wuser_15_reg;   
wire [31:0]             desc_12_wuser_1_reg;    
wire [31:0]             desc_12_wuser_2_reg;    
wire [31:0]             desc_12_wuser_3_reg;    
wire [31:0]             desc_12_wuser_4_reg;    
wire [31:0]             desc_12_wuser_5_reg;    
wire [31:0]             desc_12_wuser_6_reg;    
wire [31:0]             desc_12_wuser_7_reg;    
wire [31:0]             desc_12_wuser_8_reg;    
wire [31:0]             desc_12_wuser_9_reg;    
wire [31:0]             desc_12_xuser_0_reg;    
wire [31:0]             desc_12_xuser_10_reg;   
wire [31:0]             desc_12_xuser_11_reg;   
wire [31:0]             desc_12_xuser_12_reg;   
wire [31:0]             desc_12_xuser_13_reg;   
wire [31:0]             desc_12_xuser_14_reg;   
wire [31:0]             desc_12_xuser_15_reg;   
wire [31:0]             desc_12_xuser_1_reg;    
wire [31:0]             desc_12_xuser_2_reg;    
wire [31:0]             desc_12_xuser_3_reg;    
wire [31:0]             desc_12_xuser_4_reg;    
wire [31:0]             desc_12_xuser_5_reg;    
wire [31:0]             desc_12_xuser_6_reg;    
wire [31:0]             desc_12_xuser_7_reg;    
wire [31:0]             desc_12_xuser_8_reg;    
wire [31:0]             desc_12_xuser_9_reg;    
wire [31:0]             desc_13_attr_reg;       
wire [31:0]             desc_13_axaddr_0_reg;   
wire [31:0]             desc_13_axaddr_1_reg;   
wire [31:0]             desc_13_axaddr_2_reg;   
wire [31:0]             desc_13_axaddr_3_reg;   
wire [31:0]             desc_13_axid_0_reg;     
wire [31:0]             desc_13_axid_1_reg;     
wire [31:0]             desc_13_axid_2_reg;     
wire [31:0]             desc_13_axid_3_reg;     
wire [31:0]             desc_13_axsize_reg;     
wire [31:0]             desc_13_axuser_0_reg;   
wire [31:0]             desc_13_axuser_10_reg;  
wire [31:0]             desc_13_axuser_11_reg;  
wire [31:0]             desc_13_axuser_12_reg;  
wire [31:0]             desc_13_axuser_13_reg;  
wire [31:0]             desc_13_axuser_14_reg;  
wire [31:0]             desc_13_axuser_15_reg;  
wire [31:0]             desc_13_axuser_1_reg;   
wire [31:0]             desc_13_axuser_2_reg;   
wire [31:0]             desc_13_axuser_3_reg;   
wire [31:0]             desc_13_axuser_4_reg;   
wire [31:0]             desc_13_axuser_5_reg;   
wire [31:0]             desc_13_axuser_6_reg;   
wire [31:0]             desc_13_axuser_7_reg;   
wire [31:0]             desc_13_axuser_8_reg;   
wire [31:0]             desc_13_axuser_9_reg;   
wire [31:0]             desc_13_data_host_addr_0_reg;
wire [31:0]             desc_13_data_host_addr_1_reg;
wire [31:0]             desc_13_data_host_addr_2_reg;
wire [31:0]             desc_13_data_host_addr_3_reg;
wire [31:0]             desc_13_data_offset_reg;
wire [31:0]             desc_13_size_reg;       
wire [31:0]             desc_13_txn_type_reg;   
wire [31:0]             desc_13_wstrb_host_addr_0_reg;
wire [31:0]             desc_13_wstrb_host_addr_1_reg;
wire [31:0]             desc_13_wstrb_host_addr_2_reg;
wire [31:0]             desc_13_wstrb_host_addr_3_reg;
wire [31:0]             desc_13_wuser_0_reg;    
wire [31:0]             desc_13_wuser_10_reg;   
wire [31:0]             desc_13_wuser_11_reg;   
wire [31:0]             desc_13_wuser_12_reg;   
wire [31:0]             desc_13_wuser_13_reg;   
wire [31:0]             desc_13_wuser_14_reg;   
wire [31:0]             desc_13_wuser_15_reg;   
wire [31:0]             desc_13_wuser_1_reg;    
wire [31:0]             desc_13_wuser_2_reg;    
wire [31:0]             desc_13_wuser_3_reg;    
wire [31:0]             desc_13_wuser_4_reg;    
wire [31:0]             desc_13_wuser_5_reg;    
wire [31:0]             desc_13_wuser_6_reg;    
wire [31:0]             desc_13_wuser_7_reg;    
wire [31:0]             desc_13_wuser_8_reg;    
wire [31:0]             desc_13_wuser_9_reg;    
wire [31:0]             desc_13_xuser_0_reg;    
wire [31:0]             desc_13_xuser_10_reg;   
wire [31:0]             desc_13_xuser_11_reg;   
wire [31:0]             desc_13_xuser_12_reg;   
wire [31:0]             desc_13_xuser_13_reg;   
wire [31:0]             desc_13_xuser_14_reg;   
wire [31:0]             desc_13_xuser_15_reg;   
wire [31:0]             desc_13_xuser_1_reg;    
wire [31:0]             desc_13_xuser_2_reg;    
wire [31:0]             desc_13_xuser_3_reg;    
wire [31:0]             desc_13_xuser_4_reg;    
wire [31:0]             desc_13_xuser_5_reg;    
wire [31:0]             desc_13_xuser_6_reg;    
wire [31:0]             desc_13_xuser_7_reg;    
wire [31:0]             desc_13_xuser_8_reg;    
wire [31:0]             desc_13_xuser_9_reg;    
wire [31:0]             desc_14_attr_reg;       
wire [31:0]             desc_14_axaddr_0_reg;   
wire [31:0]             desc_14_axaddr_1_reg;   
wire [31:0]             desc_14_axaddr_2_reg;   
wire [31:0]             desc_14_axaddr_3_reg;   
wire [31:0]             desc_14_axid_0_reg;     
wire [31:0]             desc_14_axid_1_reg;     
wire [31:0]             desc_14_axid_2_reg;     
wire [31:0]             desc_14_axid_3_reg;     
wire [31:0]             desc_14_axsize_reg;     
wire [31:0]             desc_14_axuser_0_reg;   
wire [31:0]             desc_14_axuser_10_reg;  
wire [31:0]             desc_14_axuser_11_reg;  
wire [31:0]             desc_14_axuser_12_reg;  
wire [31:0]             desc_14_axuser_13_reg;  
wire [31:0]             desc_14_axuser_14_reg;  
wire [31:0]             desc_14_axuser_15_reg;  
wire [31:0]             desc_14_axuser_1_reg;   
wire [31:0]             desc_14_axuser_2_reg;   
wire [31:0]             desc_14_axuser_3_reg;   
wire [31:0]             desc_14_axuser_4_reg;   
wire [31:0]             desc_14_axuser_5_reg;   
wire [31:0]             desc_14_axuser_6_reg;   
wire [31:0]             desc_14_axuser_7_reg;   
wire [31:0]             desc_14_axuser_8_reg;   
wire [31:0]             desc_14_axuser_9_reg;   
wire [31:0]             desc_14_data_host_addr_0_reg;
wire [31:0]             desc_14_data_host_addr_1_reg;
wire [31:0]             desc_14_data_host_addr_2_reg;
wire [31:0]             desc_14_data_host_addr_3_reg;
wire [31:0]             desc_14_data_offset_reg;
wire [31:0]             desc_14_size_reg;       
wire [31:0]             desc_14_txn_type_reg;   
wire [31:0]             desc_14_wstrb_host_addr_0_reg;
wire [31:0]             desc_14_wstrb_host_addr_1_reg;
wire [31:0]             desc_14_wstrb_host_addr_2_reg;
wire [31:0]             desc_14_wstrb_host_addr_3_reg;
wire [31:0]             desc_14_wuser_0_reg;    
wire [31:0]             desc_14_wuser_10_reg;   
wire [31:0]             desc_14_wuser_11_reg;   
wire [31:0]             desc_14_wuser_12_reg;   
wire [31:0]             desc_14_wuser_13_reg;   
wire [31:0]             desc_14_wuser_14_reg;   
wire [31:0]             desc_14_wuser_15_reg;   
wire [31:0]             desc_14_wuser_1_reg;    
wire [31:0]             desc_14_wuser_2_reg;    
wire [31:0]             desc_14_wuser_3_reg;    
wire [31:0]             desc_14_wuser_4_reg;    
wire [31:0]             desc_14_wuser_5_reg;    
wire [31:0]             desc_14_wuser_6_reg;    
wire [31:0]             desc_14_wuser_7_reg;    
wire [31:0]             desc_14_wuser_8_reg;    
wire [31:0]             desc_14_wuser_9_reg;    
wire [31:0]             desc_14_xuser_0_reg;    
wire [31:0]             desc_14_xuser_10_reg;   
wire [31:0]             desc_14_xuser_11_reg;   
wire [31:0]             desc_14_xuser_12_reg;   
wire [31:0]             desc_14_xuser_13_reg;   
wire [31:0]             desc_14_xuser_14_reg;   
wire [31:0]             desc_14_xuser_15_reg;   
wire [31:0]             desc_14_xuser_1_reg;    
wire [31:0]             desc_14_xuser_2_reg;    
wire [31:0]             desc_14_xuser_3_reg;    
wire [31:0]             desc_14_xuser_4_reg;    
wire [31:0]             desc_14_xuser_5_reg;    
wire [31:0]             desc_14_xuser_6_reg;    
wire [31:0]             desc_14_xuser_7_reg;    
wire [31:0]             desc_14_xuser_8_reg;    
wire [31:0]             desc_14_xuser_9_reg;    
wire [31:0]             desc_15_attr_reg;       
wire [31:0]             desc_15_axaddr_0_reg;   
wire [31:0]             desc_15_axaddr_1_reg;   
wire [31:0]             desc_15_axaddr_2_reg;   
wire [31:0]             desc_15_axaddr_3_reg;   
wire [31:0]             desc_15_axid_0_reg;     
wire [31:0]             desc_15_axid_1_reg;     
wire [31:0]             desc_15_axid_2_reg;     
wire [31:0]             desc_15_axid_3_reg;     
wire [31:0]             desc_15_axsize_reg;     
wire [31:0]             desc_15_axuser_0_reg;   
wire [31:0]             desc_15_axuser_10_reg;  
wire [31:0]             desc_15_axuser_11_reg;  
wire [31:0]             desc_15_axuser_12_reg;  
wire [31:0]             desc_15_axuser_13_reg;  
wire [31:0]             desc_15_axuser_14_reg;  
wire [31:0]             desc_15_axuser_15_reg;  
wire [31:0]             desc_15_axuser_1_reg;   
wire [31:0]             desc_15_axuser_2_reg;   
wire [31:0]             desc_15_axuser_3_reg;   
wire [31:0]             desc_15_axuser_4_reg;   
wire [31:0]             desc_15_axuser_5_reg;   
wire [31:0]             desc_15_axuser_6_reg;   
wire [31:0]             desc_15_axuser_7_reg;   
wire [31:0]             desc_15_axuser_8_reg;   
wire [31:0]             desc_15_axuser_9_reg;   
wire [31:0]             desc_15_data_host_addr_0_reg;
wire [31:0]             desc_15_data_host_addr_1_reg;
wire [31:0]             desc_15_data_host_addr_2_reg;
wire [31:0]             desc_15_data_host_addr_3_reg;
wire [31:0]             desc_15_data_offset_reg;
wire [31:0]             desc_15_size_reg;       
wire [31:0]             desc_15_txn_type_reg;   
wire [31:0]             desc_15_wstrb_host_addr_0_reg;
wire [31:0]             desc_15_wstrb_host_addr_1_reg;
wire [31:0]             desc_15_wstrb_host_addr_2_reg;
wire [31:0]             desc_15_wstrb_host_addr_3_reg;
wire [31:0]             desc_15_wuser_0_reg;    
wire [31:0]             desc_15_wuser_10_reg;   
wire [31:0]             desc_15_wuser_11_reg;   
wire [31:0]             desc_15_wuser_12_reg;   
wire [31:0]             desc_15_wuser_13_reg;   
wire [31:0]             desc_15_wuser_14_reg;   
wire [31:0]             desc_15_wuser_15_reg;   
wire [31:0]             desc_15_wuser_1_reg;    
wire [31:0]             desc_15_wuser_2_reg;    
wire [31:0]             desc_15_wuser_3_reg;    
wire [31:0]             desc_15_wuser_4_reg;    
wire [31:0]             desc_15_wuser_5_reg;    
wire [31:0]             desc_15_wuser_6_reg;    
wire [31:0]             desc_15_wuser_7_reg;    
wire [31:0]             desc_15_wuser_8_reg;    
wire [31:0]             desc_15_wuser_9_reg;    
wire [31:0]             desc_15_xuser_0_reg;    
wire [31:0]             desc_15_xuser_10_reg;   
wire [31:0]             desc_15_xuser_11_reg;   
wire [31:0]             desc_15_xuser_12_reg;   
wire [31:0]             desc_15_xuser_13_reg;   
wire [31:0]             desc_15_xuser_14_reg;   
wire [31:0]             desc_15_xuser_15_reg;   
wire [31:0]             desc_15_xuser_1_reg;    
wire [31:0]             desc_15_xuser_2_reg;    
wire [31:0]             desc_15_xuser_3_reg;    
wire [31:0]             desc_15_xuser_4_reg;    
wire [31:0]             desc_15_xuser_5_reg;    
wire [31:0]             desc_15_xuser_6_reg;    
wire [31:0]             desc_15_xuser_7_reg;    
wire [31:0]             desc_15_xuser_8_reg;    
wire [31:0]             desc_15_xuser_9_reg;    
wire [31:0]             desc_1_attr_reg;        
wire [31:0]             desc_1_axaddr_0_reg;    
wire [31:0]             desc_1_axaddr_1_reg;    
wire [31:0]             desc_1_axaddr_2_reg;    
wire [31:0]             desc_1_axaddr_3_reg;    
wire [31:0]             desc_1_axid_0_reg;      
wire [31:0]             desc_1_axid_1_reg;      
wire [31:0]             desc_1_axid_2_reg;      
wire [31:0]             desc_1_axid_3_reg;      
wire [31:0]             desc_1_axsize_reg;      
wire [31:0]             desc_1_axuser_0_reg;    
wire [31:0]             desc_1_axuser_10_reg;   
wire [31:0]             desc_1_axuser_11_reg;   
wire [31:0]             desc_1_axuser_12_reg;   
wire [31:0]             desc_1_axuser_13_reg;   
wire [31:0]             desc_1_axuser_14_reg;   
wire [31:0]             desc_1_axuser_15_reg;   
wire [31:0]             desc_1_axuser_1_reg;    
wire [31:0]             desc_1_axuser_2_reg;    
wire [31:0]             desc_1_axuser_3_reg;    
wire [31:0]             desc_1_axuser_4_reg;    
wire [31:0]             desc_1_axuser_5_reg;    
wire [31:0]             desc_1_axuser_6_reg;    
wire [31:0]             desc_1_axuser_7_reg;    
wire [31:0]             desc_1_axuser_8_reg;    
wire [31:0]             desc_1_axuser_9_reg;    
wire [31:0]             desc_1_data_host_addr_0_reg;
wire [31:0]             desc_1_data_host_addr_1_reg;
wire [31:0]             desc_1_data_host_addr_2_reg;
wire [31:0]             desc_1_data_host_addr_3_reg;
wire [31:0]             desc_1_data_offset_reg; 
wire [31:0]             desc_1_size_reg;        
wire [31:0]             desc_1_txn_type_reg;    
wire [31:0]             desc_1_wstrb_host_addr_0_reg;
wire [31:0]             desc_1_wstrb_host_addr_1_reg;
wire [31:0]             desc_1_wstrb_host_addr_2_reg;
wire [31:0]             desc_1_wstrb_host_addr_3_reg;
wire [31:0]             desc_1_wuser_0_reg;     
wire [31:0]             desc_1_wuser_10_reg;    
wire [31:0]             desc_1_wuser_11_reg;    
wire [31:0]             desc_1_wuser_12_reg;    
wire [31:0]             desc_1_wuser_13_reg;    
wire [31:0]             desc_1_wuser_14_reg;    
wire [31:0]             desc_1_wuser_15_reg;    
wire [31:0]             desc_1_wuser_1_reg;     
wire [31:0]             desc_1_wuser_2_reg;     
wire [31:0]             desc_1_wuser_3_reg;     
wire [31:0]             desc_1_wuser_4_reg;     
wire [31:0]             desc_1_wuser_5_reg;     
wire [31:0]             desc_1_wuser_6_reg;     
wire [31:0]             desc_1_wuser_7_reg;     
wire [31:0]             desc_1_wuser_8_reg;     
wire [31:0]             desc_1_wuser_9_reg;     
wire [31:0]             desc_1_xuser_0_reg;     
wire [31:0]             desc_1_xuser_10_reg;    
wire [31:0]             desc_1_xuser_11_reg;    
wire [31:0]             desc_1_xuser_12_reg;    
wire [31:0]             desc_1_xuser_13_reg;    
wire [31:0]             desc_1_xuser_14_reg;    
wire [31:0]             desc_1_xuser_15_reg;    
wire [31:0]             desc_1_xuser_1_reg;     
wire [31:0]             desc_1_xuser_2_reg;     
wire [31:0]             desc_1_xuser_3_reg;     
wire [31:0]             desc_1_xuser_4_reg;     
wire [31:0]             desc_1_xuser_5_reg;     
wire [31:0]             desc_1_xuser_6_reg;     
wire [31:0]             desc_1_xuser_7_reg;     
wire [31:0]             desc_1_xuser_8_reg;     
wire [31:0]             desc_1_xuser_9_reg;     
wire [31:0]             desc_2_attr_reg;        
wire [31:0]             desc_2_axaddr_0_reg;    
wire [31:0]             desc_2_axaddr_1_reg;    
wire [31:0]             desc_2_axaddr_2_reg;    
wire [31:0]             desc_2_axaddr_3_reg;    
wire [31:0]             desc_2_axid_0_reg;      
wire [31:0]             desc_2_axid_1_reg;      
wire [31:0]             desc_2_axid_2_reg;      
wire [31:0]             desc_2_axid_3_reg;      
wire [31:0]             desc_2_axsize_reg;      
wire [31:0]             desc_2_axuser_0_reg;    
wire [31:0]             desc_2_axuser_10_reg;   
wire [31:0]             desc_2_axuser_11_reg;   
wire [31:0]             desc_2_axuser_12_reg;   
wire [31:0]             desc_2_axuser_13_reg;   
wire [31:0]             desc_2_axuser_14_reg;   
wire [31:0]             desc_2_axuser_15_reg;   
wire [31:0]             desc_2_axuser_1_reg;    
wire [31:0]             desc_2_axuser_2_reg;    
wire [31:0]             desc_2_axuser_3_reg;    
wire [31:0]             desc_2_axuser_4_reg;    
wire [31:0]             desc_2_axuser_5_reg;    
wire [31:0]             desc_2_axuser_6_reg;    
wire [31:0]             desc_2_axuser_7_reg;    
wire [31:0]             desc_2_axuser_8_reg;    
wire [31:0]             desc_2_axuser_9_reg;    
wire [31:0]             desc_2_data_host_addr_0_reg;
wire [31:0]             desc_2_data_host_addr_1_reg;
wire [31:0]             desc_2_data_host_addr_2_reg;
wire [31:0]             desc_2_data_host_addr_3_reg;
wire [31:0]             desc_2_data_offset_reg; 
wire [31:0]             desc_2_size_reg;        
wire [31:0]             desc_2_txn_type_reg;    
wire [31:0]             desc_2_wstrb_host_addr_0_reg;
wire [31:0]             desc_2_wstrb_host_addr_1_reg;
wire [31:0]             desc_2_wstrb_host_addr_2_reg;
wire [31:0]             desc_2_wstrb_host_addr_3_reg;
wire [31:0]             desc_2_wuser_0_reg;     
wire [31:0]             desc_2_wuser_10_reg;    
wire [31:0]             desc_2_wuser_11_reg;    
wire [31:0]             desc_2_wuser_12_reg;    
wire [31:0]             desc_2_wuser_13_reg;    
wire [31:0]             desc_2_wuser_14_reg;    
wire [31:0]             desc_2_wuser_15_reg;    
wire [31:0]             desc_2_wuser_1_reg;     
wire [31:0]             desc_2_wuser_2_reg;     
wire [31:0]             desc_2_wuser_3_reg;     
wire [31:0]             desc_2_wuser_4_reg;     
wire [31:0]             desc_2_wuser_5_reg;     
wire [31:0]             desc_2_wuser_6_reg;     
wire [31:0]             desc_2_wuser_7_reg;     
wire [31:0]             desc_2_wuser_8_reg;     
wire [31:0]             desc_2_wuser_9_reg;     
wire [31:0]             desc_2_xuser_0_reg;     
wire [31:0]             desc_2_xuser_10_reg;    
wire [31:0]             desc_2_xuser_11_reg;    
wire [31:0]             desc_2_xuser_12_reg;    
wire [31:0]             desc_2_xuser_13_reg;    
wire [31:0]             desc_2_xuser_14_reg;    
wire [31:0]             desc_2_xuser_15_reg;    
wire [31:0]             desc_2_xuser_1_reg;     
wire [31:0]             desc_2_xuser_2_reg;     
wire [31:0]             desc_2_xuser_3_reg;     
wire [31:0]             desc_2_xuser_4_reg;     
wire [31:0]             desc_2_xuser_5_reg;     
wire [31:0]             desc_2_xuser_6_reg;     
wire [31:0]             desc_2_xuser_7_reg;     
wire [31:0]             desc_2_xuser_8_reg;     
wire [31:0]             desc_2_xuser_9_reg;     
wire [31:0]             desc_3_attr_reg;        
wire [31:0]             desc_3_axaddr_0_reg;    
wire [31:0]             desc_3_axaddr_1_reg;    
wire [31:0]             desc_3_axaddr_2_reg;    
wire [31:0]             desc_3_axaddr_3_reg;    
wire [31:0]             desc_3_axid_0_reg;      
wire [31:0]             desc_3_axid_1_reg;      
wire [31:0]             desc_3_axid_2_reg;      
wire [31:0]             desc_3_axid_3_reg;      
wire [31:0]             desc_3_axsize_reg;      
wire [31:0]             desc_3_axuser_0_reg;    
wire [31:0]             desc_3_axuser_10_reg;   
wire [31:0]             desc_3_axuser_11_reg;   
wire [31:0]             desc_3_axuser_12_reg;   
wire [31:0]             desc_3_axuser_13_reg;   
wire [31:0]             desc_3_axuser_14_reg;   
wire [31:0]             desc_3_axuser_15_reg;   
wire [31:0]             desc_3_axuser_1_reg;    
wire [31:0]             desc_3_axuser_2_reg;    
wire [31:0]             desc_3_axuser_3_reg;    
wire [31:0]             desc_3_axuser_4_reg;    
wire [31:0]             desc_3_axuser_5_reg;    
wire [31:0]             desc_3_axuser_6_reg;    
wire [31:0]             desc_3_axuser_7_reg;    
wire [31:0]             desc_3_axuser_8_reg;    
wire [31:0]             desc_3_axuser_9_reg;    
wire [31:0]             desc_3_data_host_addr_0_reg;
wire [31:0]             desc_3_data_host_addr_1_reg;
wire [31:0]             desc_3_data_host_addr_2_reg;
wire [31:0]             desc_3_data_host_addr_3_reg;
wire [31:0]             desc_3_data_offset_reg; 
wire [31:0]             desc_3_size_reg;        
wire [31:0]             desc_3_txn_type_reg;    
wire [31:0]             desc_3_wstrb_host_addr_0_reg;
wire [31:0]             desc_3_wstrb_host_addr_1_reg;
wire [31:0]             desc_3_wstrb_host_addr_2_reg;
wire [31:0]             desc_3_wstrb_host_addr_3_reg;
wire [31:0]             desc_3_wuser_0_reg;     
wire [31:0]             desc_3_wuser_10_reg;    
wire [31:0]             desc_3_wuser_11_reg;    
wire [31:0]             desc_3_wuser_12_reg;    
wire [31:0]             desc_3_wuser_13_reg;    
wire [31:0]             desc_3_wuser_14_reg;    
wire [31:0]             desc_3_wuser_15_reg;    
wire [31:0]             desc_3_wuser_1_reg;     
wire [31:0]             desc_3_wuser_2_reg;     
wire [31:0]             desc_3_wuser_3_reg;     
wire [31:0]             desc_3_wuser_4_reg;     
wire [31:0]             desc_3_wuser_5_reg;     
wire [31:0]             desc_3_wuser_6_reg;     
wire [31:0]             desc_3_wuser_7_reg;     
wire [31:0]             desc_3_wuser_8_reg;     
wire [31:0]             desc_3_wuser_9_reg;     
wire [31:0]             desc_3_xuser_0_reg;     
wire [31:0]             desc_3_xuser_10_reg;    
wire [31:0]             desc_3_xuser_11_reg;    
wire [31:0]             desc_3_xuser_12_reg;    
wire [31:0]             desc_3_xuser_13_reg;    
wire [31:0]             desc_3_xuser_14_reg;    
wire [31:0]             desc_3_xuser_15_reg;    
wire [31:0]             desc_3_xuser_1_reg;     
wire [31:0]             desc_3_xuser_2_reg;     
wire [31:0]             desc_3_xuser_3_reg;     
wire [31:0]             desc_3_xuser_4_reg;     
wire [31:0]             desc_3_xuser_5_reg;     
wire [31:0]             desc_3_xuser_6_reg;     
wire [31:0]             desc_3_xuser_7_reg;     
wire [31:0]             desc_3_xuser_8_reg;     
wire [31:0]             desc_3_xuser_9_reg;     
wire [31:0]             desc_4_attr_reg;        
wire [31:0]             desc_4_axaddr_0_reg;    
wire [31:0]             desc_4_axaddr_1_reg;    
wire [31:0]             desc_4_axaddr_2_reg;    
wire [31:0]             desc_4_axaddr_3_reg;    
wire [31:0]             desc_4_axid_0_reg;      
wire [31:0]             desc_4_axid_1_reg;      
wire [31:0]             desc_4_axid_2_reg;      
wire [31:0]             desc_4_axid_3_reg;      
wire [31:0]             desc_4_axsize_reg;      
wire [31:0]             desc_4_axuser_0_reg;    
wire [31:0]             desc_4_axuser_10_reg;   
wire [31:0]             desc_4_axuser_11_reg;   
wire [31:0]             desc_4_axuser_12_reg;   
wire [31:0]             desc_4_axuser_13_reg;   
wire [31:0]             desc_4_axuser_14_reg;   
wire [31:0]             desc_4_axuser_15_reg;   
wire [31:0]             desc_4_axuser_1_reg;    
wire [31:0]             desc_4_axuser_2_reg;    
wire [31:0]             desc_4_axuser_3_reg;    
wire [31:0]             desc_4_axuser_4_reg;    
wire [31:0]             desc_4_axuser_5_reg;    
wire [31:0]             desc_4_axuser_6_reg;    
wire [31:0]             desc_4_axuser_7_reg;    
wire [31:0]             desc_4_axuser_8_reg;    
wire [31:0]             desc_4_axuser_9_reg;    
wire [31:0]             desc_4_data_host_addr_0_reg;
wire [31:0]             desc_4_data_host_addr_1_reg;
wire [31:0]             desc_4_data_host_addr_2_reg;
wire [31:0]             desc_4_data_host_addr_3_reg;
wire [31:0]             desc_4_data_offset_reg; 
wire [31:0]             desc_4_size_reg;        
wire [31:0]             desc_4_txn_type_reg;    
wire [31:0]             desc_4_wstrb_host_addr_0_reg;
wire [31:0]             desc_4_wstrb_host_addr_1_reg;
wire [31:0]             desc_4_wstrb_host_addr_2_reg;
wire [31:0]             desc_4_wstrb_host_addr_3_reg;
wire [31:0]             desc_4_wuser_0_reg;     
wire [31:0]             desc_4_wuser_10_reg;    
wire [31:0]             desc_4_wuser_11_reg;    
wire [31:0]             desc_4_wuser_12_reg;    
wire [31:0]             desc_4_wuser_13_reg;    
wire [31:0]             desc_4_wuser_14_reg;    
wire [31:0]             desc_4_wuser_15_reg;    
wire [31:0]             desc_4_wuser_1_reg;     
wire [31:0]             desc_4_wuser_2_reg;     
wire [31:0]             desc_4_wuser_3_reg;     
wire [31:0]             desc_4_wuser_4_reg;     
wire [31:0]             desc_4_wuser_5_reg;     
wire [31:0]             desc_4_wuser_6_reg;     
wire [31:0]             desc_4_wuser_7_reg;     
wire [31:0]             desc_4_wuser_8_reg;     
wire [31:0]             desc_4_wuser_9_reg;     
wire [31:0]             desc_4_xuser_0_reg;     
wire [31:0]             desc_4_xuser_10_reg;    
wire [31:0]             desc_4_xuser_11_reg;    
wire [31:0]             desc_4_xuser_12_reg;    
wire [31:0]             desc_4_xuser_13_reg;    
wire [31:0]             desc_4_xuser_14_reg;    
wire [31:0]             desc_4_xuser_15_reg;    
wire [31:0]             desc_4_xuser_1_reg;     
wire [31:0]             desc_4_xuser_2_reg;     
wire [31:0]             desc_4_xuser_3_reg;     
wire [31:0]             desc_4_xuser_4_reg;     
wire [31:0]             desc_4_xuser_5_reg;     
wire [31:0]             desc_4_xuser_6_reg;     
wire [31:0]             desc_4_xuser_7_reg;     
wire [31:0]             desc_4_xuser_8_reg;     
wire [31:0]             desc_4_xuser_9_reg;     
wire [31:0]             desc_5_attr_reg;        
wire [31:0]             desc_5_axaddr_0_reg;    
wire [31:0]             desc_5_axaddr_1_reg;    
wire [31:0]             desc_5_axaddr_2_reg;    
wire [31:0]             desc_5_axaddr_3_reg;    
wire [31:0]             desc_5_axid_0_reg;      
wire [31:0]             desc_5_axid_1_reg;      
wire [31:0]             desc_5_axid_2_reg;      
wire [31:0]             desc_5_axid_3_reg;      
wire [31:0]             desc_5_axsize_reg;      
wire [31:0]             desc_5_axuser_0_reg;    
wire [31:0]             desc_5_axuser_10_reg;   
wire [31:0]             desc_5_axuser_11_reg;   
wire [31:0]             desc_5_axuser_12_reg;   
wire [31:0]             desc_5_axuser_13_reg;   
wire [31:0]             desc_5_axuser_14_reg;   
wire [31:0]             desc_5_axuser_15_reg;   
wire [31:0]             desc_5_axuser_1_reg;    
wire [31:0]             desc_5_axuser_2_reg;    
wire [31:0]             desc_5_axuser_3_reg;    
wire [31:0]             desc_5_axuser_4_reg;    
wire [31:0]             desc_5_axuser_5_reg;    
wire [31:0]             desc_5_axuser_6_reg;    
wire [31:0]             desc_5_axuser_7_reg;    
wire [31:0]             desc_5_axuser_8_reg;    
wire [31:0]             desc_5_axuser_9_reg;    
wire [31:0]             desc_5_data_host_addr_0_reg;
wire [31:0]             desc_5_data_host_addr_1_reg;
wire [31:0]             desc_5_data_host_addr_2_reg;
wire [31:0]             desc_5_data_host_addr_3_reg;
wire [31:0]             desc_5_data_offset_reg; 
wire [31:0]             desc_5_size_reg;        
wire [31:0]             desc_5_txn_type_reg;    
wire [31:0]             desc_5_wstrb_host_addr_0_reg;
wire [31:0]             desc_5_wstrb_host_addr_1_reg;
wire [31:0]             desc_5_wstrb_host_addr_2_reg;
wire [31:0]             desc_5_wstrb_host_addr_3_reg;
wire [31:0]             desc_5_wuser_0_reg;     
wire [31:0]             desc_5_wuser_10_reg;    
wire [31:0]             desc_5_wuser_11_reg;    
wire [31:0]             desc_5_wuser_12_reg;    
wire [31:0]             desc_5_wuser_13_reg;    
wire [31:0]             desc_5_wuser_14_reg;    
wire [31:0]             desc_5_wuser_15_reg;    
wire [31:0]             desc_5_wuser_1_reg;     
wire [31:0]             desc_5_wuser_2_reg;     
wire [31:0]             desc_5_wuser_3_reg;     
wire [31:0]             desc_5_wuser_4_reg;     
wire [31:0]             desc_5_wuser_5_reg;     
wire [31:0]             desc_5_wuser_6_reg;     
wire [31:0]             desc_5_wuser_7_reg;     
wire [31:0]             desc_5_wuser_8_reg;     
wire [31:0]             desc_5_wuser_9_reg;     
wire [31:0]             desc_5_xuser_0_reg;     
wire [31:0]             desc_5_xuser_10_reg;    
wire [31:0]             desc_5_xuser_11_reg;    
wire [31:0]             desc_5_xuser_12_reg;    
wire [31:0]             desc_5_xuser_13_reg;    
wire [31:0]             desc_5_xuser_14_reg;    
wire [31:0]             desc_5_xuser_15_reg;    
wire [31:0]             desc_5_xuser_1_reg;     
wire [31:0]             desc_5_xuser_2_reg;     
wire [31:0]             desc_5_xuser_3_reg;     
wire [31:0]             desc_5_xuser_4_reg;     
wire [31:0]             desc_5_xuser_5_reg;     
wire [31:0]             desc_5_xuser_6_reg;     
wire [31:0]             desc_5_xuser_7_reg;     
wire [31:0]             desc_5_xuser_8_reg;     
wire [31:0]             desc_5_xuser_9_reg;     
wire [31:0]             desc_6_attr_reg;        
wire [31:0]             desc_6_axaddr_0_reg;    
wire [31:0]             desc_6_axaddr_1_reg;    
wire [31:0]             desc_6_axaddr_2_reg;    
wire [31:0]             desc_6_axaddr_3_reg;    
wire [31:0]             desc_6_axid_0_reg;      
wire [31:0]             desc_6_axid_1_reg;      
wire [31:0]             desc_6_axid_2_reg;      
wire [31:0]             desc_6_axid_3_reg;      
wire [31:0]             desc_6_axsize_reg;      
wire [31:0]             desc_6_axuser_0_reg;    
wire [31:0]             desc_6_axuser_10_reg;   
wire [31:0]             desc_6_axuser_11_reg;   
wire [31:0]             desc_6_axuser_12_reg;   
wire [31:0]             desc_6_axuser_13_reg;   
wire [31:0]             desc_6_axuser_14_reg;   
wire [31:0]             desc_6_axuser_15_reg;   
wire [31:0]             desc_6_axuser_1_reg;    
wire [31:0]             desc_6_axuser_2_reg;    
wire [31:0]             desc_6_axuser_3_reg;    
wire [31:0]             desc_6_axuser_4_reg;    
wire [31:0]             desc_6_axuser_5_reg;    
wire [31:0]             desc_6_axuser_6_reg;    
wire [31:0]             desc_6_axuser_7_reg;    
wire [31:0]             desc_6_axuser_8_reg;    
wire [31:0]             desc_6_axuser_9_reg;    
wire [31:0]             desc_6_data_host_addr_0_reg;
wire [31:0]             desc_6_data_host_addr_1_reg;
wire [31:0]             desc_6_data_host_addr_2_reg;
wire [31:0]             desc_6_data_host_addr_3_reg;
wire [31:0]             desc_6_data_offset_reg; 
wire [31:0]             desc_6_size_reg;        
wire [31:0]             desc_6_txn_type_reg;    
wire [31:0]             desc_6_wstrb_host_addr_0_reg;
wire [31:0]             desc_6_wstrb_host_addr_1_reg;
wire [31:0]             desc_6_wstrb_host_addr_2_reg;
wire [31:0]             desc_6_wstrb_host_addr_3_reg;
wire [31:0]             desc_6_wuser_0_reg;     
wire [31:0]             desc_6_wuser_10_reg;    
wire [31:0]             desc_6_wuser_11_reg;    
wire [31:0]             desc_6_wuser_12_reg;    
wire [31:0]             desc_6_wuser_13_reg;    
wire [31:0]             desc_6_wuser_14_reg;    
wire [31:0]             desc_6_wuser_15_reg;    
wire [31:0]             desc_6_wuser_1_reg;     
wire [31:0]             desc_6_wuser_2_reg;     
wire [31:0]             desc_6_wuser_3_reg;     
wire [31:0]             desc_6_wuser_4_reg;     
wire [31:0]             desc_6_wuser_5_reg;     
wire [31:0]             desc_6_wuser_6_reg;     
wire [31:0]             desc_6_wuser_7_reg;     
wire [31:0]             desc_6_wuser_8_reg;     
wire [31:0]             desc_6_wuser_9_reg;     
wire [31:0]             desc_6_xuser_0_reg;     
wire [31:0]             desc_6_xuser_10_reg;    
wire [31:0]             desc_6_xuser_11_reg;    
wire [31:0]             desc_6_xuser_12_reg;    
wire [31:0]             desc_6_xuser_13_reg;    
wire [31:0]             desc_6_xuser_14_reg;    
wire [31:0]             desc_6_xuser_15_reg;    
wire [31:0]             desc_6_xuser_1_reg;     
wire [31:0]             desc_6_xuser_2_reg;     
wire [31:0]             desc_6_xuser_3_reg;     
wire [31:0]             desc_6_xuser_4_reg;     
wire [31:0]             desc_6_xuser_5_reg;     
wire [31:0]             desc_6_xuser_6_reg;     
wire [31:0]             desc_6_xuser_7_reg;     
wire [31:0]             desc_6_xuser_8_reg;     
wire [31:0]             desc_6_xuser_9_reg;     
wire [31:0]             desc_7_attr_reg;        
wire [31:0]             desc_7_axaddr_0_reg;    
wire [31:0]             desc_7_axaddr_1_reg;    
wire [31:0]             desc_7_axaddr_2_reg;    
wire [31:0]             desc_7_axaddr_3_reg;    
wire [31:0]             desc_7_axid_0_reg;      
wire [31:0]             desc_7_axid_1_reg;      
wire [31:0]             desc_7_axid_2_reg;      
wire [31:0]             desc_7_axid_3_reg;      
wire [31:0]             desc_7_axsize_reg;      
wire [31:0]             desc_7_axuser_0_reg;    
wire [31:0]             desc_7_axuser_10_reg;   
wire [31:0]             desc_7_axuser_11_reg;   
wire [31:0]             desc_7_axuser_12_reg;   
wire [31:0]             desc_7_axuser_13_reg;   
wire [31:0]             desc_7_axuser_14_reg;   
wire [31:0]             desc_7_axuser_15_reg;   
wire [31:0]             desc_7_axuser_1_reg;    
wire [31:0]             desc_7_axuser_2_reg;    
wire [31:0]             desc_7_axuser_3_reg;    
wire [31:0]             desc_7_axuser_4_reg;    
wire [31:0]             desc_7_axuser_5_reg;    
wire [31:0]             desc_7_axuser_6_reg;    
wire [31:0]             desc_7_axuser_7_reg;    
wire [31:0]             desc_7_axuser_8_reg;    
wire [31:0]             desc_7_axuser_9_reg;    
wire [31:0]             desc_7_data_host_addr_0_reg;
wire [31:0]             desc_7_data_host_addr_1_reg;
wire [31:0]             desc_7_data_host_addr_2_reg;
wire [31:0]             desc_7_data_host_addr_3_reg;
wire [31:0]             desc_7_data_offset_reg; 
wire [31:0]             desc_7_size_reg;        
wire [31:0]             desc_7_txn_type_reg;    
wire [31:0]             desc_7_wstrb_host_addr_0_reg;
wire [31:0]             desc_7_wstrb_host_addr_1_reg;
wire [31:0]             desc_7_wstrb_host_addr_2_reg;
wire [31:0]             desc_7_wstrb_host_addr_3_reg;
wire [31:0]             desc_7_wuser_0_reg;     
wire [31:0]             desc_7_wuser_10_reg;    
wire [31:0]             desc_7_wuser_11_reg;    
wire [31:0]             desc_7_wuser_12_reg;    
wire [31:0]             desc_7_wuser_13_reg;    
wire [31:0]             desc_7_wuser_14_reg;    
wire [31:0]             desc_7_wuser_15_reg;    
wire [31:0]             desc_7_wuser_1_reg;     
wire [31:0]             desc_7_wuser_2_reg;     
wire [31:0]             desc_7_wuser_3_reg;     
wire [31:0]             desc_7_wuser_4_reg;     
wire [31:0]             desc_7_wuser_5_reg;     
wire [31:0]             desc_7_wuser_6_reg;     
wire [31:0]             desc_7_wuser_7_reg;     
wire [31:0]             desc_7_wuser_8_reg;     
wire [31:0]             desc_7_wuser_9_reg;     
wire [31:0]             desc_7_xuser_0_reg;     
wire [31:0]             desc_7_xuser_10_reg;    
wire [31:0]             desc_7_xuser_11_reg;    
wire [31:0]             desc_7_xuser_12_reg;    
wire [31:0]             desc_7_xuser_13_reg;    
wire [31:0]             desc_7_xuser_14_reg;    
wire [31:0]             desc_7_xuser_15_reg;    
wire [31:0]             desc_7_xuser_1_reg;     
wire [31:0]             desc_7_xuser_2_reg;     
wire [31:0]             desc_7_xuser_3_reg;     
wire [31:0]             desc_7_xuser_4_reg;     
wire [31:0]             desc_7_xuser_5_reg;     
wire [31:0]             desc_7_xuser_6_reg;     
wire [31:0]             desc_7_xuser_7_reg;     
wire [31:0]             desc_7_xuser_8_reg;     
wire [31:0]             desc_7_xuser_9_reg;     
wire [31:0]             desc_8_attr_reg;        
wire [31:0]             desc_8_axaddr_0_reg;    
wire [31:0]             desc_8_axaddr_1_reg;    
wire [31:0]             desc_8_axaddr_2_reg;    
wire [31:0]             desc_8_axaddr_3_reg;    
wire [31:0]             desc_8_axid_0_reg;      
wire [31:0]             desc_8_axid_1_reg;      
wire [31:0]             desc_8_axid_2_reg;      
wire [31:0]             desc_8_axid_3_reg;      
wire [31:0]             desc_8_axsize_reg;      
wire [31:0]             desc_8_axuser_0_reg;    
wire [31:0]             desc_8_axuser_10_reg;   
wire [31:0]             desc_8_axuser_11_reg;   
wire [31:0]             desc_8_axuser_12_reg;   
wire [31:0]             desc_8_axuser_13_reg;   
wire [31:0]             desc_8_axuser_14_reg;   
wire [31:0]             desc_8_axuser_15_reg;   
wire [31:0]             desc_8_axuser_1_reg;    
wire [31:0]             desc_8_axuser_2_reg;    
wire [31:0]             desc_8_axuser_3_reg;    
wire [31:0]             desc_8_axuser_4_reg;    
wire [31:0]             desc_8_axuser_5_reg;    
wire [31:0]             desc_8_axuser_6_reg;    
wire [31:0]             desc_8_axuser_7_reg;    
wire [31:0]             desc_8_axuser_8_reg;    
wire [31:0]             desc_8_axuser_9_reg;    
wire [31:0]             desc_8_data_host_addr_0_reg;
wire [31:0]             desc_8_data_host_addr_1_reg;
wire [31:0]             desc_8_data_host_addr_2_reg;
wire [31:0]             desc_8_data_host_addr_3_reg;
wire [31:0]             desc_8_data_offset_reg; 
wire [31:0]             desc_8_size_reg;        
wire [31:0]             desc_8_txn_type_reg;    
wire [31:0]             desc_8_wstrb_host_addr_0_reg;
wire [31:0]             desc_8_wstrb_host_addr_1_reg;
wire [31:0]             desc_8_wstrb_host_addr_2_reg;
wire [31:0]             desc_8_wstrb_host_addr_3_reg;
wire [31:0]             desc_8_wuser_0_reg;     
wire [31:0]             desc_8_wuser_10_reg;    
wire [31:0]             desc_8_wuser_11_reg;    
wire [31:0]             desc_8_wuser_12_reg;    
wire [31:0]             desc_8_wuser_13_reg;    
wire [31:0]             desc_8_wuser_14_reg;    
wire [31:0]             desc_8_wuser_15_reg;    
wire [31:0]             desc_8_wuser_1_reg;     
wire [31:0]             desc_8_wuser_2_reg;     
wire [31:0]             desc_8_wuser_3_reg;     
wire [31:0]             desc_8_wuser_4_reg;     
wire [31:0]             desc_8_wuser_5_reg;     
wire [31:0]             desc_8_wuser_6_reg;     
wire [31:0]             desc_8_wuser_7_reg;     
wire [31:0]             desc_8_wuser_8_reg;     
wire [31:0]             desc_8_wuser_9_reg;     
wire [31:0]             desc_8_xuser_0_reg;     
wire [31:0]             desc_8_xuser_10_reg;    
wire [31:0]             desc_8_xuser_11_reg;    
wire [31:0]             desc_8_xuser_12_reg;    
wire [31:0]             desc_8_xuser_13_reg;    
wire [31:0]             desc_8_xuser_14_reg;    
wire [31:0]             desc_8_xuser_15_reg;    
wire [31:0]             desc_8_xuser_1_reg;     
wire [31:0]             desc_8_xuser_2_reg;     
wire [31:0]             desc_8_xuser_3_reg;     
wire [31:0]             desc_8_xuser_4_reg;     
wire [31:0]             desc_8_xuser_5_reg;     
wire [31:0]             desc_8_xuser_6_reg;     
wire [31:0]             desc_8_xuser_7_reg;     
wire [31:0]             desc_8_xuser_8_reg;     
wire [31:0]             desc_8_xuser_9_reg;     
wire [31:0]             desc_9_attr_reg;        
wire [31:0]             desc_9_axaddr_0_reg;    
wire [31:0]             desc_9_axaddr_1_reg;    
wire [31:0]             desc_9_axaddr_2_reg;    
wire [31:0]             desc_9_axaddr_3_reg;    
wire [31:0]             desc_9_axid_0_reg;      
wire [31:0]             desc_9_axid_1_reg;      
wire [31:0]             desc_9_axid_2_reg;      
wire [31:0]             desc_9_axid_3_reg;      
wire [31:0]             desc_9_axsize_reg;      
wire [31:0]             desc_9_axuser_0_reg;    
wire [31:0]             desc_9_axuser_10_reg;   
wire [31:0]             desc_9_axuser_11_reg;   
wire [31:0]             desc_9_axuser_12_reg;   
wire [31:0]             desc_9_axuser_13_reg;   
wire [31:0]             desc_9_axuser_14_reg;   
wire [31:0]             desc_9_axuser_15_reg;   
wire [31:0]             desc_9_axuser_1_reg;    
wire [31:0]             desc_9_axuser_2_reg;    
wire [31:0]             desc_9_axuser_3_reg;    
wire [31:0]             desc_9_axuser_4_reg;    
wire [31:0]             desc_9_axuser_5_reg;    
wire [31:0]             desc_9_axuser_6_reg;    
wire [31:0]             desc_9_axuser_7_reg;    
wire [31:0]             desc_9_axuser_8_reg;    
wire [31:0]             desc_9_axuser_9_reg;    
wire [31:0]             desc_9_data_host_addr_0_reg;
wire [31:0]             desc_9_data_host_addr_1_reg;
wire [31:0]             desc_9_data_host_addr_2_reg;
wire [31:0]             desc_9_data_host_addr_3_reg;
wire [31:0]             desc_9_data_offset_reg; 
wire [31:0]             desc_9_size_reg;        
wire [31:0]             desc_9_txn_type_reg;    
wire [31:0]             desc_9_wstrb_host_addr_0_reg;
wire [31:0]             desc_9_wstrb_host_addr_1_reg;
wire [31:0]             desc_9_wstrb_host_addr_2_reg;
wire [31:0]             desc_9_wstrb_host_addr_3_reg;
wire [31:0]             desc_9_wuser_0_reg;     
wire [31:0]             desc_9_wuser_10_reg;    
wire [31:0]             desc_9_wuser_11_reg;    
wire [31:0]             desc_9_wuser_12_reg;    
wire [31:0]             desc_9_wuser_13_reg;    
wire [31:0]             desc_9_wuser_14_reg;    
wire [31:0]             desc_9_wuser_15_reg;    
wire [31:0]             desc_9_wuser_1_reg;     
wire [31:0]             desc_9_wuser_2_reg;     
wire [31:0]             desc_9_wuser_3_reg;     
wire [31:0]             desc_9_wuser_4_reg;     
wire [31:0]             desc_9_wuser_5_reg;     
wire [31:0]             desc_9_wuser_6_reg;     
wire [31:0]             desc_9_wuser_7_reg;     
wire [31:0]             desc_9_wuser_8_reg;     
wire [31:0]             desc_9_wuser_9_reg;     
wire [31:0]             desc_9_xuser_0_reg;     
wire [31:0]             desc_9_xuser_10_reg;    
wire [31:0]             desc_9_xuser_11_reg;    
wire [31:0]             desc_9_xuser_12_reg;    
wire [31:0]             desc_9_xuser_13_reg;    
wire [31:0]             desc_9_xuser_14_reg;    
wire [31:0]             desc_9_xuser_15_reg;    
wire [31:0]             desc_9_xuser_1_reg;     
wire [31:0]             desc_9_xuser_2_reg;     
wire [31:0]             desc_9_xuser_3_reg;     
wire [31:0]             desc_9_xuser_4_reg;     
wire [31:0]             desc_9_xuser_5_reg;     
wire [31:0]             desc_9_xuser_6_reg;     
wire [31:0]             desc_9_xuser_7_reg;     
wire [31:0]             desc_9_xuser_8_reg;     
wire [31:0]             desc_9_xuser_9_reg;     
wire [31:0] 			ih2rb_c2h_intr_status_0_reg   ; 
wire [31:0] 			ih2rb_c2h_intr_status_1_reg   ;
wire [31:0] 			ih2rb_intr_c2h_toggle_status_0_reg   ; 
wire [31:0] 			ih2rb_intr_c2h_toggle_status_1_reg   ; 
wire [31:0] 			ih2rb_c2h_gpio_0_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_1_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_2_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_3_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_4_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_5_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_6_reg   ;
wire [31:0] 			ih2rb_c2h_gpio_7_reg   ; 
wire [31:0] 			ih2rb_c2h_intr_status_0_reg_we; 
wire [31:0] 			ih2rb_c2h_intr_status_1_reg_we;
wire [31:0] 			ih2rb_intr_c2h_toggle_status_0_reg_we; 
wire [31:0] 			ih2rb_intr_c2h_toggle_status_1_reg_we; 
wire [31:0] 			ih2rb_c2h_gpio_0_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_1_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_2_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_3_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_4_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_5_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_6_reg_we;
wire [31:0] 			ih2rb_c2h_gpio_7_reg_we;
   
wire [31:0]             hm2rb_intr_error_status_reg_we;
wire [31:0]             hm2rb_intr_error_status_reg;
wire [(`CLOG2(RAM_SIZE/(S_AXI_USR_DATA_WIDTH/8)))-1:0] hm2rb_rd_addr;
wire [(`CLOG2(RAM_SIZE/(S_AXI_USR_DATA_WIDTH/8)))-1:0] hm2rb_wr_addr;
wire [(S_AXI_USR_DATA_WIDTH/8-1):0] hm2rb_wr_bwe;
wire [S_AXI_USR_DATA_WIDTH-1:0] hm2rb_wr_data;  
wire                    hm2rb_wr_we;            
wire [MAX_DESC-1:0]     hm2uc_done;             
wire [31:0] 			c2h_intr_status_0_reg;  
wire [31:0] 			c2h_intr_status_1_reg;
wire [31:0] 			intr_c2h_toggle_clear_0_reg;  
wire [31:0] 			intr_c2h_toggle_clear_1_reg;
wire [31:0] 			intr_c2h_toggle_status_0_reg;  
wire [31:0] 			intr_c2h_toggle_status_1_reg;
wire [31:0] 			intr_c2h_toggle_enable_0_reg;  
wire [31:0] 			intr_c2h_toggle_enable_1_reg;  
wire [31:0]             intr_error_clear_reg;   
wire [31:0]             intr_error_enable_reg;  
wire [31:0]             intr_error_status_reg;  
wire [31:0] 			h2c_intr_0_reg;         
wire [31:0] 			h2c_intr_1_reg;
wire [31:0] 			h2c_intr_2_reg;         
wire [31:0] 			h2c_intr_3_reg;         
wire [31:0]             intr_h2c_0_reg;         
wire [31:0]             intr_h2c_1_reg;         
wire [31:0]             intr_status_reg;        
wire [31:0]             intr_txn_avail_clear_reg;
wire [31:0]             intr_txn_avail_enable_reg;
wire [31:0]             intr_txn_avail_status_reg;
wire [31:0]             intr_comp_clear_reg;
wire [31:0]             intr_comp_enable_reg;
wire [31:0]             intr_comp_status_reg;
wire [31:0]             resp_fifo_free_level_reg;
wire [31:0]             resp_order_reg;
wire [31:0]             mode_select_reg;        
wire [31:0]             ownership_flip_reg;     
wire [31:0]             ownership_reg;          
wire [S_AXI_USR_DATA_WIDTH-1:0] rb2hm_rd_data;  
wire [(S_AXI_USR_DATA_WIDTH/8-1):0] rb2hm_rd_wstrb;
wire [31:0]             status_busy_reg;        
wire [31:0]             status_resp_comp_reg;   
wire [31:0]             status_resp_reg;        
wire [31:0]             trans_addr_0_reg;       
wire [31:0]             trans_addr_1_reg;       
wire [31:0]             trans_addr_2_reg;       
wire [31:0]             trans_addr_3_reg;       
wire [31:0]             trans_mask_0_reg;       
wire [31:0]             trans_mask_1_reg;       
wire [31:0]             trans_mask_2_reg;       
wire [31:0]             trans_mask_3_reg;       
wire [MAX_DESC-1:0]     uc2hm_trig;             
wire [31:0]             uc2rb_desc_0_attr_reg;  
wire [31:0]             uc2rb_desc_0_attr_reg_we;
wire [31:0]             uc2rb_desc_0_axaddr_0_reg;
wire [31:0]             uc2rb_desc_0_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_0_axaddr_1_reg;
wire [31:0]             uc2rb_desc_0_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_0_axaddr_2_reg;
wire [31:0]             uc2rb_desc_0_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_0_axaddr_3_reg;
wire [31:0]             uc2rb_desc_0_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_0_axid_0_reg;
wire [31:0]             uc2rb_desc_0_axid_0_reg_we;
wire [31:0]             uc2rb_desc_0_axid_1_reg;
wire [31:0]             uc2rb_desc_0_axid_1_reg_we;
wire [31:0]             uc2rb_desc_0_axid_2_reg;
wire [31:0]             uc2rb_desc_0_axid_2_reg_we;
wire [31:0]             uc2rb_desc_0_axid_3_reg;
wire [31:0]             uc2rb_desc_0_axid_3_reg_we;
wire [31:0]             uc2rb_desc_0_axsize_reg;
wire [31:0]             uc2rb_desc_0_axsize_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_0_reg;
wire [31:0]             uc2rb_desc_0_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_10_reg;
wire [31:0]             uc2rb_desc_0_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_11_reg;
wire [31:0]             uc2rb_desc_0_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_12_reg;
wire [31:0]             uc2rb_desc_0_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_13_reg;
wire [31:0]             uc2rb_desc_0_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_14_reg;
wire [31:0]             uc2rb_desc_0_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_15_reg;
wire [31:0]             uc2rb_desc_0_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_1_reg;
wire [31:0]             uc2rb_desc_0_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_2_reg;
wire [31:0]             uc2rb_desc_0_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_3_reg;
wire [31:0]             uc2rb_desc_0_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_4_reg;
wire [31:0]             uc2rb_desc_0_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_5_reg;
wire [31:0]             uc2rb_desc_0_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_6_reg;
wire [31:0]             uc2rb_desc_0_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_7_reg;
wire [31:0]             uc2rb_desc_0_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_8_reg;
wire [31:0]             uc2rb_desc_0_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_0_axuser_9_reg;
wire [31:0]             uc2rb_desc_0_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_0_data_offset_reg;
wire [31:0]             uc2rb_desc_0_data_offset_reg_we;
wire [31:0]             uc2rb_desc_0_size_reg;  
wire [31:0]             uc2rb_desc_0_size_reg_we;
wire [31:0]             uc2rb_desc_0_txn_type_reg;
wire [31:0]             uc2rb_desc_0_txn_type_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_0_reg;
wire [31:0]             uc2rb_desc_0_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_10_reg;
wire [31:0]             uc2rb_desc_0_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_11_reg;
wire [31:0]             uc2rb_desc_0_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_12_reg;
wire [31:0]             uc2rb_desc_0_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_13_reg;
wire [31:0]             uc2rb_desc_0_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_14_reg;
wire [31:0]             uc2rb_desc_0_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_15_reg;
wire [31:0]             uc2rb_desc_0_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_1_reg;
wire [31:0]             uc2rb_desc_0_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_2_reg;
wire [31:0]             uc2rb_desc_0_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_3_reg;
wire [31:0]             uc2rb_desc_0_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_4_reg;
wire [31:0]             uc2rb_desc_0_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_5_reg;
wire [31:0]             uc2rb_desc_0_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_6_reg;
wire [31:0]             uc2rb_desc_0_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_7_reg;
wire [31:0]             uc2rb_desc_0_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_8_reg;
wire [31:0]             uc2rb_desc_0_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_0_wuser_9_reg;
wire [31:0]             uc2rb_desc_0_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_10_attr_reg; 
wire [31:0]             uc2rb_desc_10_attr_reg_we;
wire [31:0]             uc2rb_desc_10_axaddr_0_reg;
wire [31:0]             uc2rb_desc_10_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_10_axaddr_1_reg;
wire [31:0]             uc2rb_desc_10_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_10_axaddr_2_reg;
wire [31:0]             uc2rb_desc_10_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_10_axaddr_3_reg;
wire [31:0]             uc2rb_desc_10_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_10_axid_0_reg;
wire [31:0]             uc2rb_desc_10_axid_0_reg_we;
wire [31:0]             uc2rb_desc_10_axid_1_reg;
wire [31:0]             uc2rb_desc_10_axid_1_reg_we;
wire [31:0]             uc2rb_desc_10_axid_2_reg;
wire [31:0]             uc2rb_desc_10_axid_2_reg_we;
wire [31:0]             uc2rb_desc_10_axid_3_reg;
wire [31:0]             uc2rb_desc_10_axid_3_reg_we;
wire [31:0]             uc2rb_desc_10_axsize_reg;
wire [31:0]             uc2rb_desc_10_axsize_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_0_reg;
wire [31:0]             uc2rb_desc_10_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_10_reg;
wire [31:0]             uc2rb_desc_10_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_11_reg;
wire [31:0]             uc2rb_desc_10_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_12_reg;
wire [31:0]             uc2rb_desc_10_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_13_reg;
wire [31:0]             uc2rb_desc_10_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_14_reg;
wire [31:0]             uc2rb_desc_10_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_15_reg;
wire [31:0]             uc2rb_desc_10_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_1_reg;
wire [31:0]             uc2rb_desc_10_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_2_reg;
wire [31:0]             uc2rb_desc_10_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_3_reg;
wire [31:0]             uc2rb_desc_10_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_4_reg;
wire [31:0]             uc2rb_desc_10_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_5_reg;
wire [31:0]             uc2rb_desc_10_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_6_reg;
wire [31:0]             uc2rb_desc_10_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_7_reg;
wire [31:0]             uc2rb_desc_10_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_8_reg;
wire [31:0]             uc2rb_desc_10_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_10_axuser_9_reg;
wire [31:0]             uc2rb_desc_10_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_10_data_offset_reg;
wire [31:0]             uc2rb_desc_10_data_offset_reg_we;
wire [31:0]             uc2rb_desc_10_size_reg; 
wire [31:0]             uc2rb_desc_10_size_reg_we;
wire [31:0]             uc2rb_desc_10_txn_type_reg;
wire [31:0]             uc2rb_desc_10_txn_type_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_0_reg;
wire [31:0]             uc2rb_desc_10_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_10_reg;
wire [31:0]             uc2rb_desc_10_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_11_reg;
wire [31:0]             uc2rb_desc_10_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_12_reg;
wire [31:0]             uc2rb_desc_10_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_13_reg;
wire [31:0]             uc2rb_desc_10_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_14_reg;
wire [31:0]             uc2rb_desc_10_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_15_reg;
wire [31:0]             uc2rb_desc_10_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_1_reg;
wire [31:0]             uc2rb_desc_10_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_2_reg;
wire [31:0]             uc2rb_desc_10_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_3_reg;
wire [31:0]             uc2rb_desc_10_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_4_reg;
wire [31:0]             uc2rb_desc_10_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_5_reg;
wire [31:0]             uc2rb_desc_10_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_6_reg;
wire [31:0]             uc2rb_desc_10_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_7_reg;
wire [31:0]             uc2rb_desc_10_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_8_reg;
wire [31:0]             uc2rb_desc_10_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_10_wuser_9_reg;
wire [31:0]             uc2rb_desc_10_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_11_attr_reg; 
wire [31:0]             uc2rb_desc_11_attr_reg_we;
wire [31:0]             uc2rb_desc_11_axaddr_0_reg;
wire [31:0]             uc2rb_desc_11_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_11_axaddr_1_reg;
wire [31:0]             uc2rb_desc_11_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_11_axaddr_2_reg;
wire [31:0]             uc2rb_desc_11_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_11_axaddr_3_reg;
wire [31:0]             uc2rb_desc_11_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_11_axid_0_reg;
wire [31:0]             uc2rb_desc_11_axid_0_reg_we;
wire [31:0]             uc2rb_desc_11_axid_1_reg;
wire [31:0]             uc2rb_desc_11_axid_1_reg_we;
wire [31:0]             uc2rb_desc_11_axid_2_reg;
wire [31:0]             uc2rb_desc_11_axid_2_reg_we;
wire [31:0]             uc2rb_desc_11_axid_3_reg;
wire [31:0]             uc2rb_desc_11_axid_3_reg_we;
wire [31:0]             uc2rb_desc_11_axsize_reg;
wire [31:0]             uc2rb_desc_11_axsize_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_0_reg;
wire [31:0]             uc2rb_desc_11_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_10_reg;
wire [31:0]             uc2rb_desc_11_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_11_reg;
wire [31:0]             uc2rb_desc_11_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_12_reg;
wire [31:0]             uc2rb_desc_11_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_13_reg;
wire [31:0]             uc2rb_desc_11_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_14_reg;
wire [31:0]             uc2rb_desc_11_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_15_reg;
wire [31:0]             uc2rb_desc_11_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_1_reg;
wire [31:0]             uc2rb_desc_11_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_2_reg;
wire [31:0]             uc2rb_desc_11_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_3_reg;
wire [31:0]             uc2rb_desc_11_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_4_reg;
wire [31:0]             uc2rb_desc_11_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_5_reg;
wire [31:0]             uc2rb_desc_11_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_6_reg;
wire [31:0]             uc2rb_desc_11_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_7_reg;
wire [31:0]             uc2rb_desc_11_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_8_reg;
wire [31:0]             uc2rb_desc_11_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_11_axuser_9_reg;
wire [31:0]             uc2rb_desc_11_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_11_data_offset_reg;
wire [31:0]             uc2rb_desc_11_data_offset_reg_we;
wire [31:0]             uc2rb_desc_11_size_reg; 
wire [31:0]             uc2rb_desc_11_size_reg_we;
wire [31:0]             uc2rb_desc_11_txn_type_reg;
wire [31:0]             uc2rb_desc_11_txn_type_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_0_reg;
wire [31:0]             uc2rb_desc_11_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_10_reg;
wire [31:0]             uc2rb_desc_11_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_11_reg;
wire [31:0]             uc2rb_desc_11_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_12_reg;
wire [31:0]             uc2rb_desc_11_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_13_reg;
wire [31:0]             uc2rb_desc_11_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_14_reg;
wire [31:0]             uc2rb_desc_11_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_15_reg;
wire [31:0]             uc2rb_desc_11_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_1_reg;
wire [31:0]             uc2rb_desc_11_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_2_reg;
wire [31:0]             uc2rb_desc_11_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_3_reg;
wire [31:0]             uc2rb_desc_11_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_4_reg;
wire [31:0]             uc2rb_desc_11_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_5_reg;
wire [31:0]             uc2rb_desc_11_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_6_reg;
wire [31:0]             uc2rb_desc_11_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_7_reg;
wire [31:0]             uc2rb_desc_11_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_8_reg;
wire [31:0]             uc2rb_desc_11_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_11_wuser_9_reg;
wire [31:0]             uc2rb_desc_11_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_12_attr_reg; 
wire [31:0]             uc2rb_desc_12_attr_reg_we;
wire [31:0]             uc2rb_desc_12_axaddr_0_reg;
wire [31:0]             uc2rb_desc_12_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_12_axaddr_1_reg;
wire [31:0]             uc2rb_desc_12_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_12_axaddr_2_reg;
wire [31:0]             uc2rb_desc_12_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_12_axaddr_3_reg;
wire [31:0]             uc2rb_desc_12_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_12_axid_0_reg;
wire [31:0]             uc2rb_desc_12_axid_0_reg_we;
wire [31:0]             uc2rb_desc_12_axid_1_reg;
wire [31:0]             uc2rb_desc_12_axid_1_reg_we;
wire [31:0]             uc2rb_desc_12_axid_2_reg;
wire [31:0]             uc2rb_desc_12_axid_2_reg_we;
wire [31:0]             uc2rb_desc_12_axid_3_reg;
wire [31:0]             uc2rb_desc_12_axid_3_reg_we;
wire [31:0]             uc2rb_desc_12_axsize_reg;
wire [31:0]             uc2rb_desc_12_axsize_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_0_reg;
wire [31:0]             uc2rb_desc_12_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_10_reg;
wire [31:0]             uc2rb_desc_12_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_11_reg;
wire [31:0]             uc2rb_desc_12_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_12_reg;
wire [31:0]             uc2rb_desc_12_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_13_reg;
wire [31:0]             uc2rb_desc_12_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_14_reg;
wire [31:0]             uc2rb_desc_12_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_15_reg;
wire [31:0]             uc2rb_desc_12_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_1_reg;
wire [31:0]             uc2rb_desc_12_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_2_reg;
wire [31:0]             uc2rb_desc_12_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_3_reg;
wire [31:0]             uc2rb_desc_12_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_4_reg;
wire [31:0]             uc2rb_desc_12_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_5_reg;
wire [31:0]             uc2rb_desc_12_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_6_reg;
wire [31:0]             uc2rb_desc_12_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_7_reg;
wire [31:0]             uc2rb_desc_12_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_8_reg;
wire [31:0]             uc2rb_desc_12_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_12_axuser_9_reg;
wire [31:0]             uc2rb_desc_12_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_12_data_offset_reg;
wire [31:0]             uc2rb_desc_12_data_offset_reg_we;
wire [31:0]             uc2rb_desc_12_size_reg; 
wire [31:0]             uc2rb_desc_12_size_reg_we;
wire [31:0]             uc2rb_desc_12_txn_type_reg;
wire [31:0]             uc2rb_desc_12_txn_type_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_0_reg;
wire [31:0]             uc2rb_desc_12_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_10_reg;
wire [31:0]             uc2rb_desc_12_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_11_reg;
wire [31:0]             uc2rb_desc_12_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_12_reg;
wire [31:0]             uc2rb_desc_12_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_13_reg;
wire [31:0]             uc2rb_desc_12_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_14_reg;
wire [31:0]             uc2rb_desc_12_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_15_reg;
wire [31:0]             uc2rb_desc_12_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_1_reg;
wire [31:0]             uc2rb_desc_12_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_2_reg;
wire [31:0]             uc2rb_desc_12_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_3_reg;
wire [31:0]             uc2rb_desc_12_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_4_reg;
wire [31:0]             uc2rb_desc_12_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_5_reg;
wire [31:0]             uc2rb_desc_12_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_6_reg;
wire [31:0]             uc2rb_desc_12_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_7_reg;
wire [31:0]             uc2rb_desc_12_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_8_reg;
wire [31:0]             uc2rb_desc_12_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_12_wuser_9_reg;
wire [31:0]             uc2rb_desc_12_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_13_attr_reg; 
wire [31:0]             uc2rb_desc_13_attr_reg_we;
wire [31:0]             uc2rb_desc_13_axaddr_0_reg;
wire [31:0]             uc2rb_desc_13_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_13_axaddr_1_reg;
wire [31:0]             uc2rb_desc_13_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_13_axaddr_2_reg;
wire [31:0]             uc2rb_desc_13_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_13_axaddr_3_reg;
wire [31:0]             uc2rb_desc_13_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_13_axid_0_reg;
wire [31:0]             uc2rb_desc_13_axid_0_reg_we;
wire [31:0]             uc2rb_desc_13_axid_1_reg;
wire [31:0]             uc2rb_desc_13_axid_1_reg_we;
wire [31:0]             uc2rb_desc_13_axid_2_reg;
wire [31:0]             uc2rb_desc_13_axid_2_reg_we;
wire [31:0]             uc2rb_desc_13_axid_3_reg;
wire [31:0]             uc2rb_desc_13_axid_3_reg_we;
wire [31:0]             uc2rb_desc_13_axsize_reg;
wire [31:0]             uc2rb_desc_13_axsize_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_0_reg;
wire [31:0]             uc2rb_desc_13_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_10_reg;
wire [31:0]             uc2rb_desc_13_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_11_reg;
wire [31:0]             uc2rb_desc_13_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_12_reg;
wire [31:0]             uc2rb_desc_13_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_13_reg;
wire [31:0]             uc2rb_desc_13_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_14_reg;
wire [31:0]             uc2rb_desc_13_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_15_reg;
wire [31:0]             uc2rb_desc_13_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_1_reg;
wire [31:0]             uc2rb_desc_13_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_2_reg;
wire [31:0]             uc2rb_desc_13_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_3_reg;
wire [31:0]             uc2rb_desc_13_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_4_reg;
wire [31:0]             uc2rb_desc_13_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_5_reg;
wire [31:0]             uc2rb_desc_13_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_6_reg;
wire [31:0]             uc2rb_desc_13_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_7_reg;
wire [31:0]             uc2rb_desc_13_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_8_reg;
wire [31:0]             uc2rb_desc_13_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_13_axuser_9_reg;
wire [31:0]             uc2rb_desc_13_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_13_data_offset_reg;
wire [31:0]             uc2rb_desc_13_data_offset_reg_we;
wire [31:0]             uc2rb_desc_13_size_reg; 
wire [31:0]             uc2rb_desc_13_size_reg_we;
wire [31:0]             uc2rb_desc_13_txn_type_reg;
wire [31:0]             uc2rb_desc_13_txn_type_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_0_reg;
wire [31:0]             uc2rb_desc_13_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_10_reg;
wire [31:0]             uc2rb_desc_13_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_11_reg;
wire [31:0]             uc2rb_desc_13_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_12_reg;
wire [31:0]             uc2rb_desc_13_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_13_reg;
wire [31:0]             uc2rb_desc_13_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_14_reg;
wire [31:0]             uc2rb_desc_13_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_15_reg;
wire [31:0]             uc2rb_desc_13_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_1_reg;
wire [31:0]             uc2rb_desc_13_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_2_reg;
wire [31:0]             uc2rb_desc_13_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_3_reg;
wire [31:0]             uc2rb_desc_13_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_4_reg;
wire [31:0]             uc2rb_desc_13_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_5_reg;
wire [31:0]             uc2rb_desc_13_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_6_reg;
wire [31:0]             uc2rb_desc_13_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_7_reg;
wire [31:0]             uc2rb_desc_13_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_8_reg;
wire [31:0]             uc2rb_desc_13_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_13_wuser_9_reg;
wire [31:0]             uc2rb_desc_13_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_14_attr_reg; 
wire [31:0]             uc2rb_desc_14_attr_reg_we;
wire [31:0]             uc2rb_desc_14_axaddr_0_reg;
wire [31:0]             uc2rb_desc_14_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_14_axaddr_1_reg;
wire [31:0]             uc2rb_desc_14_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_14_axaddr_2_reg;
wire [31:0]             uc2rb_desc_14_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_14_axaddr_3_reg;
wire [31:0]             uc2rb_desc_14_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_14_axid_0_reg;
wire [31:0]             uc2rb_desc_14_axid_0_reg_we;
wire [31:0]             uc2rb_desc_14_axid_1_reg;
wire [31:0]             uc2rb_desc_14_axid_1_reg_we;
wire [31:0]             uc2rb_desc_14_axid_2_reg;
wire [31:0]             uc2rb_desc_14_axid_2_reg_we;
wire [31:0]             uc2rb_desc_14_axid_3_reg;
wire [31:0]             uc2rb_desc_14_axid_3_reg_we;
wire [31:0]             uc2rb_desc_14_axsize_reg;
wire [31:0]             uc2rb_desc_14_axsize_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_0_reg;
wire [31:0]             uc2rb_desc_14_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_10_reg;
wire [31:0]             uc2rb_desc_14_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_11_reg;
wire [31:0]             uc2rb_desc_14_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_12_reg;
wire [31:0]             uc2rb_desc_14_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_13_reg;
wire [31:0]             uc2rb_desc_14_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_14_reg;
wire [31:0]             uc2rb_desc_14_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_15_reg;
wire [31:0]             uc2rb_desc_14_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_1_reg;
wire [31:0]             uc2rb_desc_14_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_2_reg;
wire [31:0]             uc2rb_desc_14_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_3_reg;
wire [31:0]             uc2rb_desc_14_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_4_reg;
wire [31:0]             uc2rb_desc_14_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_5_reg;
wire [31:0]             uc2rb_desc_14_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_6_reg;
wire [31:0]             uc2rb_desc_14_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_7_reg;
wire [31:0]             uc2rb_desc_14_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_8_reg;
wire [31:0]             uc2rb_desc_14_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_14_axuser_9_reg;
wire [31:0]             uc2rb_desc_14_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_14_data_offset_reg;
wire [31:0]             uc2rb_desc_14_data_offset_reg_we;
wire [31:0]             uc2rb_desc_14_size_reg; 
wire [31:0]             uc2rb_desc_14_size_reg_we;
wire [31:0]             uc2rb_desc_14_txn_type_reg;
wire [31:0]             uc2rb_desc_14_txn_type_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_0_reg;
wire [31:0]             uc2rb_desc_14_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_10_reg;
wire [31:0]             uc2rb_desc_14_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_11_reg;
wire [31:0]             uc2rb_desc_14_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_12_reg;
wire [31:0]             uc2rb_desc_14_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_13_reg;
wire [31:0]             uc2rb_desc_14_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_14_reg;
wire [31:0]             uc2rb_desc_14_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_15_reg;
wire [31:0]             uc2rb_desc_14_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_1_reg;
wire [31:0]             uc2rb_desc_14_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_2_reg;
wire [31:0]             uc2rb_desc_14_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_3_reg;
wire [31:0]             uc2rb_desc_14_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_4_reg;
wire [31:0]             uc2rb_desc_14_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_5_reg;
wire [31:0]             uc2rb_desc_14_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_6_reg;
wire [31:0]             uc2rb_desc_14_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_7_reg;
wire [31:0]             uc2rb_desc_14_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_8_reg;
wire [31:0]             uc2rb_desc_14_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_14_wuser_9_reg;
wire [31:0]             uc2rb_desc_14_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_15_attr_reg; 
wire [31:0]             uc2rb_desc_15_attr_reg_we;
wire [31:0]             uc2rb_desc_15_axaddr_0_reg;
wire [31:0]             uc2rb_desc_15_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_15_axaddr_1_reg;
wire [31:0]             uc2rb_desc_15_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_15_axaddr_2_reg;
wire [31:0]             uc2rb_desc_15_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_15_axaddr_3_reg;
wire [31:0]             uc2rb_desc_15_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_15_axid_0_reg;
wire [31:0]             uc2rb_desc_15_axid_0_reg_we;
wire [31:0]             uc2rb_desc_15_axid_1_reg;
wire [31:0]             uc2rb_desc_15_axid_1_reg_we;
wire [31:0]             uc2rb_desc_15_axid_2_reg;
wire [31:0]             uc2rb_desc_15_axid_2_reg_we;
wire [31:0]             uc2rb_desc_15_axid_3_reg;
wire [31:0]             uc2rb_desc_15_axid_3_reg_we;
wire [31:0]             uc2rb_desc_15_axsize_reg;
wire [31:0]             uc2rb_desc_15_axsize_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_0_reg;
wire [31:0]             uc2rb_desc_15_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_10_reg;
wire [31:0]             uc2rb_desc_15_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_11_reg;
wire [31:0]             uc2rb_desc_15_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_12_reg;
wire [31:0]             uc2rb_desc_15_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_13_reg;
wire [31:0]             uc2rb_desc_15_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_14_reg;
wire [31:0]             uc2rb_desc_15_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_15_reg;
wire [31:0]             uc2rb_desc_15_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_1_reg;
wire [31:0]             uc2rb_desc_15_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_2_reg;
wire [31:0]             uc2rb_desc_15_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_3_reg;
wire [31:0]             uc2rb_desc_15_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_4_reg;
wire [31:0]             uc2rb_desc_15_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_5_reg;
wire [31:0]             uc2rb_desc_15_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_6_reg;
wire [31:0]             uc2rb_desc_15_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_7_reg;
wire [31:0]             uc2rb_desc_15_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_8_reg;
wire [31:0]             uc2rb_desc_15_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_15_axuser_9_reg;
wire [31:0]             uc2rb_desc_15_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_15_data_offset_reg;
wire [31:0]             uc2rb_desc_15_data_offset_reg_we;
wire [31:0]             uc2rb_desc_15_size_reg; 
wire [31:0]             uc2rb_desc_15_size_reg_we;
wire [31:0]             uc2rb_desc_15_txn_type_reg;
wire [31:0]             uc2rb_desc_15_txn_type_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_0_reg;
wire [31:0]             uc2rb_desc_15_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_10_reg;
wire [31:0]             uc2rb_desc_15_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_11_reg;
wire [31:0]             uc2rb_desc_15_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_12_reg;
wire [31:0]             uc2rb_desc_15_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_13_reg;
wire [31:0]             uc2rb_desc_15_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_14_reg;
wire [31:0]             uc2rb_desc_15_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_15_reg;
wire [31:0]             uc2rb_desc_15_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_1_reg;
wire [31:0]             uc2rb_desc_15_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_2_reg;
wire [31:0]             uc2rb_desc_15_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_3_reg;
wire [31:0]             uc2rb_desc_15_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_4_reg;
wire [31:0]             uc2rb_desc_15_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_5_reg;
wire [31:0]             uc2rb_desc_15_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_6_reg;
wire [31:0]             uc2rb_desc_15_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_7_reg;
wire [31:0]             uc2rb_desc_15_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_8_reg;
wire [31:0]             uc2rb_desc_15_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_15_wuser_9_reg;
wire [31:0]             uc2rb_desc_15_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_1_attr_reg;  
wire [31:0]             uc2rb_desc_1_attr_reg_we;
wire [31:0]             uc2rb_desc_1_axaddr_0_reg;
wire [31:0]             uc2rb_desc_1_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_1_axaddr_1_reg;
wire [31:0]             uc2rb_desc_1_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_1_axaddr_2_reg;
wire [31:0]             uc2rb_desc_1_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_1_axaddr_3_reg;
wire [31:0]             uc2rb_desc_1_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_1_axid_0_reg;
wire [31:0]             uc2rb_desc_1_axid_0_reg_we;
wire [31:0]             uc2rb_desc_1_axid_1_reg;
wire [31:0]             uc2rb_desc_1_axid_1_reg_we;
wire [31:0]             uc2rb_desc_1_axid_2_reg;
wire [31:0]             uc2rb_desc_1_axid_2_reg_we;
wire [31:0]             uc2rb_desc_1_axid_3_reg;
wire [31:0]             uc2rb_desc_1_axid_3_reg_we;
wire [31:0]             uc2rb_desc_1_axsize_reg;
wire [31:0]             uc2rb_desc_1_axsize_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_0_reg;
wire [31:0]             uc2rb_desc_1_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_10_reg;
wire [31:0]             uc2rb_desc_1_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_11_reg;
wire [31:0]             uc2rb_desc_1_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_12_reg;
wire [31:0]             uc2rb_desc_1_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_13_reg;
wire [31:0]             uc2rb_desc_1_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_14_reg;
wire [31:0]             uc2rb_desc_1_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_15_reg;
wire [31:0]             uc2rb_desc_1_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_1_reg;
wire [31:0]             uc2rb_desc_1_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_2_reg;
wire [31:0]             uc2rb_desc_1_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_3_reg;
wire [31:0]             uc2rb_desc_1_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_4_reg;
wire [31:0]             uc2rb_desc_1_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_5_reg;
wire [31:0]             uc2rb_desc_1_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_6_reg;
wire [31:0]             uc2rb_desc_1_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_7_reg;
wire [31:0]             uc2rb_desc_1_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_8_reg;
wire [31:0]             uc2rb_desc_1_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_1_axuser_9_reg;
wire [31:0]             uc2rb_desc_1_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_1_data_offset_reg;
wire [31:0]             uc2rb_desc_1_data_offset_reg_we;
wire [31:0]             uc2rb_desc_1_size_reg;  
wire [31:0]             uc2rb_desc_1_size_reg_we;
wire [31:0]             uc2rb_desc_1_txn_type_reg;
wire [31:0]             uc2rb_desc_1_txn_type_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_0_reg;
wire [31:0]             uc2rb_desc_1_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_10_reg;
wire [31:0]             uc2rb_desc_1_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_11_reg;
wire [31:0]             uc2rb_desc_1_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_12_reg;
wire [31:0]             uc2rb_desc_1_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_13_reg;
wire [31:0]             uc2rb_desc_1_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_14_reg;
wire [31:0]             uc2rb_desc_1_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_15_reg;
wire [31:0]             uc2rb_desc_1_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_1_reg;
wire [31:0]             uc2rb_desc_1_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_2_reg;
wire [31:0]             uc2rb_desc_1_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_3_reg;
wire [31:0]             uc2rb_desc_1_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_4_reg;
wire [31:0]             uc2rb_desc_1_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_5_reg;
wire [31:0]             uc2rb_desc_1_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_6_reg;
wire [31:0]             uc2rb_desc_1_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_7_reg;
wire [31:0]             uc2rb_desc_1_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_8_reg;
wire [31:0]             uc2rb_desc_1_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_1_wuser_9_reg;
wire [31:0]             uc2rb_desc_1_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_2_attr_reg;  
wire [31:0]             uc2rb_desc_2_attr_reg_we;
wire [31:0]             uc2rb_desc_2_axaddr_0_reg;
wire [31:0]             uc2rb_desc_2_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_2_axaddr_1_reg;
wire [31:0]             uc2rb_desc_2_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_2_axaddr_2_reg;
wire [31:0]             uc2rb_desc_2_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_2_axaddr_3_reg;
wire [31:0]             uc2rb_desc_2_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_2_axid_0_reg;
wire [31:0]             uc2rb_desc_2_axid_0_reg_we;
wire [31:0]             uc2rb_desc_2_axid_1_reg;
wire [31:0]             uc2rb_desc_2_axid_1_reg_we;
wire [31:0]             uc2rb_desc_2_axid_2_reg;
wire [31:0]             uc2rb_desc_2_axid_2_reg_we;
wire [31:0]             uc2rb_desc_2_axid_3_reg;
wire [31:0]             uc2rb_desc_2_axid_3_reg_we;
wire [31:0]             uc2rb_desc_2_axsize_reg;
wire [31:0]             uc2rb_desc_2_axsize_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_0_reg;
wire [31:0]             uc2rb_desc_2_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_10_reg;
wire [31:0]             uc2rb_desc_2_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_11_reg;
wire [31:0]             uc2rb_desc_2_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_12_reg;
wire [31:0]             uc2rb_desc_2_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_13_reg;
wire [31:0]             uc2rb_desc_2_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_14_reg;
wire [31:0]             uc2rb_desc_2_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_15_reg;
wire [31:0]             uc2rb_desc_2_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_1_reg;
wire [31:0]             uc2rb_desc_2_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_2_reg;
wire [31:0]             uc2rb_desc_2_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_3_reg;
wire [31:0]             uc2rb_desc_2_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_4_reg;
wire [31:0]             uc2rb_desc_2_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_5_reg;
wire [31:0]             uc2rb_desc_2_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_6_reg;
wire [31:0]             uc2rb_desc_2_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_7_reg;
wire [31:0]             uc2rb_desc_2_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_8_reg;
wire [31:0]             uc2rb_desc_2_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_2_axuser_9_reg;
wire [31:0]             uc2rb_desc_2_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_2_data_offset_reg;
wire [31:0]             uc2rb_desc_2_data_offset_reg_we;
wire [31:0]             uc2rb_desc_2_size_reg;  
wire [31:0]             uc2rb_desc_2_size_reg_we;
wire [31:0]             uc2rb_desc_2_txn_type_reg;
wire [31:0]             uc2rb_desc_2_txn_type_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_0_reg;
wire [31:0]             uc2rb_desc_2_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_10_reg;
wire [31:0]             uc2rb_desc_2_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_11_reg;
wire [31:0]             uc2rb_desc_2_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_12_reg;
wire [31:0]             uc2rb_desc_2_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_13_reg;
wire [31:0]             uc2rb_desc_2_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_14_reg;
wire [31:0]             uc2rb_desc_2_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_15_reg;
wire [31:0]             uc2rb_desc_2_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_1_reg;
wire [31:0]             uc2rb_desc_2_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_2_reg;
wire [31:0]             uc2rb_desc_2_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_3_reg;
wire [31:0]             uc2rb_desc_2_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_4_reg;
wire [31:0]             uc2rb_desc_2_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_5_reg;
wire [31:0]             uc2rb_desc_2_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_6_reg;
wire [31:0]             uc2rb_desc_2_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_7_reg;
wire [31:0]             uc2rb_desc_2_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_8_reg;
wire [31:0]             uc2rb_desc_2_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_2_wuser_9_reg;
wire [31:0]             uc2rb_desc_2_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_3_attr_reg;  
wire [31:0]             uc2rb_desc_3_attr_reg_we;
wire [31:0]             uc2rb_desc_3_axaddr_0_reg;
wire [31:0]             uc2rb_desc_3_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_3_axaddr_1_reg;
wire [31:0]             uc2rb_desc_3_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_3_axaddr_2_reg;
wire [31:0]             uc2rb_desc_3_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_3_axaddr_3_reg;
wire [31:0]             uc2rb_desc_3_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_3_axid_0_reg;
wire [31:0]             uc2rb_desc_3_axid_0_reg_we;
wire [31:0]             uc2rb_desc_3_axid_1_reg;
wire [31:0]             uc2rb_desc_3_axid_1_reg_we;
wire [31:0]             uc2rb_desc_3_axid_2_reg;
wire [31:0]             uc2rb_desc_3_axid_2_reg_we;
wire [31:0]             uc2rb_desc_3_axid_3_reg;
wire [31:0]             uc2rb_desc_3_axid_3_reg_we;
wire [31:0]             uc2rb_desc_3_axsize_reg;
wire [31:0]             uc2rb_desc_3_axsize_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_0_reg;
wire [31:0]             uc2rb_desc_3_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_10_reg;
wire [31:0]             uc2rb_desc_3_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_11_reg;
wire [31:0]             uc2rb_desc_3_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_12_reg;
wire [31:0]             uc2rb_desc_3_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_13_reg;
wire [31:0]             uc2rb_desc_3_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_14_reg;
wire [31:0]             uc2rb_desc_3_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_15_reg;
wire [31:0]             uc2rb_desc_3_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_1_reg;
wire [31:0]             uc2rb_desc_3_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_2_reg;
wire [31:0]             uc2rb_desc_3_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_3_reg;
wire [31:0]             uc2rb_desc_3_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_4_reg;
wire [31:0]             uc2rb_desc_3_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_5_reg;
wire [31:0]             uc2rb_desc_3_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_6_reg;
wire [31:0]             uc2rb_desc_3_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_7_reg;
wire [31:0]             uc2rb_desc_3_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_8_reg;
wire [31:0]             uc2rb_desc_3_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_3_axuser_9_reg;
wire [31:0]             uc2rb_desc_3_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_3_data_offset_reg;
wire [31:0]             uc2rb_desc_3_data_offset_reg_we;
wire [31:0]             uc2rb_desc_3_size_reg;  
wire [31:0]             uc2rb_desc_3_size_reg_we;
wire [31:0]             uc2rb_desc_3_txn_type_reg;
wire [31:0]             uc2rb_desc_3_txn_type_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_0_reg;
wire [31:0]             uc2rb_desc_3_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_10_reg;
wire [31:0]             uc2rb_desc_3_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_11_reg;
wire [31:0]             uc2rb_desc_3_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_12_reg;
wire [31:0]             uc2rb_desc_3_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_13_reg;
wire [31:0]             uc2rb_desc_3_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_14_reg;
wire [31:0]             uc2rb_desc_3_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_15_reg;
wire [31:0]             uc2rb_desc_3_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_1_reg;
wire [31:0]             uc2rb_desc_3_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_2_reg;
wire [31:0]             uc2rb_desc_3_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_3_reg;
wire [31:0]             uc2rb_desc_3_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_4_reg;
wire [31:0]             uc2rb_desc_3_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_5_reg;
wire [31:0]             uc2rb_desc_3_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_6_reg;
wire [31:0]             uc2rb_desc_3_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_7_reg;
wire [31:0]             uc2rb_desc_3_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_8_reg;
wire [31:0]             uc2rb_desc_3_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_3_wuser_9_reg;
wire [31:0]             uc2rb_desc_3_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_4_attr_reg;  
wire [31:0]             uc2rb_desc_4_attr_reg_we;
wire [31:0]             uc2rb_desc_4_axaddr_0_reg;
wire [31:0]             uc2rb_desc_4_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_4_axaddr_1_reg;
wire [31:0]             uc2rb_desc_4_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_4_axaddr_2_reg;
wire [31:0]             uc2rb_desc_4_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_4_axaddr_3_reg;
wire [31:0]             uc2rb_desc_4_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_4_axid_0_reg;
wire [31:0]             uc2rb_desc_4_axid_0_reg_we;
wire [31:0]             uc2rb_desc_4_axid_1_reg;
wire [31:0]             uc2rb_desc_4_axid_1_reg_we;
wire [31:0]             uc2rb_desc_4_axid_2_reg;
wire [31:0]             uc2rb_desc_4_axid_2_reg_we;
wire [31:0]             uc2rb_desc_4_axid_3_reg;
wire [31:0]             uc2rb_desc_4_axid_3_reg_we;
wire [31:0]             uc2rb_desc_4_axsize_reg;
wire [31:0]             uc2rb_desc_4_axsize_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_0_reg;
wire [31:0]             uc2rb_desc_4_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_10_reg;
wire [31:0]             uc2rb_desc_4_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_11_reg;
wire [31:0]             uc2rb_desc_4_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_12_reg;
wire [31:0]             uc2rb_desc_4_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_13_reg;
wire [31:0]             uc2rb_desc_4_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_14_reg;
wire [31:0]             uc2rb_desc_4_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_15_reg;
wire [31:0]             uc2rb_desc_4_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_1_reg;
wire [31:0]             uc2rb_desc_4_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_2_reg;
wire [31:0]             uc2rb_desc_4_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_3_reg;
wire [31:0]             uc2rb_desc_4_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_4_reg;
wire [31:0]             uc2rb_desc_4_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_5_reg;
wire [31:0]             uc2rb_desc_4_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_6_reg;
wire [31:0]             uc2rb_desc_4_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_7_reg;
wire [31:0]             uc2rb_desc_4_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_8_reg;
wire [31:0]             uc2rb_desc_4_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_4_axuser_9_reg;
wire [31:0]             uc2rb_desc_4_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_4_data_offset_reg;
wire [31:0]             uc2rb_desc_4_data_offset_reg_we;
wire [31:0]             uc2rb_desc_4_size_reg;  
wire [31:0]             uc2rb_desc_4_size_reg_we;
wire [31:0]             uc2rb_desc_4_txn_type_reg;
wire [31:0]             uc2rb_desc_4_txn_type_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_0_reg;
wire [31:0]             uc2rb_desc_4_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_10_reg;
wire [31:0]             uc2rb_desc_4_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_11_reg;
wire [31:0]             uc2rb_desc_4_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_12_reg;
wire [31:0]             uc2rb_desc_4_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_13_reg;
wire [31:0]             uc2rb_desc_4_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_14_reg;
wire [31:0]             uc2rb_desc_4_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_15_reg;
wire [31:0]             uc2rb_desc_4_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_1_reg;
wire [31:0]             uc2rb_desc_4_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_2_reg;
wire [31:0]             uc2rb_desc_4_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_3_reg;
wire [31:0]             uc2rb_desc_4_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_4_reg;
wire [31:0]             uc2rb_desc_4_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_5_reg;
wire [31:0]             uc2rb_desc_4_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_6_reg;
wire [31:0]             uc2rb_desc_4_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_7_reg;
wire [31:0]             uc2rb_desc_4_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_8_reg;
wire [31:0]             uc2rb_desc_4_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_4_wuser_9_reg;
wire [31:0]             uc2rb_desc_4_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_5_attr_reg;  
wire [31:0]             uc2rb_desc_5_attr_reg_we;
wire [31:0]             uc2rb_desc_5_axaddr_0_reg;
wire [31:0]             uc2rb_desc_5_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_5_axaddr_1_reg;
wire [31:0]             uc2rb_desc_5_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_5_axaddr_2_reg;
wire [31:0]             uc2rb_desc_5_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_5_axaddr_3_reg;
wire [31:0]             uc2rb_desc_5_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_5_axid_0_reg;
wire [31:0]             uc2rb_desc_5_axid_0_reg_we;
wire [31:0]             uc2rb_desc_5_axid_1_reg;
wire [31:0]             uc2rb_desc_5_axid_1_reg_we;
wire [31:0]             uc2rb_desc_5_axid_2_reg;
wire [31:0]             uc2rb_desc_5_axid_2_reg_we;
wire [31:0]             uc2rb_desc_5_axid_3_reg;
wire [31:0]             uc2rb_desc_5_axid_3_reg_we;
wire [31:0]             uc2rb_desc_5_axsize_reg;
wire [31:0]             uc2rb_desc_5_axsize_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_0_reg;
wire [31:0]             uc2rb_desc_5_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_10_reg;
wire [31:0]             uc2rb_desc_5_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_11_reg;
wire [31:0]             uc2rb_desc_5_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_12_reg;
wire [31:0]             uc2rb_desc_5_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_13_reg;
wire [31:0]             uc2rb_desc_5_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_14_reg;
wire [31:0]             uc2rb_desc_5_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_15_reg;
wire [31:0]             uc2rb_desc_5_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_1_reg;
wire [31:0]             uc2rb_desc_5_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_2_reg;
wire [31:0]             uc2rb_desc_5_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_3_reg;
wire [31:0]             uc2rb_desc_5_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_4_reg;
wire [31:0]             uc2rb_desc_5_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_5_reg;
wire [31:0]             uc2rb_desc_5_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_6_reg;
wire [31:0]             uc2rb_desc_5_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_7_reg;
wire [31:0]             uc2rb_desc_5_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_8_reg;
wire [31:0]             uc2rb_desc_5_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_5_axuser_9_reg;
wire [31:0]             uc2rb_desc_5_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_5_data_offset_reg;
wire [31:0]             uc2rb_desc_5_data_offset_reg_we;
wire [31:0]             uc2rb_desc_5_size_reg;  
wire [31:0]             uc2rb_desc_5_size_reg_we;
wire [31:0]             uc2rb_desc_5_txn_type_reg;
wire [31:0]             uc2rb_desc_5_txn_type_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_0_reg;
wire [31:0]             uc2rb_desc_5_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_10_reg;
wire [31:0]             uc2rb_desc_5_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_11_reg;
wire [31:0]             uc2rb_desc_5_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_12_reg;
wire [31:0]             uc2rb_desc_5_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_13_reg;
wire [31:0]             uc2rb_desc_5_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_14_reg;
wire [31:0]             uc2rb_desc_5_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_15_reg;
wire [31:0]             uc2rb_desc_5_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_1_reg;
wire [31:0]             uc2rb_desc_5_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_2_reg;
wire [31:0]             uc2rb_desc_5_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_3_reg;
wire [31:0]             uc2rb_desc_5_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_4_reg;
wire [31:0]             uc2rb_desc_5_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_5_reg;
wire [31:0]             uc2rb_desc_5_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_6_reg;
wire [31:0]             uc2rb_desc_5_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_7_reg;
wire [31:0]             uc2rb_desc_5_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_8_reg;
wire [31:0]             uc2rb_desc_5_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_5_wuser_9_reg;
wire [31:0]             uc2rb_desc_5_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_6_attr_reg;  
wire [31:0]             uc2rb_desc_6_attr_reg_we;
wire [31:0]             uc2rb_desc_6_axaddr_0_reg;
wire [31:0]             uc2rb_desc_6_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_6_axaddr_1_reg;
wire [31:0]             uc2rb_desc_6_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_6_axaddr_2_reg;
wire [31:0]             uc2rb_desc_6_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_6_axaddr_3_reg;
wire [31:0]             uc2rb_desc_6_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_6_axid_0_reg;
wire [31:0]             uc2rb_desc_6_axid_0_reg_we;
wire [31:0]             uc2rb_desc_6_axid_1_reg;
wire [31:0]             uc2rb_desc_6_axid_1_reg_we;
wire [31:0]             uc2rb_desc_6_axid_2_reg;
wire [31:0]             uc2rb_desc_6_axid_2_reg_we;
wire [31:0]             uc2rb_desc_6_axid_3_reg;
wire [31:0]             uc2rb_desc_6_axid_3_reg_we;
wire [31:0]             uc2rb_desc_6_axsize_reg;
wire [31:0]             uc2rb_desc_6_axsize_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_0_reg;
wire [31:0]             uc2rb_desc_6_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_10_reg;
wire [31:0]             uc2rb_desc_6_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_11_reg;
wire [31:0]             uc2rb_desc_6_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_12_reg;
wire [31:0]             uc2rb_desc_6_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_13_reg;
wire [31:0]             uc2rb_desc_6_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_14_reg;
wire [31:0]             uc2rb_desc_6_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_15_reg;
wire [31:0]             uc2rb_desc_6_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_1_reg;
wire [31:0]             uc2rb_desc_6_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_2_reg;
wire [31:0]             uc2rb_desc_6_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_3_reg;
wire [31:0]             uc2rb_desc_6_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_4_reg;
wire [31:0]             uc2rb_desc_6_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_5_reg;
wire [31:0]             uc2rb_desc_6_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_6_reg;
wire [31:0]             uc2rb_desc_6_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_7_reg;
wire [31:0]             uc2rb_desc_6_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_8_reg;
wire [31:0]             uc2rb_desc_6_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_6_axuser_9_reg;
wire [31:0]             uc2rb_desc_6_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_6_data_offset_reg;
wire [31:0]             uc2rb_desc_6_data_offset_reg_we;
wire [31:0]             uc2rb_desc_6_size_reg;  
wire [31:0]             uc2rb_desc_6_size_reg_we;
wire [31:0]             uc2rb_desc_6_txn_type_reg;
wire [31:0]             uc2rb_desc_6_txn_type_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_0_reg;
wire [31:0]             uc2rb_desc_6_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_10_reg;
wire [31:0]             uc2rb_desc_6_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_11_reg;
wire [31:0]             uc2rb_desc_6_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_12_reg;
wire [31:0]             uc2rb_desc_6_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_13_reg;
wire [31:0]             uc2rb_desc_6_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_14_reg;
wire [31:0]             uc2rb_desc_6_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_15_reg;
wire [31:0]             uc2rb_desc_6_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_1_reg;
wire [31:0]             uc2rb_desc_6_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_2_reg;
wire [31:0]             uc2rb_desc_6_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_3_reg;
wire [31:0]             uc2rb_desc_6_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_4_reg;
wire [31:0]             uc2rb_desc_6_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_5_reg;
wire [31:0]             uc2rb_desc_6_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_6_reg;
wire [31:0]             uc2rb_desc_6_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_7_reg;
wire [31:0]             uc2rb_desc_6_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_8_reg;
wire [31:0]             uc2rb_desc_6_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_6_wuser_9_reg;
wire [31:0]             uc2rb_desc_6_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_7_attr_reg;  
wire [31:0]             uc2rb_desc_7_attr_reg_we;
wire [31:0]             uc2rb_desc_7_axaddr_0_reg;
wire [31:0]             uc2rb_desc_7_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_7_axaddr_1_reg;
wire [31:0]             uc2rb_desc_7_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_7_axaddr_2_reg;
wire [31:0]             uc2rb_desc_7_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_7_axaddr_3_reg;
wire [31:0]             uc2rb_desc_7_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_7_axid_0_reg;
wire [31:0]             uc2rb_desc_7_axid_0_reg_we;
wire [31:0]             uc2rb_desc_7_axid_1_reg;
wire [31:0]             uc2rb_desc_7_axid_1_reg_we;
wire [31:0]             uc2rb_desc_7_axid_2_reg;
wire [31:0]             uc2rb_desc_7_axid_2_reg_we;
wire [31:0]             uc2rb_desc_7_axid_3_reg;
wire [31:0]             uc2rb_desc_7_axid_3_reg_we;
wire [31:0]             uc2rb_desc_7_axsize_reg;
wire [31:0]             uc2rb_desc_7_axsize_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_0_reg;
wire [31:0]             uc2rb_desc_7_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_10_reg;
wire [31:0]             uc2rb_desc_7_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_11_reg;
wire [31:0]             uc2rb_desc_7_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_12_reg;
wire [31:0]             uc2rb_desc_7_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_13_reg;
wire [31:0]             uc2rb_desc_7_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_14_reg;
wire [31:0]             uc2rb_desc_7_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_15_reg;
wire [31:0]             uc2rb_desc_7_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_1_reg;
wire [31:0]             uc2rb_desc_7_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_2_reg;
wire [31:0]             uc2rb_desc_7_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_3_reg;
wire [31:0]             uc2rb_desc_7_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_4_reg;
wire [31:0]             uc2rb_desc_7_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_5_reg;
wire [31:0]             uc2rb_desc_7_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_6_reg;
wire [31:0]             uc2rb_desc_7_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_7_reg;
wire [31:0]             uc2rb_desc_7_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_8_reg;
wire [31:0]             uc2rb_desc_7_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_7_axuser_9_reg;
wire [31:0]             uc2rb_desc_7_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_7_data_offset_reg;
wire [31:0]             uc2rb_desc_7_data_offset_reg_we;
wire [31:0]             uc2rb_desc_7_size_reg;  
wire [31:0]             uc2rb_desc_7_size_reg_we;
wire [31:0]             uc2rb_desc_7_txn_type_reg;
wire [31:0]             uc2rb_desc_7_txn_type_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_0_reg;
wire [31:0]             uc2rb_desc_7_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_10_reg;
wire [31:0]             uc2rb_desc_7_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_11_reg;
wire [31:0]             uc2rb_desc_7_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_12_reg;
wire [31:0]             uc2rb_desc_7_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_13_reg;
wire [31:0]             uc2rb_desc_7_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_14_reg;
wire [31:0]             uc2rb_desc_7_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_15_reg;
wire [31:0]             uc2rb_desc_7_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_1_reg;
wire [31:0]             uc2rb_desc_7_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_2_reg;
wire [31:0]             uc2rb_desc_7_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_3_reg;
wire [31:0]             uc2rb_desc_7_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_4_reg;
wire [31:0]             uc2rb_desc_7_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_5_reg;
wire [31:0]             uc2rb_desc_7_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_6_reg;
wire [31:0]             uc2rb_desc_7_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_7_reg;
wire [31:0]             uc2rb_desc_7_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_8_reg;
wire [31:0]             uc2rb_desc_7_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_7_wuser_9_reg;
wire [31:0]             uc2rb_desc_7_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_8_attr_reg;  
wire [31:0]             uc2rb_desc_8_attr_reg_we;
wire [31:0]             uc2rb_desc_8_axaddr_0_reg;
wire [31:0]             uc2rb_desc_8_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_8_axaddr_1_reg;
wire [31:0]             uc2rb_desc_8_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_8_axaddr_2_reg;
wire [31:0]             uc2rb_desc_8_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_8_axaddr_3_reg;
wire [31:0]             uc2rb_desc_8_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_8_axid_0_reg;
wire [31:0]             uc2rb_desc_8_axid_0_reg_we;
wire [31:0]             uc2rb_desc_8_axid_1_reg;
wire [31:0]             uc2rb_desc_8_axid_1_reg_we;
wire [31:0]             uc2rb_desc_8_axid_2_reg;
wire [31:0]             uc2rb_desc_8_axid_2_reg_we;
wire [31:0]             uc2rb_desc_8_axid_3_reg;
wire [31:0]             uc2rb_desc_8_axid_3_reg_we;
wire [31:0]             uc2rb_desc_8_axsize_reg;
wire [31:0]             uc2rb_desc_8_axsize_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_0_reg;
wire [31:0]             uc2rb_desc_8_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_10_reg;
wire [31:0]             uc2rb_desc_8_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_11_reg;
wire [31:0]             uc2rb_desc_8_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_12_reg;
wire [31:0]             uc2rb_desc_8_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_13_reg;
wire [31:0]             uc2rb_desc_8_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_14_reg;
wire [31:0]             uc2rb_desc_8_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_15_reg;
wire [31:0]             uc2rb_desc_8_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_1_reg;
wire [31:0]             uc2rb_desc_8_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_2_reg;
wire [31:0]             uc2rb_desc_8_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_3_reg;
wire [31:0]             uc2rb_desc_8_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_4_reg;
wire [31:0]             uc2rb_desc_8_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_5_reg;
wire [31:0]             uc2rb_desc_8_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_6_reg;
wire [31:0]             uc2rb_desc_8_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_7_reg;
wire [31:0]             uc2rb_desc_8_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_8_reg;
wire [31:0]             uc2rb_desc_8_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_8_axuser_9_reg;
wire [31:0]             uc2rb_desc_8_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_8_data_offset_reg;
wire [31:0]             uc2rb_desc_8_data_offset_reg_we;
wire [31:0]             uc2rb_desc_8_size_reg;  
wire [31:0]             uc2rb_desc_8_size_reg_we;
wire [31:0]             uc2rb_desc_8_txn_type_reg;
wire [31:0]             uc2rb_desc_8_txn_type_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_0_reg;
wire [31:0]             uc2rb_desc_8_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_10_reg;
wire [31:0]             uc2rb_desc_8_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_11_reg;
wire [31:0]             uc2rb_desc_8_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_12_reg;
wire [31:0]             uc2rb_desc_8_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_13_reg;
wire [31:0]             uc2rb_desc_8_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_14_reg;
wire [31:0]             uc2rb_desc_8_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_15_reg;
wire [31:0]             uc2rb_desc_8_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_1_reg;
wire [31:0]             uc2rb_desc_8_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_2_reg;
wire [31:0]             uc2rb_desc_8_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_3_reg;
wire [31:0]             uc2rb_desc_8_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_4_reg;
wire [31:0]             uc2rb_desc_8_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_5_reg;
wire [31:0]             uc2rb_desc_8_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_6_reg;
wire [31:0]             uc2rb_desc_8_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_7_reg;
wire [31:0]             uc2rb_desc_8_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_8_reg;
wire [31:0]             uc2rb_desc_8_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_8_wuser_9_reg;
wire [31:0]             uc2rb_desc_8_wuser_9_reg_we;
wire [31:0]             uc2rb_desc_9_attr_reg;  
wire [31:0]             uc2rb_desc_9_attr_reg_we;
wire [31:0]             uc2rb_desc_9_axaddr_0_reg;
wire [31:0]             uc2rb_desc_9_axaddr_0_reg_we;
wire [31:0]             uc2rb_desc_9_axaddr_1_reg;
wire [31:0]             uc2rb_desc_9_axaddr_1_reg_we;
wire [31:0]             uc2rb_desc_9_axaddr_2_reg;
wire [31:0]             uc2rb_desc_9_axaddr_2_reg_we;
wire [31:0]             uc2rb_desc_9_axaddr_3_reg;
wire [31:0]             uc2rb_desc_9_axaddr_3_reg_we;
wire [31:0]             uc2rb_desc_9_axid_0_reg;
wire [31:0]             uc2rb_desc_9_axid_0_reg_we;
wire [31:0]             uc2rb_desc_9_axid_1_reg;
wire [31:0]             uc2rb_desc_9_axid_1_reg_we;
wire [31:0]             uc2rb_desc_9_axid_2_reg;
wire [31:0]             uc2rb_desc_9_axid_2_reg_we;
wire [31:0]             uc2rb_desc_9_axid_3_reg;
wire [31:0]             uc2rb_desc_9_axid_3_reg_we;
wire [31:0]             uc2rb_desc_9_axsize_reg;
wire [31:0]             uc2rb_desc_9_axsize_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_0_reg;
wire [31:0]             uc2rb_desc_9_axuser_0_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_10_reg;
wire [31:0]             uc2rb_desc_9_axuser_10_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_11_reg;
wire [31:0]             uc2rb_desc_9_axuser_11_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_12_reg;
wire [31:0]             uc2rb_desc_9_axuser_12_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_13_reg;
wire [31:0]             uc2rb_desc_9_axuser_13_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_14_reg;
wire [31:0]             uc2rb_desc_9_axuser_14_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_15_reg;
wire [31:0]             uc2rb_desc_9_axuser_15_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_1_reg;
wire [31:0]             uc2rb_desc_9_axuser_1_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_2_reg;
wire [31:0]             uc2rb_desc_9_axuser_2_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_3_reg;
wire [31:0]             uc2rb_desc_9_axuser_3_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_4_reg;
wire [31:0]             uc2rb_desc_9_axuser_4_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_5_reg;
wire [31:0]             uc2rb_desc_9_axuser_5_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_6_reg;
wire [31:0]             uc2rb_desc_9_axuser_6_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_7_reg;
wire [31:0]             uc2rb_desc_9_axuser_7_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_8_reg;
wire [31:0]             uc2rb_desc_9_axuser_8_reg_we;
wire [31:0]             uc2rb_desc_9_axuser_9_reg;
wire [31:0]             uc2rb_desc_9_axuser_9_reg_we;
wire [31:0]             uc2rb_desc_9_data_offset_reg;
wire [31:0]             uc2rb_desc_9_data_offset_reg_we;
wire [31:0]             uc2rb_desc_9_size_reg;  
wire [31:0]             uc2rb_desc_9_size_reg_we;
wire [31:0]             uc2rb_desc_9_txn_type_reg;
wire [31:0]             uc2rb_desc_9_txn_type_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_0_reg;
wire [31:0]             uc2rb_desc_9_wuser_0_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_10_reg;
wire [31:0]             uc2rb_desc_9_wuser_10_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_11_reg;
wire [31:0]             uc2rb_desc_9_wuser_11_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_12_reg;
wire [31:0]             uc2rb_desc_9_wuser_12_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_13_reg;
wire [31:0]             uc2rb_desc_9_wuser_13_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_14_reg;
wire [31:0]             uc2rb_desc_9_wuser_14_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_15_reg;
wire [31:0]             uc2rb_desc_9_wuser_15_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_1_reg;
wire [31:0]             uc2rb_desc_9_wuser_1_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_2_reg;
wire [31:0]             uc2rb_desc_9_wuser_2_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_3_reg;
wire [31:0]             uc2rb_desc_9_wuser_3_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_4_reg;
wire [31:0]             uc2rb_desc_9_wuser_4_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_5_reg;
wire [31:0]             uc2rb_desc_9_wuser_5_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_6_reg;
wire [31:0]             uc2rb_desc_9_wuser_6_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_7_reg;
wire [31:0]             uc2rb_desc_9_wuser_7_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_8_reg;
wire [31:0]             uc2rb_desc_9_wuser_8_reg_we;
wire [31:0]             uc2rb_desc_9_wuser_9_reg;
wire [31:0]             uc2rb_desc_9_wuser_9_reg_we;
wire [31:0]             uc2rb_intr_error_status_reg;
wire [31:0]             uc2rb_intr_error_status_reg_we;
wire [31:0]             uc2rb_intr_txn_avail_status_reg;
wire [31:0]             uc2rb_intr_txn_avail_status_reg_we;
wire [31:0]             uc2rb_intr_comp_status_reg;
wire [31:0]             uc2rb_intr_comp_status_reg_we;
wire [31:0]             uc2rb_ownership_reg;    
wire [31:0]             uc2rb_ownership_reg_we; 
wire [(`CLOG2((RAM_SIZE*8)/S_AXI_USR_DATA_WIDTH))-1:0] uc2rb_rd_addr;
wire [S_AXI_USR_DATA_WIDTH-1:0]                        rb2uc_rd_data;
wire [31:0]             uc2rb_status_busy_reg;  
wire [31:0]             uc2rb_status_busy_reg_we;
wire [31:0]             uc2rb_resp_fifo_free_level_reg;  
wire [31:0]             uc2rb_resp_fifo_free_level_reg_we;
wire [(`CLOG2((RAM_SIZE*8)/S_AXI_USR_DATA_WIDTH))-1:0] uc2rb_wr_addr;
wire [(S_AXI_USR_DATA_WIDTH/8)-1:0] uc2rb_wr_bwe;
wire [S_AXI_USR_DATA_WIDTH-1:0] uc2rb_wr_data;  
wire                    uc2rb_wr_we;            
wire [(S_AXI_USR_DATA_WIDTH/8)-1:0] uc2rb_wr_wstrb;
wire [31:0]             version_reg;            
// End of automatics

   user_slave_control #(
                            .EN_INTFS_AXI4          (EN_INTFS_AXI4       ),
                            .EN_INTFS_AXI4LITE      (EN_INTFS_AXI4LITE   ),
                            .EN_INTFS_AXI3          (EN_INTFS_AXI3       ),
                            .S_AXI_USR_ADDR_WIDTH   (S_AXI_USR_ADDR_WIDTH), 
                            .S_AXI_USR_DATA_WIDTH   (S_AXI_USR_DATA_WIDTH), 
                            .S_AXI_USR_ID_WIDTH     (S_AXI_USR_ID_WIDTH  ), 
                            .S_AXI_USR_AWUSER_WIDTH (S_AXI_USR_AWUSER_WIDTH),
                            .S_AXI_USR_WUSER_WIDTH  (S_AXI_USR_WUSER_WIDTH),
                            .S_AXI_USR_BUSER_WIDTH  (S_AXI_USR_BUSER_WIDTH),
                            .S_AXI_USR_ARUSER_WIDTH (S_AXI_USR_ARUSER_WIDTH),
                            .S_AXI_USR_RUSER_WIDTH  (S_AXI_USR_RUSER_WIDTH),
                            .RAM_SIZE               (RAM_SIZE            ), 
                            .MAX_DESC               (MAX_DESC            ),
	                    .FORCE_RESP_ORDER       (FORCE_RESP_ORDER)
                        )
   

user_slave_control_inst (/*AUTO*INST*/
                                               // Outputs
                                               .uc2rb_intr_error_status_reg(uc2rb_intr_error_status_reg),
                                               .uc2rb_ownership_reg(uc2rb_ownership_reg),
                                               .uc2rb_intr_txn_avail_status_reg(uc2rb_intr_txn_avail_status_reg),
                                               .uc2rb_intr_comp_status_reg(uc2rb_intr_comp_status_reg),
                                               .uc2rb_status_busy_reg(uc2rb_status_busy_reg),
                                               .uc2rb_resp_fifo_free_level_reg(uc2rb_resp_fifo_free_level_reg),
                                               .uc2rb_desc_0_txn_type_reg(uc2rb_desc_0_txn_type_reg),
                                               .uc2rb_desc_0_size_reg(uc2rb_desc_0_size_reg),
                                               .uc2rb_desc_0_data_offset_reg(uc2rb_desc_0_data_offset_reg),
                                               .uc2rb_desc_0_axsize_reg(uc2rb_desc_0_axsize_reg),
                                               .uc2rb_desc_0_attr_reg(uc2rb_desc_0_attr_reg),
                                               .uc2rb_desc_0_axaddr_0_reg(uc2rb_desc_0_axaddr_0_reg),
                                               .uc2rb_desc_0_axaddr_1_reg(uc2rb_desc_0_axaddr_1_reg),
                                               .uc2rb_desc_0_axaddr_2_reg(uc2rb_desc_0_axaddr_2_reg),
                                               .uc2rb_desc_0_axaddr_3_reg(uc2rb_desc_0_axaddr_3_reg),
                                               .uc2rb_desc_0_axid_0_reg(uc2rb_desc_0_axid_0_reg),
                                               .uc2rb_desc_0_axid_1_reg(uc2rb_desc_0_axid_1_reg),
                                               .uc2rb_desc_0_axid_2_reg(uc2rb_desc_0_axid_2_reg),
                                               .uc2rb_desc_0_axid_3_reg(uc2rb_desc_0_axid_3_reg),
                                               .uc2rb_desc_0_axuser_0_reg(uc2rb_desc_0_axuser_0_reg),
                                               .uc2rb_desc_0_axuser_1_reg(uc2rb_desc_0_axuser_1_reg),
                                               .uc2rb_desc_0_axuser_2_reg(uc2rb_desc_0_axuser_2_reg),
                                               .uc2rb_desc_0_axuser_3_reg(uc2rb_desc_0_axuser_3_reg),
                                               .uc2rb_desc_0_axuser_4_reg(uc2rb_desc_0_axuser_4_reg),
                                               .uc2rb_desc_0_axuser_5_reg(uc2rb_desc_0_axuser_5_reg),
                                               .uc2rb_desc_0_axuser_6_reg(uc2rb_desc_0_axuser_6_reg),
                                               .uc2rb_desc_0_axuser_7_reg(uc2rb_desc_0_axuser_7_reg),
                                               .uc2rb_desc_0_axuser_8_reg(uc2rb_desc_0_axuser_8_reg),
                                               .uc2rb_desc_0_axuser_9_reg(uc2rb_desc_0_axuser_9_reg),
                                               .uc2rb_desc_0_axuser_10_reg(uc2rb_desc_0_axuser_10_reg),
                                               .uc2rb_desc_0_axuser_11_reg(uc2rb_desc_0_axuser_11_reg),
                                               .uc2rb_desc_0_axuser_12_reg(uc2rb_desc_0_axuser_12_reg),
                                               .uc2rb_desc_0_axuser_13_reg(uc2rb_desc_0_axuser_13_reg),
                                               .uc2rb_desc_0_axuser_14_reg(uc2rb_desc_0_axuser_14_reg),
                                               .uc2rb_desc_0_axuser_15_reg(uc2rb_desc_0_axuser_15_reg),
                                               .uc2rb_desc_0_wuser_0_reg(uc2rb_desc_0_wuser_0_reg),
                                               .uc2rb_desc_0_wuser_1_reg(uc2rb_desc_0_wuser_1_reg),
                                               .uc2rb_desc_0_wuser_2_reg(uc2rb_desc_0_wuser_2_reg),
                                               .uc2rb_desc_0_wuser_3_reg(uc2rb_desc_0_wuser_3_reg),
                                               .uc2rb_desc_0_wuser_4_reg(uc2rb_desc_0_wuser_4_reg),
                                               .uc2rb_desc_0_wuser_5_reg(uc2rb_desc_0_wuser_5_reg),
                                               .uc2rb_desc_0_wuser_6_reg(uc2rb_desc_0_wuser_6_reg),
                                               .uc2rb_desc_0_wuser_7_reg(uc2rb_desc_0_wuser_7_reg),
                                               .uc2rb_desc_0_wuser_8_reg(uc2rb_desc_0_wuser_8_reg),
                                               .uc2rb_desc_0_wuser_9_reg(uc2rb_desc_0_wuser_9_reg),
                                               .uc2rb_desc_0_wuser_10_reg(uc2rb_desc_0_wuser_10_reg),
                                               .uc2rb_desc_0_wuser_11_reg(uc2rb_desc_0_wuser_11_reg),
                                               .uc2rb_desc_0_wuser_12_reg(uc2rb_desc_0_wuser_12_reg),
                                               .uc2rb_desc_0_wuser_13_reg(uc2rb_desc_0_wuser_13_reg),
                                               .uc2rb_desc_0_wuser_14_reg(uc2rb_desc_0_wuser_14_reg),
                                               .uc2rb_desc_0_wuser_15_reg(uc2rb_desc_0_wuser_15_reg),
                                               .uc2rb_desc_1_txn_type_reg(uc2rb_desc_1_txn_type_reg),
                                               .uc2rb_desc_1_size_reg(uc2rb_desc_1_size_reg),
                                               .uc2rb_desc_1_data_offset_reg(uc2rb_desc_1_data_offset_reg),
                                               .uc2rb_desc_1_axsize_reg(uc2rb_desc_1_axsize_reg),
                                               .uc2rb_desc_1_attr_reg(uc2rb_desc_1_attr_reg),
                                               .uc2rb_desc_1_axaddr_0_reg(uc2rb_desc_1_axaddr_0_reg),
                                               .uc2rb_desc_1_axaddr_1_reg(uc2rb_desc_1_axaddr_1_reg),
                                               .uc2rb_desc_1_axaddr_2_reg(uc2rb_desc_1_axaddr_2_reg),
                                               .uc2rb_desc_1_axaddr_3_reg(uc2rb_desc_1_axaddr_3_reg),
                                               .uc2rb_desc_1_axid_0_reg(uc2rb_desc_1_axid_0_reg),
                                               .uc2rb_desc_1_axid_1_reg(uc2rb_desc_1_axid_1_reg),
                                               .uc2rb_desc_1_axid_2_reg(uc2rb_desc_1_axid_2_reg),
                                               .uc2rb_desc_1_axid_3_reg(uc2rb_desc_1_axid_3_reg),
                                               .uc2rb_desc_1_axuser_0_reg(uc2rb_desc_1_axuser_0_reg),
                                               .uc2rb_desc_1_axuser_1_reg(uc2rb_desc_1_axuser_1_reg),
                                               .uc2rb_desc_1_axuser_2_reg(uc2rb_desc_1_axuser_2_reg),
                                               .uc2rb_desc_1_axuser_3_reg(uc2rb_desc_1_axuser_3_reg),
                                               .uc2rb_desc_1_axuser_4_reg(uc2rb_desc_1_axuser_4_reg),
                                               .uc2rb_desc_1_axuser_5_reg(uc2rb_desc_1_axuser_5_reg),
                                               .uc2rb_desc_1_axuser_6_reg(uc2rb_desc_1_axuser_6_reg),
                                               .uc2rb_desc_1_axuser_7_reg(uc2rb_desc_1_axuser_7_reg),
                                               .uc2rb_desc_1_axuser_8_reg(uc2rb_desc_1_axuser_8_reg),
                                               .uc2rb_desc_1_axuser_9_reg(uc2rb_desc_1_axuser_9_reg),
                                               .uc2rb_desc_1_axuser_10_reg(uc2rb_desc_1_axuser_10_reg),
                                               .uc2rb_desc_1_axuser_11_reg(uc2rb_desc_1_axuser_11_reg),
                                               .uc2rb_desc_1_axuser_12_reg(uc2rb_desc_1_axuser_12_reg),
                                               .uc2rb_desc_1_axuser_13_reg(uc2rb_desc_1_axuser_13_reg),
                                               .uc2rb_desc_1_axuser_14_reg(uc2rb_desc_1_axuser_14_reg),
                                               .uc2rb_desc_1_axuser_15_reg(uc2rb_desc_1_axuser_15_reg),
                                               .uc2rb_desc_1_wuser_0_reg(uc2rb_desc_1_wuser_0_reg),
                                               .uc2rb_desc_1_wuser_1_reg(uc2rb_desc_1_wuser_1_reg),
                                               .uc2rb_desc_1_wuser_2_reg(uc2rb_desc_1_wuser_2_reg),
                                               .uc2rb_desc_1_wuser_3_reg(uc2rb_desc_1_wuser_3_reg),
                                               .uc2rb_desc_1_wuser_4_reg(uc2rb_desc_1_wuser_4_reg),
                                               .uc2rb_desc_1_wuser_5_reg(uc2rb_desc_1_wuser_5_reg),
                                               .uc2rb_desc_1_wuser_6_reg(uc2rb_desc_1_wuser_6_reg),
                                               .uc2rb_desc_1_wuser_7_reg(uc2rb_desc_1_wuser_7_reg),
                                               .uc2rb_desc_1_wuser_8_reg(uc2rb_desc_1_wuser_8_reg),
                                               .uc2rb_desc_1_wuser_9_reg(uc2rb_desc_1_wuser_9_reg),
                                               .uc2rb_desc_1_wuser_10_reg(uc2rb_desc_1_wuser_10_reg),
                                               .uc2rb_desc_1_wuser_11_reg(uc2rb_desc_1_wuser_11_reg),
                                               .uc2rb_desc_1_wuser_12_reg(uc2rb_desc_1_wuser_12_reg),
                                               .uc2rb_desc_1_wuser_13_reg(uc2rb_desc_1_wuser_13_reg),
                                               .uc2rb_desc_1_wuser_14_reg(uc2rb_desc_1_wuser_14_reg),
                                               .uc2rb_desc_1_wuser_15_reg(uc2rb_desc_1_wuser_15_reg),
                                               .uc2rb_desc_2_txn_type_reg(uc2rb_desc_2_txn_type_reg),
                                               .uc2rb_desc_2_size_reg(uc2rb_desc_2_size_reg),
                                               .uc2rb_desc_2_data_offset_reg(uc2rb_desc_2_data_offset_reg),
                                               .uc2rb_desc_2_axsize_reg(uc2rb_desc_2_axsize_reg),
                                               .uc2rb_desc_2_attr_reg(uc2rb_desc_2_attr_reg),
                                               .uc2rb_desc_2_axaddr_0_reg(uc2rb_desc_2_axaddr_0_reg),
                                               .uc2rb_desc_2_axaddr_1_reg(uc2rb_desc_2_axaddr_1_reg),
                                               .uc2rb_desc_2_axaddr_2_reg(uc2rb_desc_2_axaddr_2_reg),
                                               .uc2rb_desc_2_axaddr_3_reg(uc2rb_desc_2_axaddr_3_reg),
                                               .uc2rb_desc_2_axid_0_reg(uc2rb_desc_2_axid_0_reg),
                                               .uc2rb_desc_2_axid_1_reg(uc2rb_desc_2_axid_1_reg),
                                               .uc2rb_desc_2_axid_2_reg(uc2rb_desc_2_axid_2_reg),
                                               .uc2rb_desc_2_axid_3_reg(uc2rb_desc_2_axid_3_reg),
                                               .uc2rb_desc_2_axuser_0_reg(uc2rb_desc_2_axuser_0_reg),
                                               .uc2rb_desc_2_axuser_1_reg(uc2rb_desc_2_axuser_1_reg),
                                               .uc2rb_desc_2_axuser_2_reg(uc2rb_desc_2_axuser_2_reg),
                                               .uc2rb_desc_2_axuser_3_reg(uc2rb_desc_2_axuser_3_reg),
                                               .uc2rb_desc_2_axuser_4_reg(uc2rb_desc_2_axuser_4_reg),
                                               .uc2rb_desc_2_axuser_5_reg(uc2rb_desc_2_axuser_5_reg),
                                               .uc2rb_desc_2_axuser_6_reg(uc2rb_desc_2_axuser_6_reg),
                                               .uc2rb_desc_2_axuser_7_reg(uc2rb_desc_2_axuser_7_reg),
                                               .uc2rb_desc_2_axuser_8_reg(uc2rb_desc_2_axuser_8_reg),
                                               .uc2rb_desc_2_axuser_9_reg(uc2rb_desc_2_axuser_9_reg),
                                               .uc2rb_desc_2_axuser_10_reg(uc2rb_desc_2_axuser_10_reg),
                                               .uc2rb_desc_2_axuser_11_reg(uc2rb_desc_2_axuser_11_reg),
                                               .uc2rb_desc_2_axuser_12_reg(uc2rb_desc_2_axuser_12_reg),
                                               .uc2rb_desc_2_axuser_13_reg(uc2rb_desc_2_axuser_13_reg),
                                               .uc2rb_desc_2_axuser_14_reg(uc2rb_desc_2_axuser_14_reg),
                                               .uc2rb_desc_2_axuser_15_reg(uc2rb_desc_2_axuser_15_reg),
                                               .uc2rb_desc_2_wuser_0_reg(uc2rb_desc_2_wuser_0_reg),
                                               .uc2rb_desc_2_wuser_1_reg(uc2rb_desc_2_wuser_1_reg),
                                               .uc2rb_desc_2_wuser_2_reg(uc2rb_desc_2_wuser_2_reg),
                                               .uc2rb_desc_2_wuser_3_reg(uc2rb_desc_2_wuser_3_reg),
                                               .uc2rb_desc_2_wuser_4_reg(uc2rb_desc_2_wuser_4_reg),
                                               .uc2rb_desc_2_wuser_5_reg(uc2rb_desc_2_wuser_5_reg),
                                               .uc2rb_desc_2_wuser_6_reg(uc2rb_desc_2_wuser_6_reg),
                                               .uc2rb_desc_2_wuser_7_reg(uc2rb_desc_2_wuser_7_reg),
                                               .uc2rb_desc_2_wuser_8_reg(uc2rb_desc_2_wuser_8_reg),
                                               .uc2rb_desc_2_wuser_9_reg(uc2rb_desc_2_wuser_9_reg),
                                               .uc2rb_desc_2_wuser_10_reg(uc2rb_desc_2_wuser_10_reg),
                                               .uc2rb_desc_2_wuser_11_reg(uc2rb_desc_2_wuser_11_reg),
                                               .uc2rb_desc_2_wuser_12_reg(uc2rb_desc_2_wuser_12_reg),
                                               .uc2rb_desc_2_wuser_13_reg(uc2rb_desc_2_wuser_13_reg),
                                               .uc2rb_desc_2_wuser_14_reg(uc2rb_desc_2_wuser_14_reg),
                                               .uc2rb_desc_2_wuser_15_reg(uc2rb_desc_2_wuser_15_reg),
                                               .uc2rb_desc_3_txn_type_reg(uc2rb_desc_3_txn_type_reg),
                                               .uc2rb_desc_3_size_reg(uc2rb_desc_3_size_reg),
                                               .uc2rb_desc_3_data_offset_reg(uc2rb_desc_3_data_offset_reg),
                                               .uc2rb_desc_3_axsize_reg(uc2rb_desc_3_axsize_reg),
                                               .uc2rb_desc_3_attr_reg(uc2rb_desc_3_attr_reg),
                                               .uc2rb_desc_3_axaddr_0_reg(uc2rb_desc_3_axaddr_0_reg),
                                               .uc2rb_desc_3_axaddr_1_reg(uc2rb_desc_3_axaddr_1_reg),
                                               .uc2rb_desc_3_axaddr_2_reg(uc2rb_desc_3_axaddr_2_reg),
                                               .uc2rb_desc_3_axaddr_3_reg(uc2rb_desc_3_axaddr_3_reg),
                                               .uc2rb_desc_3_axid_0_reg(uc2rb_desc_3_axid_0_reg),
                                               .uc2rb_desc_3_axid_1_reg(uc2rb_desc_3_axid_1_reg),
                                               .uc2rb_desc_3_axid_2_reg(uc2rb_desc_3_axid_2_reg),
                                               .uc2rb_desc_3_axid_3_reg(uc2rb_desc_3_axid_3_reg),
                                               .uc2rb_desc_3_axuser_0_reg(uc2rb_desc_3_axuser_0_reg),
                                               .uc2rb_desc_3_axuser_1_reg(uc2rb_desc_3_axuser_1_reg),
                                               .uc2rb_desc_3_axuser_2_reg(uc2rb_desc_3_axuser_2_reg),
                                               .uc2rb_desc_3_axuser_3_reg(uc2rb_desc_3_axuser_3_reg),
                                               .uc2rb_desc_3_axuser_4_reg(uc2rb_desc_3_axuser_4_reg),
                                               .uc2rb_desc_3_axuser_5_reg(uc2rb_desc_3_axuser_5_reg),
                                               .uc2rb_desc_3_axuser_6_reg(uc2rb_desc_3_axuser_6_reg),
                                               .uc2rb_desc_3_axuser_7_reg(uc2rb_desc_3_axuser_7_reg),
                                               .uc2rb_desc_3_axuser_8_reg(uc2rb_desc_3_axuser_8_reg),
                                               .uc2rb_desc_3_axuser_9_reg(uc2rb_desc_3_axuser_9_reg),
                                               .uc2rb_desc_3_axuser_10_reg(uc2rb_desc_3_axuser_10_reg),
                                               .uc2rb_desc_3_axuser_11_reg(uc2rb_desc_3_axuser_11_reg),
                                               .uc2rb_desc_3_axuser_12_reg(uc2rb_desc_3_axuser_12_reg),
                                               .uc2rb_desc_3_axuser_13_reg(uc2rb_desc_3_axuser_13_reg),
                                               .uc2rb_desc_3_axuser_14_reg(uc2rb_desc_3_axuser_14_reg),
                                               .uc2rb_desc_3_axuser_15_reg(uc2rb_desc_3_axuser_15_reg),
                                               .uc2rb_desc_3_wuser_0_reg(uc2rb_desc_3_wuser_0_reg),
                                               .uc2rb_desc_3_wuser_1_reg(uc2rb_desc_3_wuser_1_reg),
                                               .uc2rb_desc_3_wuser_2_reg(uc2rb_desc_3_wuser_2_reg),
                                               .uc2rb_desc_3_wuser_3_reg(uc2rb_desc_3_wuser_3_reg),
                                               .uc2rb_desc_3_wuser_4_reg(uc2rb_desc_3_wuser_4_reg),
                                               .uc2rb_desc_3_wuser_5_reg(uc2rb_desc_3_wuser_5_reg),
                                               .uc2rb_desc_3_wuser_6_reg(uc2rb_desc_3_wuser_6_reg),
                                               .uc2rb_desc_3_wuser_7_reg(uc2rb_desc_3_wuser_7_reg),
                                               .uc2rb_desc_3_wuser_8_reg(uc2rb_desc_3_wuser_8_reg),
                                               .uc2rb_desc_3_wuser_9_reg(uc2rb_desc_3_wuser_9_reg),
                                               .uc2rb_desc_3_wuser_10_reg(uc2rb_desc_3_wuser_10_reg),
                                               .uc2rb_desc_3_wuser_11_reg(uc2rb_desc_3_wuser_11_reg),
                                               .uc2rb_desc_3_wuser_12_reg(uc2rb_desc_3_wuser_12_reg),
                                               .uc2rb_desc_3_wuser_13_reg(uc2rb_desc_3_wuser_13_reg),
                                               .uc2rb_desc_3_wuser_14_reg(uc2rb_desc_3_wuser_14_reg),
                                               .uc2rb_desc_3_wuser_15_reg(uc2rb_desc_3_wuser_15_reg),
                                               .uc2rb_desc_4_txn_type_reg(uc2rb_desc_4_txn_type_reg),
                                               .uc2rb_desc_4_size_reg(uc2rb_desc_4_size_reg),
                                               .uc2rb_desc_4_data_offset_reg(uc2rb_desc_4_data_offset_reg),
                                               .uc2rb_desc_4_axsize_reg(uc2rb_desc_4_axsize_reg),
                                               .uc2rb_desc_4_attr_reg(uc2rb_desc_4_attr_reg),
                                               .uc2rb_desc_4_axaddr_0_reg(uc2rb_desc_4_axaddr_0_reg),
                                               .uc2rb_desc_4_axaddr_1_reg(uc2rb_desc_4_axaddr_1_reg),
                                               .uc2rb_desc_4_axaddr_2_reg(uc2rb_desc_4_axaddr_2_reg),
                                               .uc2rb_desc_4_axaddr_3_reg(uc2rb_desc_4_axaddr_3_reg),
                                               .uc2rb_desc_4_axid_0_reg(uc2rb_desc_4_axid_0_reg),
                                               .uc2rb_desc_4_axid_1_reg(uc2rb_desc_4_axid_1_reg),
                                               .uc2rb_desc_4_axid_2_reg(uc2rb_desc_4_axid_2_reg),
                                               .uc2rb_desc_4_axid_3_reg(uc2rb_desc_4_axid_3_reg),
                                               .uc2rb_desc_4_axuser_0_reg(uc2rb_desc_4_axuser_0_reg),
                                               .uc2rb_desc_4_axuser_1_reg(uc2rb_desc_4_axuser_1_reg),
                                               .uc2rb_desc_4_axuser_2_reg(uc2rb_desc_4_axuser_2_reg),
                                               .uc2rb_desc_4_axuser_3_reg(uc2rb_desc_4_axuser_3_reg),
                                               .uc2rb_desc_4_axuser_4_reg(uc2rb_desc_4_axuser_4_reg),
                                               .uc2rb_desc_4_axuser_5_reg(uc2rb_desc_4_axuser_5_reg),
                                               .uc2rb_desc_4_axuser_6_reg(uc2rb_desc_4_axuser_6_reg),
                                               .uc2rb_desc_4_axuser_7_reg(uc2rb_desc_4_axuser_7_reg),
                                               .uc2rb_desc_4_axuser_8_reg(uc2rb_desc_4_axuser_8_reg),
                                               .uc2rb_desc_4_axuser_9_reg(uc2rb_desc_4_axuser_9_reg),
                                               .uc2rb_desc_4_axuser_10_reg(uc2rb_desc_4_axuser_10_reg),
                                               .uc2rb_desc_4_axuser_11_reg(uc2rb_desc_4_axuser_11_reg),
                                               .uc2rb_desc_4_axuser_12_reg(uc2rb_desc_4_axuser_12_reg),
                                               .uc2rb_desc_4_axuser_13_reg(uc2rb_desc_4_axuser_13_reg),
                                               .uc2rb_desc_4_axuser_14_reg(uc2rb_desc_4_axuser_14_reg),
                                               .uc2rb_desc_4_axuser_15_reg(uc2rb_desc_4_axuser_15_reg),
                                               .uc2rb_desc_4_wuser_0_reg(uc2rb_desc_4_wuser_0_reg),
                                               .uc2rb_desc_4_wuser_1_reg(uc2rb_desc_4_wuser_1_reg),
                                               .uc2rb_desc_4_wuser_2_reg(uc2rb_desc_4_wuser_2_reg),
                                               .uc2rb_desc_4_wuser_3_reg(uc2rb_desc_4_wuser_3_reg),
                                               .uc2rb_desc_4_wuser_4_reg(uc2rb_desc_4_wuser_4_reg),
                                               .uc2rb_desc_4_wuser_5_reg(uc2rb_desc_4_wuser_5_reg),
                                               .uc2rb_desc_4_wuser_6_reg(uc2rb_desc_4_wuser_6_reg),
                                               .uc2rb_desc_4_wuser_7_reg(uc2rb_desc_4_wuser_7_reg),
                                               .uc2rb_desc_4_wuser_8_reg(uc2rb_desc_4_wuser_8_reg),
                                               .uc2rb_desc_4_wuser_9_reg(uc2rb_desc_4_wuser_9_reg),
                                               .uc2rb_desc_4_wuser_10_reg(uc2rb_desc_4_wuser_10_reg),
                                               .uc2rb_desc_4_wuser_11_reg(uc2rb_desc_4_wuser_11_reg),
                                               .uc2rb_desc_4_wuser_12_reg(uc2rb_desc_4_wuser_12_reg),
                                               .uc2rb_desc_4_wuser_13_reg(uc2rb_desc_4_wuser_13_reg),
                                               .uc2rb_desc_4_wuser_14_reg(uc2rb_desc_4_wuser_14_reg),
                                               .uc2rb_desc_4_wuser_15_reg(uc2rb_desc_4_wuser_15_reg),
                                               .uc2rb_desc_5_txn_type_reg(uc2rb_desc_5_txn_type_reg),
                                               .uc2rb_desc_5_size_reg(uc2rb_desc_5_size_reg),
                                               .uc2rb_desc_5_data_offset_reg(uc2rb_desc_5_data_offset_reg),
                                               .uc2rb_desc_5_axsize_reg(uc2rb_desc_5_axsize_reg),
                                               .uc2rb_desc_5_attr_reg(uc2rb_desc_5_attr_reg),
                                               .uc2rb_desc_5_axaddr_0_reg(uc2rb_desc_5_axaddr_0_reg),
                                               .uc2rb_desc_5_axaddr_1_reg(uc2rb_desc_5_axaddr_1_reg),
                                               .uc2rb_desc_5_axaddr_2_reg(uc2rb_desc_5_axaddr_2_reg),
                                               .uc2rb_desc_5_axaddr_3_reg(uc2rb_desc_5_axaddr_3_reg),
                                               .uc2rb_desc_5_axid_0_reg(uc2rb_desc_5_axid_0_reg),
                                               .uc2rb_desc_5_axid_1_reg(uc2rb_desc_5_axid_1_reg),
                                               .uc2rb_desc_5_axid_2_reg(uc2rb_desc_5_axid_2_reg),
                                               .uc2rb_desc_5_axid_3_reg(uc2rb_desc_5_axid_3_reg),
                                               .uc2rb_desc_5_axuser_0_reg(uc2rb_desc_5_axuser_0_reg),
                                               .uc2rb_desc_5_axuser_1_reg(uc2rb_desc_5_axuser_1_reg),
                                               .uc2rb_desc_5_axuser_2_reg(uc2rb_desc_5_axuser_2_reg),
                                               .uc2rb_desc_5_axuser_3_reg(uc2rb_desc_5_axuser_3_reg),
                                               .uc2rb_desc_5_axuser_4_reg(uc2rb_desc_5_axuser_4_reg),
                                               .uc2rb_desc_5_axuser_5_reg(uc2rb_desc_5_axuser_5_reg),
                                               .uc2rb_desc_5_axuser_6_reg(uc2rb_desc_5_axuser_6_reg),
                                               .uc2rb_desc_5_axuser_7_reg(uc2rb_desc_5_axuser_7_reg),
                                               .uc2rb_desc_5_axuser_8_reg(uc2rb_desc_5_axuser_8_reg),
                                               .uc2rb_desc_5_axuser_9_reg(uc2rb_desc_5_axuser_9_reg),
                                               .uc2rb_desc_5_axuser_10_reg(uc2rb_desc_5_axuser_10_reg),
                                               .uc2rb_desc_5_axuser_11_reg(uc2rb_desc_5_axuser_11_reg),
                                               .uc2rb_desc_5_axuser_12_reg(uc2rb_desc_5_axuser_12_reg),
                                               .uc2rb_desc_5_axuser_13_reg(uc2rb_desc_5_axuser_13_reg),
                                               .uc2rb_desc_5_axuser_14_reg(uc2rb_desc_5_axuser_14_reg),
                                               .uc2rb_desc_5_axuser_15_reg(uc2rb_desc_5_axuser_15_reg),
                                               .uc2rb_desc_5_wuser_0_reg(uc2rb_desc_5_wuser_0_reg),
                                               .uc2rb_desc_5_wuser_1_reg(uc2rb_desc_5_wuser_1_reg),
                                               .uc2rb_desc_5_wuser_2_reg(uc2rb_desc_5_wuser_2_reg),
                                               .uc2rb_desc_5_wuser_3_reg(uc2rb_desc_5_wuser_3_reg),
                                               .uc2rb_desc_5_wuser_4_reg(uc2rb_desc_5_wuser_4_reg),
                                               .uc2rb_desc_5_wuser_5_reg(uc2rb_desc_5_wuser_5_reg),
                                               .uc2rb_desc_5_wuser_6_reg(uc2rb_desc_5_wuser_6_reg),
                                               .uc2rb_desc_5_wuser_7_reg(uc2rb_desc_5_wuser_7_reg),
                                               .uc2rb_desc_5_wuser_8_reg(uc2rb_desc_5_wuser_8_reg),
                                               .uc2rb_desc_5_wuser_9_reg(uc2rb_desc_5_wuser_9_reg),
                                               .uc2rb_desc_5_wuser_10_reg(uc2rb_desc_5_wuser_10_reg),
                                               .uc2rb_desc_5_wuser_11_reg(uc2rb_desc_5_wuser_11_reg),
                                               .uc2rb_desc_5_wuser_12_reg(uc2rb_desc_5_wuser_12_reg),
                                               .uc2rb_desc_5_wuser_13_reg(uc2rb_desc_5_wuser_13_reg),
                                               .uc2rb_desc_5_wuser_14_reg(uc2rb_desc_5_wuser_14_reg),
                                               .uc2rb_desc_5_wuser_15_reg(uc2rb_desc_5_wuser_15_reg),
                                               .uc2rb_desc_6_txn_type_reg(uc2rb_desc_6_txn_type_reg),
                                               .uc2rb_desc_6_size_reg(uc2rb_desc_6_size_reg),
                                               .uc2rb_desc_6_data_offset_reg(uc2rb_desc_6_data_offset_reg),
                                               .uc2rb_desc_6_axsize_reg(uc2rb_desc_6_axsize_reg),
                                               .uc2rb_desc_6_attr_reg(uc2rb_desc_6_attr_reg),
                                               .uc2rb_desc_6_axaddr_0_reg(uc2rb_desc_6_axaddr_0_reg),
                                               .uc2rb_desc_6_axaddr_1_reg(uc2rb_desc_6_axaddr_1_reg),
                                               .uc2rb_desc_6_axaddr_2_reg(uc2rb_desc_6_axaddr_2_reg),
                                               .uc2rb_desc_6_axaddr_3_reg(uc2rb_desc_6_axaddr_3_reg),
                                               .uc2rb_desc_6_axid_0_reg(uc2rb_desc_6_axid_0_reg),
                                               .uc2rb_desc_6_axid_1_reg(uc2rb_desc_6_axid_1_reg),
                                               .uc2rb_desc_6_axid_2_reg(uc2rb_desc_6_axid_2_reg),
                                               .uc2rb_desc_6_axid_3_reg(uc2rb_desc_6_axid_3_reg),
                                               .uc2rb_desc_6_axuser_0_reg(uc2rb_desc_6_axuser_0_reg),
                                               .uc2rb_desc_6_axuser_1_reg(uc2rb_desc_6_axuser_1_reg),
                                               .uc2rb_desc_6_axuser_2_reg(uc2rb_desc_6_axuser_2_reg),
                                               .uc2rb_desc_6_axuser_3_reg(uc2rb_desc_6_axuser_3_reg),
                                               .uc2rb_desc_6_axuser_4_reg(uc2rb_desc_6_axuser_4_reg),
                                               .uc2rb_desc_6_axuser_5_reg(uc2rb_desc_6_axuser_5_reg),
                                               .uc2rb_desc_6_axuser_6_reg(uc2rb_desc_6_axuser_6_reg),
                                               .uc2rb_desc_6_axuser_7_reg(uc2rb_desc_6_axuser_7_reg),
                                               .uc2rb_desc_6_axuser_8_reg(uc2rb_desc_6_axuser_8_reg),
                                               .uc2rb_desc_6_axuser_9_reg(uc2rb_desc_6_axuser_9_reg),
                                               .uc2rb_desc_6_axuser_10_reg(uc2rb_desc_6_axuser_10_reg),
                                               .uc2rb_desc_6_axuser_11_reg(uc2rb_desc_6_axuser_11_reg),
                                               .uc2rb_desc_6_axuser_12_reg(uc2rb_desc_6_axuser_12_reg),
                                               .uc2rb_desc_6_axuser_13_reg(uc2rb_desc_6_axuser_13_reg),
                                               .uc2rb_desc_6_axuser_14_reg(uc2rb_desc_6_axuser_14_reg),
                                               .uc2rb_desc_6_axuser_15_reg(uc2rb_desc_6_axuser_15_reg),
                                               .uc2rb_desc_6_wuser_0_reg(uc2rb_desc_6_wuser_0_reg),
                                               .uc2rb_desc_6_wuser_1_reg(uc2rb_desc_6_wuser_1_reg),
                                               .uc2rb_desc_6_wuser_2_reg(uc2rb_desc_6_wuser_2_reg),
                                               .uc2rb_desc_6_wuser_3_reg(uc2rb_desc_6_wuser_3_reg),
                                               .uc2rb_desc_6_wuser_4_reg(uc2rb_desc_6_wuser_4_reg),
                                               .uc2rb_desc_6_wuser_5_reg(uc2rb_desc_6_wuser_5_reg),
                                               .uc2rb_desc_6_wuser_6_reg(uc2rb_desc_6_wuser_6_reg),
                                               .uc2rb_desc_6_wuser_7_reg(uc2rb_desc_6_wuser_7_reg),
                                               .uc2rb_desc_6_wuser_8_reg(uc2rb_desc_6_wuser_8_reg),
                                               .uc2rb_desc_6_wuser_9_reg(uc2rb_desc_6_wuser_9_reg),
                                               .uc2rb_desc_6_wuser_10_reg(uc2rb_desc_6_wuser_10_reg),
                                               .uc2rb_desc_6_wuser_11_reg(uc2rb_desc_6_wuser_11_reg),
                                               .uc2rb_desc_6_wuser_12_reg(uc2rb_desc_6_wuser_12_reg),
                                               .uc2rb_desc_6_wuser_13_reg(uc2rb_desc_6_wuser_13_reg),
                                               .uc2rb_desc_6_wuser_14_reg(uc2rb_desc_6_wuser_14_reg),
                                               .uc2rb_desc_6_wuser_15_reg(uc2rb_desc_6_wuser_15_reg),
                                               .uc2rb_desc_7_txn_type_reg(uc2rb_desc_7_txn_type_reg),
                                               .uc2rb_desc_7_size_reg(uc2rb_desc_7_size_reg),
                                               .uc2rb_desc_7_data_offset_reg(uc2rb_desc_7_data_offset_reg),
                                               .uc2rb_desc_7_axsize_reg(uc2rb_desc_7_axsize_reg),
                                               .uc2rb_desc_7_attr_reg(uc2rb_desc_7_attr_reg),
                                               .uc2rb_desc_7_axaddr_0_reg(uc2rb_desc_7_axaddr_0_reg),
                                               .uc2rb_desc_7_axaddr_1_reg(uc2rb_desc_7_axaddr_1_reg),
                                               .uc2rb_desc_7_axaddr_2_reg(uc2rb_desc_7_axaddr_2_reg),
                                               .uc2rb_desc_7_axaddr_3_reg(uc2rb_desc_7_axaddr_3_reg),
                                               .uc2rb_desc_7_axid_0_reg(uc2rb_desc_7_axid_0_reg),
                                               .uc2rb_desc_7_axid_1_reg(uc2rb_desc_7_axid_1_reg),
                                               .uc2rb_desc_7_axid_2_reg(uc2rb_desc_7_axid_2_reg),
                                               .uc2rb_desc_7_axid_3_reg(uc2rb_desc_7_axid_3_reg),
                                               .uc2rb_desc_7_axuser_0_reg(uc2rb_desc_7_axuser_0_reg),
                                               .uc2rb_desc_7_axuser_1_reg(uc2rb_desc_7_axuser_1_reg),
                                               .uc2rb_desc_7_axuser_2_reg(uc2rb_desc_7_axuser_2_reg),
                                               .uc2rb_desc_7_axuser_3_reg(uc2rb_desc_7_axuser_3_reg),
                                               .uc2rb_desc_7_axuser_4_reg(uc2rb_desc_7_axuser_4_reg),
                                               .uc2rb_desc_7_axuser_5_reg(uc2rb_desc_7_axuser_5_reg),
                                               .uc2rb_desc_7_axuser_6_reg(uc2rb_desc_7_axuser_6_reg),
                                               .uc2rb_desc_7_axuser_7_reg(uc2rb_desc_7_axuser_7_reg),
                                               .uc2rb_desc_7_axuser_8_reg(uc2rb_desc_7_axuser_8_reg),
                                               .uc2rb_desc_7_axuser_9_reg(uc2rb_desc_7_axuser_9_reg),
                                               .uc2rb_desc_7_axuser_10_reg(uc2rb_desc_7_axuser_10_reg),
                                               .uc2rb_desc_7_axuser_11_reg(uc2rb_desc_7_axuser_11_reg),
                                               .uc2rb_desc_7_axuser_12_reg(uc2rb_desc_7_axuser_12_reg),
                                               .uc2rb_desc_7_axuser_13_reg(uc2rb_desc_7_axuser_13_reg),
                                               .uc2rb_desc_7_axuser_14_reg(uc2rb_desc_7_axuser_14_reg),
                                               .uc2rb_desc_7_axuser_15_reg(uc2rb_desc_7_axuser_15_reg),
                                               .uc2rb_desc_7_wuser_0_reg(uc2rb_desc_7_wuser_0_reg),
                                               .uc2rb_desc_7_wuser_1_reg(uc2rb_desc_7_wuser_1_reg),
                                               .uc2rb_desc_7_wuser_2_reg(uc2rb_desc_7_wuser_2_reg),
                                               .uc2rb_desc_7_wuser_3_reg(uc2rb_desc_7_wuser_3_reg),
                                               .uc2rb_desc_7_wuser_4_reg(uc2rb_desc_7_wuser_4_reg),
                                               .uc2rb_desc_7_wuser_5_reg(uc2rb_desc_7_wuser_5_reg),
                                               .uc2rb_desc_7_wuser_6_reg(uc2rb_desc_7_wuser_6_reg),
                                               .uc2rb_desc_7_wuser_7_reg(uc2rb_desc_7_wuser_7_reg),
                                               .uc2rb_desc_7_wuser_8_reg(uc2rb_desc_7_wuser_8_reg),
                                               .uc2rb_desc_7_wuser_9_reg(uc2rb_desc_7_wuser_9_reg),
                                               .uc2rb_desc_7_wuser_10_reg(uc2rb_desc_7_wuser_10_reg),
                                               .uc2rb_desc_7_wuser_11_reg(uc2rb_desc_7_wuser_11_reg),
                                               .uc2rb_desc_7_wuser_12_reg(uc2rb_desc_7_wuser_12_reg),
                                               .uc2rb_desc_7_wuser_13_reg(uc2rb_desc_7_wuser_13_reg),
                                               .uc2rb_desc_7_wuser_14_reg(uc2rb_desc_7_wuser_14_reg),
                                               .uc2rb_desc_7_wuser_15_reg(uc2rb_desc_7_wuser_15_reg),
                                               .uc2rb_desc_8_txn_type_reg(uc2rb_desc_8_txn_type_reg),
                                               .uc2rb_desc_8_size_reg(uc2rb_desc_8_size_reg),
                                               .uc2rb_desc_8_data_offset_reg(uc2rb_desc_8_data_offset_reg),
                                               .uc2rb_desc_8_axsize_reg(uc2rb_desc_8_axsize_reg),
                                               .uc2rb_desc_8_attr_reg(uc2rb_desc_8_attr_reg),
                                               .uc2rb_desc_8_axaddr_0_reg(uc2rb_desc_8_axaddr_0_reg),
                                               .uc2rb_desc_8_axaddr_1_reg(uc2rb_desc_8_axaddr_1_reg),
                                               .uc2rb_desc_8_axaddr_2_reg(uc2rb_desc_8_axaddr_2_reg),
                                               .uc2rb_desc_8_axaddr_3_reg(uc2rb_desc_8_axaddr_3_reg),
                                               .uc2rb_desc_8_axid_0_reg(uc2rb_desc_8_axid_0_reg),
                                               .uc2rb_desc_8_axid_1_reg(uc2rb_desc_8_axid_1_reg),
                                               .uc2rb_desc_8_axid_2_reg(uc2rb_desc_8_axid_2_reg),
                                               .uc2rb_desc_8_axid_3_reg(uc2rb_desc_8_axid_3_reg),
                                               .uc2rb_desc_8_axuser_0_reg(uc2rb_desc_8_axuser_0_reg),
                                               .uc2rb_desc_8_axuser_1_reg(uc2rb_desc_8_axuser_1_reg),
                                               .uc2rb_desc_8_axuser_2_reg(uc2rb_desc_8_axuser_2_reg),
                                               .uc2rb_desc_8_axuser_3_reg(uc2rb_desc_8_axuser_3_reg),
                                               .uc2rb_desc_8_axuser_4_reg(uc2rb_desc_8_axuser_4_reg),
                                               .uc2rb_desc_8_axuser_5_reg(uc2rb_desc_8_axuser_5_reg),
                                               .uc2rb_desc_8_axuser_6_reg(uc2rb_desc_8_axuser_6_reg),
                                               .uc2rb_desc_8_axuser_7_reg(uc2rb_desc_8_axuser_7_reg),
                                               .uc2rb_desc_8_axuser_8_reg(uc2rb_desc_8_axuser_8_reg),
                                               .uc2rb_desc_8_axuser_9_reg(uc2rb_desc_8_axuser_9_reg),
                                               .uc2rb_desc_8_axuser_10_reg(uc2rb_desc_8_axuser_10_reg),
                                               .uc2rb_desc_8_axuser_11_reg(uc2rb_desc_8_axuser_11_reg),
                                               .uc2rb_desc_8_axuser_12_reg(uc2rb_desc_8_axuser_12_reg),
                                               .uc2rb_desc_8_axuser_13_reg(uc2rb_desc_8_axuser_13_reg),
                                               .uc2rb_desc_8_axuser_14_reg(uc2rb_desc_8_axuser_14_reg),
                                               .uc2rb_desc_8_axuser_15_reg(uc2rb_desc_8_axuser_15_reg),
                                               .uc2rb_desc_8_wuser_0_reg(uc2rb_desc_8_wuser_0_reg),
                                               .uc2rb_desc_8_wuser_1_reg(uc2rb_desc_8_wuser_1_reg),
                                               .uc2rb_desc_8_wuser_2_reg(uc2rb_desc_8_wuser_2_reg),
                                               .uc2rb_desc_8_wuser_3_reg(uc2rb_desc_8_wuser_3_reg),
                                               .uc2rb_desc_8_wuser_4_reg(uc2rb_desc_8_wuser_4_reg),
                                               .uc2rb_desc_8_wuser_5_reg(uc2rb_desc_8_wuser_5_reg),
                                               .uc2rb_desc_8_wuser_6_reg(uc2rb_desc_8_wuser_6_reg),
                                               .uc2rb_desc_8_wuser_7_reg(uc2rb_desc_8_wuser_7_reg),
                                               .uc2rb_desc_8_wuser_8_reg(uc2rb_desc_8_wuser_8_reg),
                                               .uc2rb_desc_8_wuser_9_reg(uc2rb_desc_8_wuser_9_reg),
                                               .uc2rb_desc_8_wuser_10_reg(uc2rb_desc_8_wuser_10_reg),
                                               .uc2rb_desc_8_wuser_11_reg(uc2rb_desc_8_wuser_11_reg),
                                               .uc2rb_desc_8_wuser_12_reg(uc2rb_desc_8_wuser_12_reg),
                                               .uc2rb_desc_8_wuser_13_reg(uc2rb_desc_8_wuser_13_reg),
                                               .uc2rb_desc_8_wuser_14_reg(uc2rb_desc_8_wuser_14_reg),
                                               .uc2rb_desc_8_wuser_15_reg(uc2rb_desc_8_wuser_15_reg),
                                               .uc2rb_desc_9_txn_type_reg(uc2rb_desc_9_txn_type_reg),
                                               .uc2rb_desc_9_size_reg(uc2rb_desc_9_size_reg),
                                               .uc2rb_desc_9_data_offset_reg(uc2rb_desc_9_data_offset_reg),
                                               .uc2rb_desc_9_axsize_reg(uc2rb_desc_9_axsize_reg),
                                               .uc2rb_desc_9_attr_reg(uc2rb_desc_9_attr_reg),
                                               .uc2rb_desc_9_axaddr_0_reg(uc2rb_desc_9_axaddr_0_reg),
                                               .uc2rb_desc_9_axaddr_1_reg(uc2rb_desc_9_axaddr_1_reg),
                                               .uc2rb_desc_9_axaddr_2_reg(uc2rb_desc_9_axaddr_2_reg),
                                               .uc2rb_desc_9_axaddr_3_reg(uc2rb_desc_9_axaddr_3_reg),
                                               .uc2rb_desc_9_axid_0_reg(uc2rb_desc_9_axid_0_reg),
                                               .uc2rb_desc_9_axid_1_reg(uc2rb_desc_9_axid_1_reg),
                                               .uc2rb_desc_9_axid_2_reg(uc2rb_desc_9_axid_2_reg),
                                               .uc2rb_desc_9_axid_3_reg(uc2rb_desc_9_axid_3_reg),
                                               .uc2rb_desc_9_axuser_0_reg(uc2rb_desc_9_axuser_0_reg),
                                               .uc2rb_desc_9_axuser_1_reg(uc2rb_desc_9_axuser_1_reg),
                                               .uc2rb_desc_9_axuser_2_reg(uc2rb_desc_9_axuser_2_reg),
                                               .uc2rb_desc_9_axuser_3_reg(uc2rb_desc_9_axuser_3_reg),
                                               .uc2rb_desc_9_axuser_4_reg(uc2rb_desc_9_axuser_4_reg),
                                               .uc2rb_desc_9_axuser_5_reg(uc2rb_desc_9_axuser_5_reg),
                                               .uc2rb_desc_9_axuser_6_reg(uc2rb_desc_9_axuser_6_reg),
                                               .uc2rb_desc_9_axuser_7_reg(uc2rb_desc_9_axuser_7_reg),
                                               .uc2rb_desc_9_axuser_8_reg(uc2rb_desc_9_axuser_8_reg),
                                               .uc2rb_desc_9_axuser_9_reg(uc2rb_desc_9_axuser_9_reg),
                                               .uc2rb_desc_9_axuser_10_reg(uc2rb_desc_9_axuser_10_reg),
                                               .uc2rb_desc_9_axuser_11_reg(uc2rb_desc_9_axuser_11_reg),
                                               .uc2rb_desc_9_axuser_12_reg(uc2rb_desc_9_axuser_12_reg),
                                               .uc2rb_desc_9_axuser_13_reg(uc2rb_desc_9_axuser_13_reg),
                                               .uc2rb_desc_9_axuser_14_reg(uc2rb_desc_9_axuser_14_reg),
                                               .uc2rb_desc_9_axuser_15_reg(uc2rb_desc_9_axuser_15_reg),
                                               .uc2rb_desc_9_wuser_0_reg(uc2rb_desc_9_wuser_0_reg),
                                               .uc2rb_desc_9_wuser_1_reg(uc2rb_desc_9_wuser_1_reg),
                                               .uc2rb_desc_9_wuser_2_reg(uc2rb_desc_9_wuser_2_reg),
                                               .uc2rb_desc_9_wuser_3_reg(uc2rb_desc_9_wuser_3_reg),
                                               .uc2rb_desc_9_wuser_4_reg(uc2rb_desc_9_wuser_4_reg),
                                               .uc2rb_desc_9_wuser_5_reg(uc2rb_desc_9_wuser_5_reg),
                                               .uc2rb_desc_9_wuser_6_reg(uc2rb_desc_9_wuser_6_reg),
                                               .uc2rb_desc_9_wuser_7_reg(uc2rb_desc_9_wuser_7_reg),
                                               .uc2rb_desc_9_wuser_8_reg(uc2rb_desc_9_wuser_8_reg),
                                               .uc2rb_desc_9_wuser_9_reg(uc2rb_desc_9_wuser_9_reg),
                                               .uc2rb_desc_9_wuser_10_reg(uc2rb_desc_9_wuser_10_reg),
                                               .uc2rb_desc_9_wuser_11_reg(uc2rb_desc_9_wuser_11_reg),
                                               .uc2rb_desc_9_wuser_12_reg(uc2rb_desc_9_wuser_12_reg),
                                               .uc2rb_desc_9_wuser_13_reg(uc2rb_desc_9_wuser_13_reg),
                                               .uc2rb_desc_9_wuser_14_reg(uc2rb_desc_9_wuser_14_reg),
                                               .uc2rb_desc_9_wuser_15_reg(uc2rb_desc_9_wuser_15_reg),
                                               .uc2rb_desc_10_txn_type_reg(uc2rb_desc_10_txn_type_reg),
                                               .uc2rb_desc_10_size_reg(uc2rb_desc_10_size_reg),
                                               .uc2rb_desc_10_data_offset_reg(uc2rb_desc_10_data_offset_reg),
                                               .uc2rb_desc_10_axsize_reg(uc2rb_desc_10_axsize_reg),
                                               .uc2rb_desc_10_attr_reg(uc2rb_desc_10_attr_reg),
                                               .uc2rb_desc_10_axaddr_0_reg(uc2rb_desc_10_axaddr_0_reg),
                                               .uc2rb_desc_10_axaddr_1_reg(uc2rb_desc_10_axaddr_1_reg),
                                               .uc2rb_desc_10_axaddr_2_reg(uc2rb_desc_10_axaddr_2_reg),
                                               .uc2rb_desc_10_axaddr_3_reg(uc2rb_desc_10_axaddr_3_reg),
                                               .uc2rb_desc_10_axid_0_reg(uc2rb_desc_10_axid_0_reg),
                                               .uc2rb_desc_10_axid_1_reg(uc2rb_desc_10_axid_1_reg),
                                               .uc2rb_desc_10_axid_2_reg(uc2rb_desc_10_axid_2_reg),
                                               .uc2rb_desc_10_axid_3_reg(uc2rb_desc_10_axid_3_reg),
                                               .uc2rb_desc_10_axuser_0_reg(uc2rb_desc_10_axuser_0_reg),
                                               .uc2rb_desc_10_axuser_1_reg(uc2rb_desc_10_axuser_1_reg),
                                               .uc2rb_desc_10_axuser_2_reg(uc2rb_desc_10_axuser_2_reg),
                                               .uc2rb_desc_10_axuser_3_reg(uc2rb_desc_10_axuser_3_reg),
                                               .uc2rb_desc_10_axuser_4_reg(uc2rb_desc_10_axuser_4_reg),
                                               .uc2rb_desc_10_axuser_5_reg(uc2rb_desc_10_axuser_5_reg),
                                               .uc2rb_desc_10_axuser_6_reg(uc2rb_desc_10_axuser_6_reg),
                                               .uc2rb_desc_10_axuser_7_reg(uc2rb_desc_10_axuser_7_reg),
                                               .uc2rb_desc_10_axuser_8_reg(uc2rb_desc_10_axuser_8_reg),
                                               .uc2rb_desc_10_axuser_9_reg(uc2rb_desc_10_axuser_9_reg),
                                               .uc2rb_desc_10_axuser_10_reg(uc2rb_desc_10_axuser_10_reg),
                                               .uc2rb_desc_10_axuser_11_reg(uc2rb_desc_10_axuser_11_reg),
                                               .uc2rb_desc_10_axuser_12_reg(uc2rb_desc_10_axuser_12_reg),
                                               .uc2rb_desc_10_axuser_13_reg(uc2rb_desc_10_axuser_13_reg),
                                               .uc2rb_desc_10_axuser_14_reg(uc2rb_desc_10_axuser_14_reg),
                                               .uc2rb_desc_10_axuser_15_reg(uc2rb_desc_10_axuser_15_reg),
                                               .uc2rb_desc_10_wuser_0_reg(uc2rb_desc_10_wuser_0_reg),
                                               .uc2rb_desc_10_wuser_1_reg(uc2rb_desc_10_wuser_1_reg),
                                               .uc2rb_desc_10_wuser_2_reg(uc2rb_desc_10_wuser_2_reg),
                                               .uc2rb_desc_10_wuser_3_reg(uc2rb_desc_10_wuser_3_reg),
                                               .uc2rb_desc_10_wuser_4_reg(uc2rb_desc_10_wuser_4_reg),
                                               .uc2rb_desc_10_wuser_5_reg(uc2rb_desc_10_wuser_5_reg),
                                               .uc2rb_desc_10_wuser_6_reg(uc2rb_desc_10_wuser_6_reg),
                                               .uc2rb_desc_10_wuser_7_reg(uc2rb_desc_10_wuser_7_reg),
                                               .uc2rb_desc_10_wuser_8_reg(uc2rb_desc_10_wuser_8_reg),
                                               .uc2rb_desc_10_wuser_9_reg(uc2rb_desc_10_wuser_9_reg),
                                               .uc2rb_desc_10_wuser_10_reg(uc2rb_desc_10_wuser_10_reg),
                                               .uc2rb_desc_10_wuser_11_reg(uc2rb_desc_10_wuser_11_reg),
                                               .uc2rb_desc_10_wuser_12_reg(uc2rb_desc_10_wuser_12_reg),
                                               .uc2rb_desc_10_wuser_13_reg(uc2rb_desc_10_wuser_13_reg),
                                               .uc2rb_desc_10_wuser_14_reg(uc2rb_desc_10_wuser_14_reg),
                                               .uc2rb_desc_10_wuser_15_reg(uc2rb_desc_10_wuser_15_reg),
                                               .uc2rb_desc_11_txn_type_reg(uc2rb_desc_11_txn_type_reg),
                                               .uc2rb_desc_11_size_reg(uc2rb_desc_11_size_reg),
                                               .uc2rb_desc_11_data_offset_reg(uc2rb_desc_11_data_offset_reg),
                                               .uc2rb_desc_11_axsize_reg(uc2rb_desc_11_axsize_reg),
                                               .uc2rb_desc_11_attr_reg(uc2rb_desc_11_attr_reg),
                                               .uc2rb_desc_11_axaddr_0_reg(uc2rb_desc_11_axaddr_0_reg),
                                               .uc2rb_desc_11_axaddr_1_reg(uc2rb_desc_11_axaddr_1_reg),
                                               .uc2rb_desc_11_axaddr_2_reg(uc2rb_desc_11_axaddr_2_reg),
                                               .uc2rb_desc_11_axaddr_3_reg(uc2rb_desc_11_axaddr_3_reg),
                                               .uc2rb_desc_11_axid_0_reg(uc2rb_desc_11_axid_0_reg),
                                               .uc2rb_desc_11_axid_1_reg(uc2rb_desc_11_axid_1_reg),
                                               .uc2rb_desc_11_axid_2_reg(uc2rb_desc_11_axid_2_reg),
                                               .uc2rb_desc_11_axid_3_reg(uc2rb_desc_11_axid_3_reg),
                                               .uc2rb_desc_11_axuser_0_reg(uc2rb_desc_11_axuser_0_reg),
                                               .uc2rb_desc_11_axuser_1_reg(uc2rb_desc_11_axuser_1_reg),
                                               .uc2rb_desc_11_axuser_2_reg(uc2rb_desc_11_axuser_2_reg),
                                               .uc2rb_desc_11_axuser_3_reg(uc2rb_desc_11_axuser_3_reg),
                                               .uc2rb_desc_11_axuser_4_reg(uc2rb_desc_11_axuser_4_reg),
                                               .uc2rb_desc_11_axuser_5_reg(uc2rb_desc_11_axuser_5_reg),
                                               .uc2rb_desc_11_axuser_6_reg(uc2rb_desc_11_axuser_6_reg),
                                               .uc2rb_desc_11_axuser_7_reg(uc2rb_desc_11_axuser_7_reg),
                                               .uc2rb_desc_11_axuser_8_reg(uc2rb_desc_11_axuser_8_reg),
                                               .uc2rb_desc_11_axuser_9_reg(uc2rb_desc_11_axuser_9_reg),
                                               .uc2rb_desc_11_axuser_10_reg(uc2rb_desc_11_axuser_10_reg),
                                               .uc2rb_desc_11_axuser_11_reg(uc2rb_desc_11_axuser_11_reg),
                                               .uc2rb_desc_11_axuser_12_reg(uc2rb_desc_11_axuser_12_reg),
                                               .uc2rb_desc_11_axuser_13_reg(uc2rb_desc_11_axuser_13_reg),
                                               .uc2rb_desc_11_axuser_14_reg(uc2rb_desc_11_axuser_14_reg),
                                               .uc2rb_desc_11_axuser_15_reg(uc2rb_desc_11_axuser_15_reg),
                                               .uc2rb_desc_11_wuser_0_reg(uc2rb_desc_11_wuser_0_reg),
                                               .uc2rb_desc_11_wuser_1_reg(uc2rb_desc_11_wuser_1_reg),
                                               .uc2rb_desc_11_wuser_2_reg(uc2rb_desc_11_wuser_2_reg),
                                               .uc2rb_desc_11_wuser_3_reg(uc2rb_desc_11_wuser_3_reg),
                                               .uc2rb_desc_11_wuser_4_reg(uc2rb_desc_11_wuser_4_reg),
                                               .uc2rb_desc_11_wuser_5_reg(uc2rb_desc_11_wuser_5_reg),
                                               .uc2rb_desc_11_wuser_6_reg(uc2rb_desc_11_wuser_6_reg),
                                               .uc2rb_desc_11_wuser_7_reg(uc2rb_desc_11_wuser_7_reg),
                                               .uc2rb_desc_11_wuser_8_reg(uc2rb_desc_11_wuser_8_reg),
                                               .uc2rb_desc_11_wuser_9_reg(uc2rb_desc_11_wuser_9_reg),
                                               .uc2rb_desc_11_wuser_10_reg(uc2rb_desc_11_wuser_10_reg),
                                               .uc2rb_desc_11_wuser_11_reg(uc2rb_desc_11_wuser_11_reg),
                                               .uc2rb_desc_11_wuser_12_reg(uc2rb_desc_11_wuser_12_reg),
                                               .uc2rb_desc_11_wuser_13_reg(uc2rb_desc_11_wuser_13_reg),
                                               .uc2rb_desc_11_wuser_14_reg(uc2rb_desc_11_wuser_14_reg),
                                               .uc2rb_desc_11_wuser_15_reg(uc2rb_desc_11_wuser_15_reg),
                                               .uc2rb_desc_12_txn_type_reg(uc2rb_desc_12_txn_type_reg),
                                               .uc2rb_desc_12_size_reg(uc2rb_desc_12_size_reg),
                                               .uc2rb_desc_12_data_offset_reg(uc2rb_desc_12_data_offset_reg),
                                               .uc2rb_desc_12_axsize_reg(uc2rb_desc_12_axsize_reg),
                                               .uc2rb_desc_12_attr_reg(uc2rb_desc_12_attr_reg),
                                               .uc2rb_desc_12_axaddr_0_reg(uc2rb_desc_12_axaddr_0_reg),
                                               .uc2rb_desc_12_axaddr_1_reg(uc2rb_desc_12_axaddr_1_reg),
                                               .uc2rb_desc_12_axaddr_2_reg(uc2rb_desc_12_axaddr_2_reg),
                                               .uc2rb_desc_12_axaddr_3_reg(uc2rb_desc_12_axaddr_3_reg),
                                               .uc2rb_desc_12_axid_0_reg(uc2rb_desc_12_axid_0_reg),
                                               .uc2rb_desc_12_axid_1_reg(uc2rb_desc_12_axid_1_reg),
                                               .uc2rb_desc_12_axid_2_reg(uc2rb_desc_12_axid_2_reg),
                                               .uc2rb_desc_12_axid_3_reg(uc2rb_desc_12_axid_3_reg),
                                               .uc2rb_desc_12_axuser_0_reg(uc2rb_desc_12_axuser_0_reg),
                                               .uc2rb_desc_12_axuser_1_reg(uc2rb_desc_12_axuser_1_reg),
                                               .uc2rb_desc_12_axuser_2_reg(uc2rb_desc_12_axuser_2_reg),
                                               .uc2rb_desc_12_axuser_3_reg(uc2rb_desc_12_axuser_3_reg),
                                               .uc2rb_desc_12_axuser_4_reg(uc2rb_desc_12_axuser_4_reg),
                                               .uc2rb_desc_12_axuser_5_reg(uc2rb_desc_12_axuser_5_reg),
                                               .uc2rb_desc_12_axuser_6_reg(uc2rb_desc_12_axuser_6_reg),
                                               .uc2rb_desc_12_axuser_7_reg(uc2rb_desc_12_axuser_7_reg),
                                               .uc2rb_desc_12_axuser_8_reg(uc2rb_desc_12_axuser_8_reg),
                                               .uc2rb_desc_12_axuser_9_reg(uc2rb_desc_12_axuser_9_reg),
                                               .uc2rb_desc_12_axuser_10_reg(uc2rb_desc_12_axuser_10_reg),
                                               .uc2rb_desc_12_axuser_11_reg(uc2rb_desc_12_axuser_11_reg),
                                               .uc2rb_desc_12_axuser_12_reg(uc2rb_desc_12_axuser_12_reg),
                                               .uc2rb_desc_12_axuser_13_reg(uc2rb_desc_12_axuser_13_reg),
                                               .uc2rb_desc_12_axuser_14_reg(uc2rb_desc_12_axuser_14_reg),
                                               .uc2rb_desc_12_axuser_15_reg(uc2rb_desc_12_axuser_15_reg),
                                               .uc2rb_desc_12_wuser_0_reg(uc2rb_desc_12_wuser_0_reg),
                                               .uc2rb_desc_12_wuser_1_reg(uc2rb_desc_12_wuser_1_reg),
                                               .uc2rb_desc_12_wuser_2_reg(uc2rb_desc_12_wuser_2_reg),
                                               .uc2rb_desc_12_wuser_3_reg(uc2rb_desc_12_wuser_3_reg),
                                               .uc2rb_desc_12_wuser_4_reg(uc2rb_desc_12_wuser_4_reg),
                                               .uc2rb_desc_12_wuser_5_reg(uc2rb_desc_12_wuser_5_reg),
                                               .uc2rb_desc_12_wuser_6_reg(uc2rb_desc_12_wuser_6_reg),
                                               .uc2rb_desc_12_wuser_7_reg(uc2rb_desc_12_wuser_7_reg),
                                               .uc2rb_desc_12_wuser_8_reg(uc2rb_desc_12_wuser_8_reg),
                                               .uc2rb_desc_12_wuser_9_reg(uc2rb_desc_12_wuser_9_reg),
                                               .uc2rb_desc_12_wuser_10_reg(uc2rb_desc_12_wuser_10_reg),
                                               .uc2rb_desc_12_wuser_11_reg(uc2rb_desc_12_wuser_11_reg),
                                               .uc2rb_desc_12_wuser_12_reg(uc2rb_desc_12_wuser_12_reg),
                                               .uc2rb_desc_12_wuser_13_reg(uc2rb_desc_12_wuser_13_reg),
                                               .uc2rb_desc_12_wuser_14_reg(uc2rb_desc_12_wuser_14_reg),
                                               .uc2rb_desc_12_wuser_15_reg(uc2rb_desc_12_wuser_15_reg),
                                               .uc2rb_desc_13_txn_type_reg(uc2rb_desc_13_txn_type_reg),
                                               .uc2rb_desc_13_size_reg(uc2rb_desc_13_size_reg),
                                               .uc2rb_desc_13_data_offset_reg(uc2rb_desc_13_data_offset_reg),
                                               .uc2rb_desc_13_axsize_reg(uc2rb_desc_13_axsize_reg),
                                               .uc2rb_desc_13_attr_reg(uc2rb_desc_13_attr_reg),
                                               .uc2rb_desc_13_axaddr_0_reg(uc2rb_desc_13_axaddr_0_reg),
                                               .uc2rb_desc_13_axaddr_1_reg(uc2rb_desc_13_axaddr_1_reg),
                                               .uc2rb_desc_13_axaddr_2_reg(uc2rb_desc_13_axaddr_2_reg),
                                               .uc2rb_desc_13_axaddr_3_reg(uc2rb_desc_13_axaddr_3_reg),
                                               .uc2rb_desc_13_axid_0_reg(uc2rb_desc_13_axid_0_reg),
                                               .uc2rb_desc_13_axid_1_reg(uc2rb_desc_13_axid_1_reg),
                                               .uc2rb_desc_13_axid_2_reg(uc2rb_desc_13_axid_2_reg),
                                               .uc2rb_desc_13_axid_3_reg(uc2rb_desc_13_axid_3_reg),
                                               .uc2rb_desc_13_axuser_0_reg(uc2rb_desc_13_axuser_0_reg),
                                               .uc2rb_desc_13_axuser_1_reg(uc2rb_desc_13_axuser_1_reg),
                                               .uc2rb_desc_13_axuser_2_reg(uc2rb_desc_13_axuser_2_reg),
                                               .uc2rb_desc_13_axuser_3_reg(uc2rb_desc_13_axuser_3_reg),
                                               .uc2rb_desc_13_axuser_4_reg(uc2rb_desc_13_axuser_4_reg),
                                               .uc2rb_desc_13_axuser_5_reg(uc2rb_desc_13_axuser_5_reg),
                                               .uc2rb_desc_13_axuser_6_reg(uc2rb_desc_13_axuser_6_reg),
                                               .uc2rb_desc_13_axuser_7_reg(uc2rb_desc_13_axuser_7_reg),
                                               .uc2rb_desc_13_axuser_8_reg(uc2rb_desc_13_axuser_8_reg),
                                               .uc2rb_desc_13_axuser_9_reg(uc2rb_desc_13_axuser_9_reg),
                                               .uc2rb_desc_13_axuser_10_reg(uc2rb_desc_13_axuser_10_reg),
                                               .uc2rb_desc_13_axuser_11_reg(uc2rb_desc_13_axuser_11_reg),
                                               .uc2rb_desc_13_axuser_12_reg(uc2rb_desc_13_axuser_12_reg),
                                               .uc2rb_desc_13_axuser_13_reg(uc2rb_desc_13_axuser_13_reg),
                                               .uc2rb_desc_13_axuser_14_reg(uc2rb_desc_13_axuser_14_reg),
                                               .uc2rb_desc_13_axuser_15_reg(uc2rb_desc_13_axuser_15_reg),
                                               .uc2rb_desc_13_wuser_0_reg(uc2rb_desc_13_wuser_0_reg),
                                               .uc2rb_desc_13_wuser_1_reg(uc2rb_desc_13_wuser_1_reg),
                                               .uc2rb_desc_13_wuser_2_reg(uc2rb_desc_13_wuser_2_reg),
                                               .uc2rb_desc_13_wuser_3_reg(uc2rb_desc_13_wuser_3_reg),
                                               .uc2rb_desc_13_wuser_4_reg(uc2rb_desc_13_wuser_4_reg),
                                               .uc2rb_desc_13_wuser_5_reg(uc2rb_desc_13_wuser_5_reg),
                                               .uc2rb_desc_13_wuser_6_reg(uc2rb_desc_13_wuser_6_reg),
                                               .uc2rb_desc_13_wuser_7_reg(uc2rb_desc_13_wuser_7_reg),
                                               .uc2rb_desc_13_wuser_8_reg(uc2rb_desc_13_wuser_8_reg),
                                               .uc2rb_desc_13_wuser_9_reg(uc2rb_desc_13_wuser_9_reg),
                                               .uc2rb_desc_13_wuser_10_reg(uc2rb_desc_13_wuser_10_reg),
                                               .uc2rb_desc_13_wuser_11_reg(uc2rb_desc_13_wuser_11_reg),
                                               .uc2rb_desc_13_wuser_12_reg(uc2rb_desc_13_wuser_12_reg),
                                               .uc2rb_desc_13_wuser_13_reg(uc2rb_desc_13_wuser_13_reg),
                                               .uc2rb_desc_13_wuser_14_reg(uc2rb_desc_13_wuser_14_reg),
                                               .uc2rb_desc_13_wuser_15_reg(uc2rb_desc_13_wuser_15_reg),
                                               .uc2rb_desc_14_txn_type_reg(uc2rb_desc_14_txn_type_reg),
                                               .uc2rb_desc_14_size_reg(uc2rb_desc_14_size_reg),
                                               .uc2rb_desc_14_data_offset_reg(uc2rb_desc_14_data_offset_reg),
                                               .uc2rb_desc_14_axsize_reg(uc2rb_desc_14_axsize_reg),
                                               .uc2rb_desc_14_attr_reg(uc2rb_desc_14_attr_reg),
                                               .uc2rb_desc_14_axaddr_0_reg(uc2rb_desc_14_axaddr_0_reg),
                                               .uc2rb_desc_14_axaddr_1_reg(uc2rb_desc_14_axaddr_1_reg),
                                               .uc2rb_desc_14_axaddr_2_reg(uc2rb_desc_14_axaddr_2_reg),
                                               .uc2rb_desc_14_axaddr_3_reg(uc2rb_desc_14_axaddr_3_reg),
                                               .uc2rb_desc_14_axid_0_reg(uc2rb_desc_14_axid_0_reg),
                                               .uc2rb_desc_14_axid_1_reg(uc2rb_desc_14_axid_1_reg),
                                               .uc2rb_desc_14_axid_2_reg(uc2rb_desc_14_axid_2_reg),
                                               .uc2rb_desc_14_axid_3_reg(uc2rb_desc_14_axid_3_reg),
                                               .uc2rb_desc_14_axuser_0_reg(uc2rb_desc_14_axuser_0_reg),
                                               .uc2rb_desc_14_axuser_1_reg(uc2rb_desc_14_axuser_1_reg),
                                               .uc2rb_desc_14_axuser_2_reg(uc2rb_desc_14_axuser_2_reg),
                                               .uc2rb_desc_14_axuser_3_reg(uc2rb_desc_14_axuser_3_reg),
                                               .uc2rb_desc_14_axuser_4_reg(uc2rb_desc_14_axuser_4_reg),
                                               .uc2rb_desc_14_axuser_5_reg(uc2rb_desc_14_axuser_5_reg),
                                               .uc2rb_desc_14_axuser_6_reg(uc2rb_desc_14_axuser_6_reg),
                                               .uc2rb_desc_14_axuser_7_reg(uc2rb_desc_14_axuser_7_reg),
                                               .uc2rb_desc_14_axuser_8_reg(uc2rb_desc_14_axuser_8_reg),
                                               .uc2rb_desc_14_axuser_9_reg(uc2rb_desc_14_axuser_9_reg),
                                               .uc2rb_desc_14_axuser_10_reg(uc2rb_desc_14_axuser_10_reg),
                                               .uc2rb_desc_14_axuser_11_reg(uc2rb_desc_14_axuser_11_reg),
                                               .uc2rb_desc_14_axuser_12_reg(uc2rb_desc_14_axuser_12_reg),
                                               .uc2rb_desc_14_axuser_13_reg(uc2rb_desc_14_axuser_13_reg),
                                               .uc2rb_desc_14_axuser_14_reg(uc2rb_desc_14_axuser_14_reg),
                                               .uc2rb_desc_14_axuser_15_reg(uc2rb_desc_14_axuser_15_reg),
                                               .uc2rb_desc_14_wuser_0_reg(uc2rb_desc_14_wuser_0_reg),
                                               .uc2rb_desc_14_wuser_1_reg(uc2rb_desc_14_wuser_1_reg),
                                               .uc2rb_desc_14_wuser_2_reg(uc2rb_desc_14_wuser_2_reg),
                                               .uc2rb_desc_14_wuser_3_reg(uc2rb_desc_14_wuser_3_reg),
                                               .uc2rb_desc_14_wuser_4_reg(uc2rb_desc_14_wuser_4_reg),
                                               .uc2rb_desc_14_wuser_5_reg(uc2rb_desc_14_wuser_5_reg),
                                               .uc2rb_desc_14_wuser_6_reg(uc2rb_desc_14_wuser_6_reg),
                                               .uc2rb_desc_14_wuser_7_reg(uc2rb_desc_14_wuser_7_reg),
                                               .uc2rb_desc_14_wuser_8_reg(uc2rb_desc_14_wuser_8_reg),
                                               .uc2rb_desc_14_wuser_9_reg(uc2rb_desc_14_wuser_9_reg),
                                               .uc2rb_desc_14_wuser_10_reg(uc2rb_desc_14_wuser_10_reg),
                                               .uc2rb_desc_14_wuser_11_reg(uc2rb_desc_14_wuser_11_reg),
                                               .uc2rb_desc_14_wuser_12_reg(uc2rb_desc_14_wuser_12_reg),
                                               .uc2rb_desc_14_wuser_13_reg(uc2rb_desc_14_wuser_13_reg),
                                               .uc2rb_desc_14_wuser_14_reg(uc2rb_desc_14_wuser_14_reg),
                                               .uc2rb_desc_14_wuser_15_reg(uc2rb_desc_14_wuser_15_reg),
                                               .uc2rb_desc_15_txn_type_reg(uc2rb_desc_15_txn_type_reg),
                                               .uc2rb_desc_15_size_reg(uc2rb_desc_15_size_reg),
                                               .uc2rb_desc_15_data_offset_reg(uc2rb_desc_15_data_offset_reg),
                                               .uc2rb_desc_15_axsize_reg(uc2rb_desc_15_axsize_reg),
                                               .uc2rb_desc_15_attr_reg(uc2rb_desc_15_attr_reg),
                                               .uc2rb_desc_15_axaddr_0_reg(uc2rb_desc_15_axaddr_0_reg),
                                               .uc2rb_desc_15_axaddr_1_reg(uc2rb_desc_15_axaddr_1_reg),
                                               .uc2rb_desc_15_axaddr_2_reg(uc2rb_desc_15_axaddr_2_reg),
                                               .uc2rb_desc_15_axaddr_3_reg(uc2rb_desc_15_axaddr_3_reg),
                                               .uc2rb_desc_15_axid_0_reg(uc2rb_desc_15_axid_0_reg),
                                               .uc2rb_desc_15_axid_1_reg(uc2rb_desc_15_axid_1_reg),
                                               .uc2rb_desc_15_axid_2_reg(uc2rb_desc_15_axid_2_reg),
                                               .uc2rb_desc_15_axid_3_reg(uc2rb_desc_15_axid_3_reg),
                                               .uc2rb_desc_15_axuser_0_reg(uc2rb_desc_15_axuser_0_reg),
                                               .uc2rb_desc_15_axuser_1_reg(uc2rb_desc_15_axuser_1_reg),
                                               .uc2rb_desc_15_axuser_2_reg(uc2rb_desc_15_axuser_2_reg),
                                               .uc2rb_desc_15_axuser_3_reg(uc2rb_desc_15_axuser_3_reg),
                                               .uc2rb_desc_15_axuser_4_reg(uc2rb_desc_15_axuser_4_reg),
                                               .uc2rb_desc_15_axuser_5_reg(uc2rb_desc_15_axuser_5_reg),
                                               .uc2rb_desc_15_axuser_6_reg(uc2rb_desc_15_axuser_6_reg),
                                               .uc2rb_desc_15_axuser_7_reg(uc2rb_desc_15_axuser_7_reg),
                                               .uc2rb_desc_15_axuser_8_reg(uc2rb_desc_15_axuser_8_reg),
                                               .uc2rb_desc_15_axuser_9_reg(uc2rb_desc_15_axuser_9_reg),
                                               .uc2rb_desc_15_axuser_10_reg(uc2rb_desc_15_axuser_10_reg),
                                               .uc2rb_desc_15_axuser_11_reg(uc2rb_desc_15_axuser_11_reg),
                                               .uc2rb_desc_15_axuser_12_reg(uc2rb_desc_15_axuser_12_reg),
                                               .uc2rb_desc_15_axuser_13_reg(uc2rb_desc_15_axuser_13_reg),
                                               .uc2rb_desc_15_axuser_14_reg(uc2rb_desc_15_axuser_14_reg),
                                               .uc2rb_desc_15_axuser_15_reg(uc2rb_desc_15_axuser_15_reg),
                                               .uc2rb_desc_15_wuser_0_reg(uc2rb_desc_15_wuser_0_reg),
                                               .uc2rb_desc_15_wuser_1_reg(uc2rb_desc_15_wuser_1_reg),
                                               .uc2rb_desc_15_wuser_2_reg(uc2rb_desc_15_wuser_2_reg),
                                               .uc2rb_desc_15_wuser_3_reg(uc2rb_desc_15_wuser_3_reg),
                                               .uc2rb_desc_15_wuser_4_reg(uc2rb_desc_15_wuser_4_reg),
                                               .uc2rb_desc_15_wuser_5_reg(uc2rb_desc_15_wuser_5_reg),
                                               .uc2rb_desc_15_wuser_6_reg(uc2rb_desc_15_wuser_6_reg),
                                               .uc2rb_desc_15_wuser_7_reg(uc2rb_desc_15_wuser_7_reg),
                                               .uc2rb_desc_15_wuser_8_reg(uc2rb_desc_15_wuser_8_reg),
                                               .uc2rb_desc_15_wuser_9_reg(uc2rb_desc_15_wuser_9_reg),
                                               .uc2rb_desc_15_wuser_10_reg(uc2rb_desc_15_wuser_10_reg),
                                               .uc2rb_desc_15_wuser_11_reg(uc2rb_desc_15_wuser_11_reg),
                                               .uc2rb_desc_15_wuser_12_reg(uc2rb_desc_15_wuser_12_reg),
                                               .uc2rb_desc_15_wuser_13_reg(uc2rb_desc_15_wuser_13_reg),
                                               .uc2rb_desc_15_wuser_14_reg(uc2rb_desc_15_wuser_14_reg),
                                               .uc2rb_desc_15_wuser_15_reg(uc2rb_desc_15_wuser_15_reg),
                                               .uc2rb_intr_error_status_reg_we(uc2rb_intr_error_status_reg_we),
                                               .uc2rb_ownership_reg_we(uc2rb_ownership_reg_we),
                                               .uc2rb_intr_txn_avail_status_reg_we(uc2rb_intr_txn_avail_status_reg_we),
                                               .uc2rb_intr_comp_status_reg_we(uc2rb_intr_comp_status_reg_we),
                                               .uc2rb_status_busy_reg_we(uc2rb_status_busy_reg_we),
                                               .uc2rb_resp_fifo_free_level_reg_we(uc2rb_resp_fifo_free_level_reg_we),
                                               .uc2rb_desc_0_txn_type_reg_we(uc2rb_desc_0_txn_type_reg_we),
                                               .uc2rb_desc_0_size_reg_we(uc2rb_desc_0_size_reg_we),
                                               .uc2rb_desc_0_data_offset_reg_we(uc2rb_desc_0_data_offset_reg_we),
                                               .uc2rb_desc_0_axsize_reg_we(uc2rb_desc_0_axsize_reg_we),
                                               .uc2rb_desc_0_attr_reg_we(uc2rb_desc_0_attr_reg_we),
                                               .uc2rb_desc_0_axaddr_0_reg_we(uc2rb_desc_0_axaddr_0_reg_we),
                                               .uc2rb_desc_0_axaddr_1_reg_we(uc2rb_desc_0_axaddr_1_reg_we),
                                               .uc2rb_desc_0_axaddr_2_reg_we(uc2rb_desc_0_axaddr_2_reg_we),
                                               .uc2rb_desc_0_axaddr_3_reg_we(uc2rb_desc_0_axaddr_3_reg_we),
                                               .uc2rb_desc_0_axid_0_reg_we(uc2rb_desc_0_axid_0_reg_we),
                                               .uc2rb_desc_0_axid_1_reg_we(uc2rb_desc_0_axid_1_reg_we),
                                               .uc2rb_desc_0_axid_2_reg_we(uc2rb_desc_0_axid_2_reg_we),
                                               .uc2rb_desc_0_axid_3_reg_we(uc2rb_desc_0_axid_3_reg_we),
                                               .uc2rb_desc_0_axuser_0_reg_we(uc2rb_desc_0_axuser_0_reg_we),
                                               .uc2rb_desc_0_axuser_1_reg_we(uc2rb_desc_0_axuser_1_reg_we),
                                               .uc2rb_desc_0_axuser_2_reg_we(uc2rb_desc_0_axuser_2_reg_we),
                                               .uc2rb_desc_0_axuser_3_reg_we(uc2rb_desc_0_axuser_3_reg_we),
                                               .uc2rb_desc_0_axuser_4_reg_we(uc2rb_desc_0_axuser_4_reg_we),
                                               .uc2rb_desc_0_axuser_5_reg_we(uc2rb_desc_0_axuser_5_reg_we),
                                               .uc2rb_desc_0_axuser_6_reg_we(uc2rb_desc_0_axuser_6_reg_we),
                                               .uc2rb_desc_0_axuser_7_reg_we(uc2rb_desc_0_axuser_7_reg_we),
                                               .uc2rb_desc_0_axuser_8_reg_we(uc2rb_desc_0_axuser_8_reg_we),
                                               .uc2rb_desc_0_axuser_9_reg_we(uc2rb_desc_0_axuser_9_reg_we),
                                               .uc2rb_desc_0_axuser_10_reg_we(uc2rb_desc_0_axuser_10_reg_we),
                                               .uc2rb_desc_0_axuser_11_reg_we(uc2rb_desc_0_axuser_11_reg_we),
                                               .uc2rb_desc_0_axuser_12_reg_we(uc2rb_desc_0_axuser_12_reg_we),
                                               .uc2rb_desc_0_axuser_13_reg_we(uc2rb_desc_0_axuser_13_reg_we),
                                               .uc2rb_desc_0_axuser_14_reg_we(uc2rb_desc_0_axuser_14_reg_we),
                                               .uc2rb_desc_0_axuser_15_reg_we(uc2rb_desc_0_axuser_15_reg_we),
                                               .uc2rb_desc_0_wuser_0_reg_we(uc2rb_desc_0_wuser_0_reg_we),
                                               .uc2rb_desc_0_wuser_1_reg_we(uc2rb_desc_0_wuser_1_reg_we),
                                               .uc2rb_desc_0_wuser_2_reg_we(uc2rb_desc_0_wuser_2_reg_we),
                                               .uc2rb_desc_0_wuser_3_reg_we(uc2rb_desc_0_wuser_3_reg_we),
                                               .uc2rb_desc_0_wuser_4_reg_we(uc2rb_desc_0_wuser_4_reg_we),
                                               .uc2rb_desc_0_wuser_5_reg_we(uc2rb_desc_0_wuser_5_reg_we),
                                               .uc2rb_desc_0_wuser_6_reg_we(uc2rb_desc_0_wuser_6_reg_we),
                                               .uc2rb_desc_0_wuser_7_reg_we(uc2rb_desc_0_wuser_7_reg_we),
                                               .uc2rb_desc_0_wuser_8_reg_we(uc2rb_desc_0_wuser_8_reg_we),
                                               .uc2rb_desc_0_wuser_9_reg_we(uc2rb_desc_0_wuser_9_reg_we),
                                               .uc2rb_desc_0_wuser_10_reg_we(uc2rb_desc_0_wuser_10_reg_we),
                                               .uc2rb_desc_0_wuser_11_reg_we(uc2rb_desc_0_wuser_11_reg_we),
                                               .uc2rb_desc_0_wuser_12_reg_we(uc2rb_desc_0_wuser_12_reg_we),
                                               .uc2rb_desc_0_wuser_13_reg_we(uc2rb_desc_0_wuser_13_reg_we),
                                               .uc2rb_desc_0_wuser_14_reg_we(uc2rb_desc_0_wuser_14_reg_we),
                                               .uc2rb_desc_0_wuser_15_reg_we(uc2rb_desc_0_wuser_15_reg_we),
                                               .uc2rb_desc_1_txn_type_reg_we(uc2rb_desc_1_txn_type_reg_we),
                                               .uc2rb_desc_1_size_reg_we(uc2rb_desc_1_size_reg_we),
                                               .uc2rb_desc_1_data_offset_reg_we(uc2rb_desc_1_data_offset_reg_we),
                                               .uc2rb_desc_1_axsize_reg_we(uc2rb_desc_1_axsize_reg_we),
                                               .uc2rb_desc_1_attr_reg_we(uc2rb_desc_1_attr_reg_we),
                                               .uc2rb_desc_1_axaddr_0_reg_we(uc2rb_desc_1_axaddr_0_reg_we),
                                               .uc2rb_desc_1_axaddr_1_reg_we(uc2rb_desc_1_axaddr_1_reg_we),
                                               .uc2rb_desc_1_axaddr_2_reg_we(uc2rb_desc_1_axaddr_2_reg_we),
                                               .uc2rb_desc_1_axaddr_3_reg_we(uc2rb_desc_1_axaddr_3_reg_we),
                                               .uc2rb_desc_1_axid_0_reg_we(uc2rb_desc_1_axid_0_reg_we),
                                               .uc2rb_desc_1_axid_1_reg_we(uc2rb_desc_1_axid_1_reg_we),
                                               .uc2rb_desc_1_axid_2_reg_we(uc2rb_desc_1_axid_2_reg_we),
                                               .uc2rb_desc_1_axid_3_reg_we(uc2rb_desc_1_axid_3_reg_we),
                                               .uc2rb_desc_1_axuser_0_reg_we(uc2rb_desc_1_axuser_0_reg_we),
                                               .uc2rb_desc_1_axuser_1_reg_we(uc2rb_desc_1_axuser_1_reg_we),
                                               .uc2rb_desc_1_axuser_2_reg_we(uc2rb_desc_1_axuser_2_reg_we),
                                               .uc2rb_desc_1_axuser_3_reg_we(uc2rb_desc_1_axuser_3_reg_we),
                                               .uc2rb_desc_1_axuser_4_reg_we(uc2rb_desc_1_axuser_4_reg_we),
                                               .uc2rb_desc_1_axuser_5_reg_we(uc2rb_desc_1_axuser_5_reg_we),
                                               .uc2rb_desc_1_axuser_6_reg_we(uc2rb_desc_1_axuser_6_reg_we),
                                               .uc2rb_desc_1_axuser_7_reg_we(uc2rb_desc_1_axuser_7_reg_we),
                                               .uc2rb_desc_1_axuser_8_reg_we(uc2rb_desc_1_axuser_8_reg_we),
                                               .uc2rb_desc_1_axuser_9_reg_we(uc2rb_desc_1_axuser_9_reg_we),
                                               .uc2rb_desc_1_axuser_10_reg_we(uc2rb_desc_1_axuser_10_reg_we),
                                               .uc2rb_desc_1_axuser_11_reg_we(uc2rb_desc_1_axuser_11_reg_we),
                                               .uc2rb_desc_1_axuser_12_reg_we(uc2rb_desc_1_axuser_12_reg_we),
                                               .uc2rb_desc_1_axuser_13_reg_we(uc2rb_desc_1_axuser_13_reg_we),
                                               .uc2rb_desc_1_axuser_14_reg_we(uc2rb_desc_1_axuser_14_reg_we),
                                               .uc2rb_desc_1_axuser_15_reg_we(uc2rb_desc_1_axuser_15_reg_we),
                                               .uc2rb_desc_1_wuser_0_reg_we(uc2rb_desc_1_wuser_0_reg_we),
                                               .uc2rb_desc_1_wuser_1_reg_we(uc2rb_desc_1_wuser_1_reg_we),
                                               .uc2rb_desc_1_wuser_2_reg_we(uc2rb_desc_1_wuser_2_reg_we),
                                               .uc2rb_desc_1_wuser_3_reg_we(uc2rb_desc_1_wuser_3_reg_we),
                                               .uc2rb_desc_1_wuser_4_reg_we(uc2rb_desc_1_wuser_4_reg_we),
                                               .uc2rb_desc_1_wuser_5_reg_we(uc2rb_desc_1_wuser_5_reg_we),
                                               .uc2rb_desc_1_wuser_6_reg_we(uc2rb_desc_1_wuser_6_reg_we),
                                               .uc2rb_desc_1_wuser_7_reg_we(uc2rb_desc_1_wuser_7_reg_we),
                                               .uc2rb_desc_1_wuser_8_reg_we(uc2rb_desc_1_wuser_8_reg_we),
                                               .uc2rb_desc_1_wuser_9_reg_we(uc2rb_desc_1_wuser_9_reg_we),
                                               .uc2rb_desc_1_wuser_10_reg_we(uc2rb_desc_1_wuser_10_reg_we),
                                               .uc2rb_desc_1_wuser_11_reg_we(uc2rb_desc_1_wuser_11_reg_we),
                                               .uc2rb_desc_1_wuser_12_reg_we(uc2rb_desc_1_wuser_12_reg_we),
                                               .uc2rb_desc_1_wuser_13_reg_we(uc2rb_desc_1_wuser_13_reg_we),
                                               .uc2rb_desc_1_wuser_14_reg_we(uc2rb_desc_1_wuser_14_reg_we),
                                               .uc2rb_desc_1_wuser_15_reg_we(uc2rb_desc_1_wuser_15_reg_we),
                                               .uc2rb_desc_2_txn_type_reg_we(uc2rb_desc_2_txn_type_reg_we),
                                               .uc2rb_desc_2_size_reg_we(uc2rb_desc_2_size_reg_we),
                                               .uc2rb_desc_2_data_offset_reg_we(uc2rb_desc_2_data_offset_reg_we),
                                               .uc2rb_desc_2_axsize_reg_we(uc2rb_desc_2_axsize_reg_we),
                                               .uc2rb_desc_2_attr_reg_we(uc2rb_desc_2_attr_reg_we),
                                               .uc2rb_desc_2_axaddr_0_reg_we(uc2rb_desc_2_axaddr_0_reg_we),
                                               .uc2rb_desc_2_axaddr_1_reg_we(uc2rb_desc_2_axaddr_1_reg_we),
                                               .uc2rb_desc_2_axaddr_2_reg_we(uc2rb_desc_2_axaddr_2_reg_we),
                                               .uc2rb_desc_2_axaddr_3_reg_we(uc2rb_desc_2_axaddr_3_reg_we),
                                               .uc2rb_desc_2_axid_0_reg_we(uc2rb_desc_2_axid_0_reg_we),
                                               .uc2rb_desc_2_axid_1_reg_we(uc2rb_desc_2_axid_1_reg_we),
                                               .uc2rb_desc_2_axid_2_reg_we(uc2rb_desc_2_axid_2_reg_we),
                                               .uc2rb_desc_2_axid_3_reg_we(uc2rb_desc_2_axid_3_reg_we),
                                               .uc2rb_desc_2_axuser_0_reg_we(uc2rb_desc_2_axuser_0_reg_we),
                                               .uc2rb_desc_2_axuser_1_reg_we(uc2rb_desc_2_axuser_1_reg_we),
                                               .uc2rb_desc_2_axuser_2_reg_we(uc2rb_desc_2_axuser_2_reg_we),
                                               .uc2rb_desc_2_axuser_3_reg_we(uc2rb_desc_2_axuser_3_reg_we),
                                               .uc2rb_desc_2_axuser_4_reg_we(uc2rb_desc_2_axuser_4_reg_we),
                                               .uc2rb_desc_2_axuser_5_reg_we(uc2rb_desc_2_axuser_5_reg_we),
                                               .uc2rb_desc_2_axuser_6_reg_we(uc2rb_desc_2_axuser_6_reg_we),
                                               .uc2rb_desc_2_axuser_7_reg_we(uc2rb_desc_2_axuser_7_reg_we),
                                               .uc2rb_desc_2_axuser_8_reg_we(uc2rb_desc_2_axuser_8_reg_we),
                                               .uc2rb_desc_2_axuser_9_reg_we(uc2rb_desc_2_axuser_9_reg_we),
                                               .uc2rb_desc_2_axuser_10_reg_we(uc2rb_desc_2_axuser_10_reg_we),
                                               .uc2rb_desc_2_axuser_11_reg_we(uc2rb_desc_2_axuser_11_reg_we),
                                               .uc2rb_desc_2_axuser_12_reg_we(uc2rb_desc_2_axuser_12_reg_we),
                                               .uc2rb_desc_2_axuser_13_reg_we(uc2rb_desc_2_axuser_13_reg_we),
                                               .uc2rb_desc_2_axuser_14_reg_we(uc2rb_desc_2_axuser_14_reg_we),
                                               .uc2rb_desc_2_axuser_15_reg_we(uc2rb_desc_2_axuser_15_reg_we),
                                               .uc2rb_desc_2_wuser_0_reg_we(uc2rb_desc_2_wuser_0_reg_we),
                                               .uc2rb_desc_2_wuser_1_reg_we(uc2rb_desc_2_wuser_1_reg_we),
                                               .uc2rb_desc_2_wuser_2_reg_we(uc2rb_desc_2_wuser_2_reg_we),
                                               .uc2rb_desc_2_wuser_3_reg_we(uc2rb_desc_2_wuser_3_reg_we),
                                               .uc2rb_desc_2_wuser_4_reg_we(uc2rb_desc_2_wuser_4_reg_we),
                                               .uc2rb_desc_2_wuser_5_reg_we(uc2rb_desc_2_wuser_5_reg_we),
                                               .uc2rb_desc_2_wuser_6_reg_we(uc2rb_desc_2_wuser_6_reg_we),
                                               .uc2rb_desc_2_wuser_7_reg_we(uc2rb_desc_2_wuser_7_reg_we),
                                               .uc2rb_desc_2_wuser_8_reg_we(uc2rb_desc_2_wuser_8_reg_we),
                                               .uc2rb_desc_2_wuser_9_reg_we(uc2rb_desc_2_wuser_9_reg_we),
                                               .uc2rb_desc_2_wuser_10_reg_we(uc2rb_desc_2_wuser_10_reg_we),
                                               .uc2rb_desc_2_wuser_11_reg_we(uc2rb_desc_2_wuser_11_reg_we),
                                               .uc2rb_desc_2_wuser_12_reg_we(uc2rb_desc_2_wuser_12_reg_we),
                                               .uc2rb_desc_2_wuser_13_reg_we(uc2rb_desc_2_wuser_13_reg_we),
                                               .uc2rb_desc_2_wuser_14_reg_we(uc2rb_desc_2_wuser_14_reg_we),
                                               .uc2rb_desc_2_wuser_15_reg_we(uc2rb_desc_2_wuser_15_reg_we),
                                               .uc2rb_desc_3_txn_type_reg_we(uc2rb_desc_3_txn_type_reg_we),
                                               .uc2rb_desc_3_size_reg_we(uc2rb_desc_3_size_reg_we),
                                               .uc2rb_desc_3_data_offset_reg_we(uc2rb_desc_3_data_offset_reg_we),
                                               .uc2rb_desc_3_axsize_reg_we(uc2rb_desc_3_axsize_reg_we),
                                               .uc2rb_desc_3_attr_reg_we(uc2rb_desc_3_attr_reg_we),
                                               .uc2rb_desc_3_axaddr_0_reg_we(uc2rb_desc_3_axaddr_0_reg_we),
                                               .uc2rb_desc_3_axaddr_1_reg_we(uc2rb_desc_3_axaddr_1_reg_we),
                                               .uc2rb_desc_3_axaddr_2_reg_we(uc2rb_desc_3_axaddr_2_reg_we),
                                               .uc2rb_desc_3_axaddr_3_reg_we(uc2rb_desc_3_axaddr_3_reg_we),
                                               .uc2rb_desc_3_axid_0_reg_we(uc2rb_desc_3_axid_0_reg_we),
                                               .uc2rb_desc_3_axid_1_reg_we(uc2rb_desc_3_axid_1_reg_we),
                                               .uc2rb_desc_3_axid_2_reg_we(uc2rb_desc_3_axid_2_reg_we),
                                               .uc2rb_desc_3_axid_3_reg_we(uc2rb_desc_3_axid_3_reg_we),
                                               .uc2rb_desc_3_axuser_0_reg_we(uc2rb_desc_3_axuser_0_reg_we),
                                               .uc2rb_desc_3_axuser_1_reg_we(uc2rb_desc_3_axuser_1_reg_we),
                                               .uc2rb_desc_3_axuser_2_reg_we(uc2rb_desc_3_axuser_2_reg_we),
                                               .uc2rb_desc_3_axuser_3_reg_we(uc2rb_desc_3_axuser_3_reg_we),
                                               .uc2rb_desc_3_axuser_4_reg_we(uc2rb_desc_3_axuser_4_reg_we),
                                               .uc2rb_desc_3_axuser_5_reg_we(uc2rb_desc_3_axuser_5_reg_we),
                                               .uc2rb_desc_3_axuser_6_reg_we(uc2rb_desc_3_axuser_6_reg_we),
                                               .uc2rb_desc_3_axuser_7_reg_we(uc2rb_desc_3_axuser_7_reg_we),
                                               .uc2rb_desc_3_axuser_8_reg_we(uc2rb_desc_3_axuser_8_reg_we),
                                               .uc2rb_desc_3_axuser_9_reg_we(uc2rb_desc_3_axuser_9_reg_we),
                                               .uc2rb_desc_3_axuser_10_reg_we(uc2rb_desc_3_axuser_10_reg_we),
                                               .uc2rb_desc_3_axuser_11_reg_we(uc2rb_desc_3_axuser_11_reg_we),
                                               .uc2rb_desc_3_axuser_12_reg_we(uc2rb_desc_3_axuser_12_reg_we),
                                               .uc2rb_desc_3_axuser_13_reg_we(uc2rb_desc_3_axuser_13_reg_we),
                                               .uc2rb_desc_3_axuser_14_reg_we(uc2rb_desc_3_axuser_14_reg_we),
                                               .uc2rb_desc_3_axuser_15_reg_we(uc2rb_desc_3_axuser_15_reg_we),
                                               .uc2rb_desc_3_wuser_0_reg_we(uc2rb_desc_3_wuser_0_reg_we),
                                               .uc2rb_desc_3_wuser_1_reg_we(uc2rb_desc_3_wuser_1_reg_we),
                                               .uc2rb_desc_3_wuser_2_reg_we(uc2rb_desc_3_wuser_2_reg_we),
                                               .uc2rb_desc_3_wuser_3_reg_we(uc2rb_desc_3_wuser_3_reg_we),
                                               .uc2rb_desc_3_wuser_4_reg_we(uc2rb_desc_3_wuser_4_reg_we),
                                               .uc2rb_desc_3_wuser_5_reg_we(uc2rb_desc_3_wuser_5_reg_we),
                                               .uc2rb_desc_3_wuser_6_reg_we(uc2rb_desc_3_wuser_6_reg_we),
                                               .uc2rb_desc_3_wuser_7_reg_we(uc2rb_desc_3_wuser_7_reg_we),
                                               .uc2rb_desc_3_wuser_8_reg_we(uc2rb_desc_3_wuser_8_reg_we),
                                               .uc2rb_desc_3_wuser_9_reg_we(uc2rb_desc_3_wuser_9_reg_we),
                                               .uc2rb_desc_3_wuser_10_reg_we(uc2rb_desc_3_wuser_10_reg_we),
                                               .uc2rb_desc_3_wuser_11_reg_we(uc2rb_desc_3_wuser_11_reg_we),
                                               .uc2rb_desc_3_wuser_12_reg_we(uc2rb_desc_3_wuser_12_reg_we),
                                               .uc2rb_desc_3_wuser_13_reg_we(uc2rb_desc_3_wuser_13_reg_we),
                                               .uc2rb_desc_3_wuser_14_reg_we(uc2rb_desc_3_wuser_14_reg_we),
                                               .uc2rb_desc_3_wuser_15_reg_we(uc2rb_desc_3_wuser_15_reg_we),
                                               .uc2rb_desc_4_txn_type_reg_we(uc2rb_desc_4_txn_type_reg_we),
                                               .uc2rb_desc_4_size_reg_we(uc2rb_desc_4_size_reg_we),
                                               .uc2rb_desc_4_data_offset_reg_we(uc2rb_desc_4_data_offset_reg_we),
                                               .uc2rb_desc_4_axsize_reg_we(uc2rb_desc_4_axsize_reg_we),
                                               .uc2rb_desc_4_attr_reg_we(uc2rb_desc_4_attr_reg_we),
                                               .uc2rb_desc_4_axaddr_0_reg_we(uc2rb_desc_4_axaddr_0_reg_we),
                                               .uc2rb_desc_4_axaddr_1_reg_we(uc2rb_desc_4_axaddr_1_reg_we),
                                               .uc2rb_desc_4_axaddr_2_reg_we(uc2rb_desc_4_axaddr_2_reg_we),
                                               .uc2rb_desc_4_axaddr_3_reg_we(uc2rb_desc_4_axaddr_3_reg_we),
                                               .uc2rb_desc_4_axid_0_reg_we(uc2rb_desc_4_axid_0_reg_we),
                                               .uc2rb_desc_4_axid_1_reg_we(uc2rb_desc_4_axid_1_reg_we),
                                               .uc2rb_desc_4_axid_2_reg_we(uc2rb_desc_4_axid_2_reg_we),
                                               .uc2rb_desc_4_axid_3_reg_we(uc2rb_desc_4_axid_3_reg_we),
                                               .uc2rb_desc_4_axuser_0_reg_we(uc2rb_desc_4_axuser_0_reg_we),
                                               .uc2rb_desc_4_axuser_1_reg_we(uc2rb_desc_4_axuser_1_reg_we),
                                               .uc2rb_desc_4_axuser_2_reg_we(uc2rb_desc_4_axuser_2_reg_we),
                                               .uc2rb_desc_4_axuser_3_reg_we(uc2rb_desc_4_axuser_3_reg_we),
                                               .uc2rb_desc_4_axuser_4_reg_we(uc2rb_desc_4_axuser_4_reg_we),
                                               .uc2rb_desc_4_axuser_5_reg_we(uc2rb_desc_4_axuser_5_reg_we),
                                               .uc2rb_desc_4_axuser_6_reg_we(uc2rb_desc_4_axuser_6_reg_we),
                                               .uc2rb_desc_4_axuser_7_reg_we(uc2rb_desc_4_axuser_7_reg_we),
                                               .uc2rb_desc_4_axuser_8_reg_we(uc2rb_desc_4_axuser_8_reg_we),
                                               .uc2rb_desc_4_axuser_9_reg_we(uc2rb_desc_4_axuser_9_reg_we),
                                               .uc2rb_desc_4_axuser_10_reg_we(uc2rb_desc_4_axuser_10_reg_we),
                                               .uc2rb_desc_4_axuser_11_reg_we(uc2rb_desc_4_axuser_11_reg_we),
                                               .uc2rb_desc_4_axuser_12_reg_we(uc2rb_desc_4_axuser_12_reg_we),
                                               .uc2rb_desc_4_axuser_13_reg_we(uc2rb_desc_4_axuser_13_reg_we),
                                               .uc2rb_desc_4_axuser_14_reg_we(uc2rb_desc_4_axuser_14_reg_we),
                                               .uc2rb_desc_4_axuser_15_reg_we(uc2rb_desc_4_axuser_15_reg_we),
                                               .uc2rb_desc_4_wuser_0_reg_we(uc2rb_desc_4_wuser_0_reg_we),
                                               .uc2rb_desc_4_wuser_1_reg_we(uc2rb_desc_4_wuser_1_reg_we),
                                               .uc2rb_desc_4_wuser_2_reg_we(uc2rb_desc_4_wuser_2_reg_we),
                                               .uc2rb_desc_4_wuser_3_reg_we(uc2rb_desc_4_wuser_3_reg_we),
                                               .uc2rb_desc_4_wuser_4_reg_we(uc2rb_desc_4_wuser_4_reg_we),
                                               .uc2rb_desc_4_wuser_5_reg_we(uc2rb_desc_4_wuser_5_reg_we),
                                               .uc2rb_desc_4_wuser_6_reg_we(uc2rb_desc_4_wuser_6_reg_we),
                                               .uc2rb_desc_4_wuser_7_reg_we(uc2rb_desc_4_wuser_7_reg_we),
                                               .uc2rb_desc_4_wuser_8_reg_we(uc2rb_desc_4_wuser_8_reg_we),
                                               .uc2rb_desc_4_wuser_9_reg_we(uc2rb_desc_4_wuser_9_reg_we),
                                               .uc2rb_desc_4_wuser_10_reg_we(uc2rb_desc_4_wuser_10_reg_we),
                                               .uc2rb_desc_4_wuser_11_reg_we(uc2rb_desc_4_wuser_11_reg_we),
                                               .uc2rb_desc_4_wuser_12_reg_we(uc2rb_desc_4_wuser_12_reg_we),
                                               .uc2rb_desc_4_wuser_13_reg_we(uc2rb_desc_4_wuser_13_reg_we),
                                               .uc2rb_desc_4_wuser_14_reg_we(uc2rb_desc_4_wuser_14_reg_we),
                                               .uc2rb_desc_4_wuser_15_reg_we(uc2rb_desc_4_wuser_15_reg_we),
                                               .uc2rb_desc_5_txn_type_reg_we(uc2rb_desc_5_txn_type_reg_we),
                                               .uc2rb_desc_5_size_reg_we(uc2rb_desc_5_size_reg_we),
                                               .uc2rb_desc_5_data_offset_reg_we(uc2rb_desc_5_data_offset_reg_we),
                                               .uc2rb_desc_5_axsize_reg_we(uc2rb_desc_5_axsize_reg_we),
                                               .uc2rb_desc_5_attr_reg_we(uc2rb_desc_5_attr_reg_we),
                                               .uc2rb_desc_5_axaddr_0_reg_we(uc2rb_desc_5_axaddr_0_reg_we),
                                               .uc2rb_desc_5_axaddr_1_reg_we(uc2rb_desc_5_axaddr_1_reg_we),
                                               .uc2rb_desc_5_axaddr_2_reg_we(uc2rb_desc_5_axaddr_2_reg_we),
                                               .uc2rb_desc_5_axaddr_3_reg_we(uc2rb_desc_5_axaddr_3_reg_we),
                                               .uc2rb_desc_5_axid_0_reg_we(uc2rb_desc_5_axid_0_reg_we),
                                               .uc2rb_desc_5_axid_1_reg_we(uc2rb_desc_5_axid_1_reg_we),
                                               .uc2rb_desc_5_axid_2_reg_we(uc2rb_desc_5_axid_2_reg_we),
                                               .uc2rb_desc_5_axid_3_reg_we(uc2rb_desc_5_axid_3_reg_we),
                                               .uc2rb_desc_5_axuser_0_reg_we(uc2rb_desc_5_axuser_0_reg_we),
                                               .uc2rb_desc_5_axuser_1_reg_we(uc2rb_desc_5_axuser_1_reg_we),
                                               .uc2rb_desc_5_axuser_2_reg_we(uc2rb_desc_5_axuser_2_reg_we),
                                               .uc2rb_desc_5_axuser_3_reg_we(uc2rb_desc_5_axuser_3_reg_we),
                                               .uc2rb_desc_5_axuser_4_reg_we(uc2rb_desc_5_axuser_4_reg_we),
                                               .uc2rb_desc_5_axuser_5_reg_we(uc2rb_desc_5_axuser_5_reg_we),
                                               .uc2rb_desc_5_axuser_6_reg_we(uc2rb_desc_5_axuser_6_reg_we),
                                               .uc2rb_desc_5_axuser_7_reg_we(uc2rb_desc_5_axuser_7_reg_we),
                                               .uc2rb_desc_5_axuser_8_reg_we(uc2rb_desc_5_axuser_8_reg_we),
                                               .uc2rb_desc_5_axuser_9_reg_we(uc2rb_desc_5_axuser_9_reg_we),
                                               .uc2rb_desc_5_axuser_10_reg_we(uc2rb_desc_5_axuser_10_reg_we),
                                               .uc2rb_desc_5_axuser_11_reg_we(uc2rb_desc_5_axuser_11_reg_we),
                                               .uc2rb_desc_5_axuser_12_reg_we(uc2rb_desc_5_axuser_12_reg_we),
                                               .uc2rb_desc_5_axuser_13_reg_we(uc2rb_desc_5_axuser_13_reg_we),
                                               .uc2rb_desc_5_axuser_14_reg_we(uc2rb_desc_5_axuser_14_reg_we),
                                               .uc2rb_desc_5_axuser_15_reg_we(uc2rb_desc_5_axuser_15_reg_we),
                                               .uc2rb_desc_5_wuser_0_reg_we(uc2rb_desc_5_wuser_0_reg_we),
                                               .uc2rb_desc_5_wuser_1_reg_we(uc2rb_desc_5_wuser_1_reg_we),
                                               .uc2rb_desc_5_wuser_2_reg_we(uc2rb_desc_5_wuser_2_reg_we),
                                               .uc2rb_desc_5_wuser_3_reg_we(uc2rb_desc_5_wuser_3_reg_we),
                                               .uc2rb_desc_5_wuser_4_reg_we(uc2rb_desc_5_wuser_4_reg_we),
                                               .uc2rb_desc_5_wuser_5_reg_we(uc2rb_desc_5_wuser_5_reg_we),
                                               .uc2rb_desc_5_wuser_6_reg_we(uc2rb_desc_5_wuser_6_reg_we),
                                               .uc2rb_desc_5_wuser_7_reg_we(uc2rb_desc_5_wuser_7_reg_we),
                                               .uc2rb_desc_5_wuser_8_reg_we(uc2rb_desc_5_wuser_8_reg_we),
                                               .uc2rb_desc_5_wuser_9_reg_we(uc2rb_desc_5_wuser_9_reg_we),
                                               .uc2rb_desc_5_wuser_10_reg_we(uc2rb_desc_5_wuser_10_reg_we),
                                               .uc2rb_desc_5_wuser_11_reg_we(uc2rb_desc_5_wuser_11_reg_we),
                                               .uc2rb_desc_5_wuser_12_reg_we(uc2rb_desc_5_wuser_12_reg_we),
                                               .uc2rb_desc_5_wuser_13_reg_we(uc2rb_desc_5_wuser_13_reg_we),
                                               .uc2rb_desc_5_wuser_14_reg_we(uc2rb_desc_5_wuser_14_reg_we),
                                               .uc2rb_desc_5_wuser_15_reg_we(uc2rb_desc_5_wuser_15_reg_we),
                                               .uc2rb_desc_6_txn_type_reg_we(uc2rb_desc_6_txn_type_reg_we),
                                               .uc2rb_desc_6_size_reg_we(uc2rb_desc_6_size_reg_we),
                                               .uc2rb_desc_6_data_offset_reg_we(uc2rb_desc_6_data_offset_reg_we),
                                               .uc2rb_desc_6_axsize_reg_we(uc2rb_desc_6_axsize_reg_we),
                                               .uc2rb_desc_6_attr_reg_we(uc2rb_desc_6_attr_reg_we),
                                               .uc2rb_desc_6_axaddr_0_reg_we(uc2rb_desc_6_axaddr_0_reg_we),
                                               .uc2rb_desc_6_axaddr_1_reg_we(uc2rb_desc_6_axaddr_1_reg_we),
                                               .uc2rb_desc_6_axaddr_2_reg_we(uc2rb_desc_6_axaddr_2_reg_we),
                                               .uc2rb_desc_6_axaddr_3_reg_we(uc2rb_desc_6_axaddr_3_reg_we),
                                               .uc2rb_desc_6_axid_0_reg_we(uc2rb_desc_6_axid_0_reg_we),
                                               .uc2rb_desc_6_axid_1_reg_we(uc2rb_desc_6_axid_1_reg_we),
                                               .uc2rb_desc_6_axid_2_reg_we(uc2rb_desc_6_axid_2_reg_we),
                                               .uc2rb_desc_6_axid_3_reg_we(uc2rb_desc_6_axid_3_reg_we),
                                               .uc2rb_desc_6_axuser_0_reg_we(uc2rb_desc_6_axuser_0_reg_we),
                                               .uc2rb_desc_6_axuser_1_reg_we(uc2rb_desc_6_axuser_1_reg_we),
                                               .uc2rb_desc_6_axuser_2_reg_we(uc2rb_desc_6_axuser_2_reg_we),
                                               .uc2rb_desc_6_axuser_3_reg_we(uc2rb_desc_6_axuser_3_reg_we),
                                               .uc2rb_desc_6_axuser_4_reg_we(uc2rb_desc_6_axuser_4_reg_we),
                                               .uc2rb_desc_6_axuser_5_reg_we(uc2rb_desc_6_axuser_5_reg_we),
                                               .uc2rb_desc_6_axuser_6_reg_we(uc2rb_desc_6_axuser_6_reg_we),
                                               .uc2rb_desc_6_axuser_7_reg_we(uc2rb_desc_6_axuser_7_reg_we),
                                               .uc2rb_desc_6_axuser_8_reg_we(uc2rb_desc_6_axuser_8_reg_we),
                                               .uc2rb_desc_6_axuser_9_reg_we(uc2rb_desc_6_axuser_9_reg_we),
                                               .uc2rb_desc_6_axuser_10_reg_we(uc2rb_desc_6_axuser_10_reg_we),
                                               .uc2rb_desc_6_axuser_11_reg_we(uc2rb_desc_6_axuser_11_reg_we),
                                               .uc2rb_desc_6_axuser_12_reg_we(uc2rb_desc_6_axuser_12_reg_we),
                                               .uc2rb_desc_6_axuser_13_reg_we(uc2rb_desc_6_axuser_13_reg_we),
                                               .uc2rb_desc_6_axuser_14_reg_we(uc2rb_desc_6_axuser_14_reg_we),
                                               .uc2rb_desc_6_axuser_15_reg_we(uc2rb_desc_6_axuser_15_reg_we),
                                               .uc2rb_desc_6_wuser_0_reg_we(uc2rb_desc_6_wuser_0_reg_we),
                                               .uc2rb_desc_6_wuser_1_reg_we(uc2rb_desc_6_wuser_1_reg_we),
                                               .uc2rb_desc_6_wuser_2_reg_we(uc2rb_desc_6_wuser_2_reg_we),
                                               .uc2rb_desc_6_wuser_3_reg_we(uc2rb_desc_6_wuser_3_reg_we),
                                               .uc2rb_desc_6_wuser_4_reg_we(uc2rb_desc_6_wuser_4_reg_we),
                                               .uc2rb_desc_6_wuser_5_reg_we(uc2rb_desc_6_wuser_5_reg_we),
                                               .uc2rb_desc_6_wuser_6_reg_we(uc2rb_desc_6_wuser_6_reg_we),
                                               .uc2rb_desc_6_wuser_7_reg_we(uc2rb_desc_6_wuser_7_reg_we),
                                               .uc2rb_desc_6_wuser_8_reg_we(uc2rb_desc_6_wuser_8_reg_we),
                                               .uc2rb_desc_6_wuser_9_reg_we(uc2rb_desc_6_wuser_9_reg_we),
                                               .uc2rb_desc_6_wuser_10_reg_we(uc2rb_desc_6_wuser_10_reg_we),
                                               .uc2rb_desc_6_wuser_11_reg_we(uc2rb_desc_6_wuser_11_reg_we),
                                               .uc2rb_desc_6_wuser_12_reg_we(uc2rb_desc_6_wuser_12_reg_we),
                                               .uc2rb_desc_6_wuser_13_reg_we(uc2rb_desc_6_wuser_13_reg_we),
                                               .uc2rb_desc_6_wuser_14_reg_we(uc2rb_desc_6_wuser_14_reg_we),
                                               .uc2rb_desc_6_wuser_15_reg_we(uc2rb_desc_6_wuser_15_reg_we),
                                               .uc2rb_desc_7_txn_type_reg_we(uc2rb_desc_7_txn_type_reg_we),
                                               .uc2rb_desc_7_size_reg_we(uc2rb_desc_7_size_reg_we),
                                               .uc2rb_desc_7_data_offset_reg_we(uc2rb_desc_7_data_offset_reg_we),
                                               .uc2rb_desc_7_axsize_reg_we(uc2rb_desc_7_axsize_reg_we),
                                               .uc2rb_desc_7_attr_reg_we(uc2rb_desc_7_attr_reg_we),
                                               .uc2rb_desc_7_axaddr_0_reg_we(uc2rb_desc_7_axaddr_0_reg_we),
                                               .uc2rb_desc_7_axaddr_1_reg_we(uc2rb_desc_7_axaddr_1_reg_we),
                                               .uc2rb_desc_7_axaddr_2_reg_we(uc2rb_desc_7_axaddr_2_reg_we),
                                               .uc2rb_desc_7_axaddr_3_reg_we(uc2rb_desc_7_axaddr_3_reg_we),
                                               .uc2rb_desc_7_axid_0_reg_we(uc2rb_desc_7_axid_0_reg_we),
                                               .uc2rb_desc_7_axid_1_reg_we(uc2rb_desc_7_axid_1_reg_we),
                                               .uc2rb_desc_7_axid_2_reg_we(uc2rb_desc_7_axid_2_reg_we),
                                               .uc2rb_desc_7_axid_3_reg_we(uc2rb_desc_7_axid_3_reg_we),
                                               .uc2rb_desc_7_axuser_0_reg_we(uc2rb_desc_7_axuser_0_reg_we),
                                               .uc2rb_desc_7_axuser_1_reg_we(uc2rb_desc_7_axuser_1_reg_we),
                                               .uc2rb_desc_7_axuser_2_reg_we(uc2rb_desc_7_axuser_2_reg_we),
                                               .uc2rb_desc_7_axuser_3_reg_we(uc2rb_desc_7_axuser_3_reg_we),
                                               .uc2rb_desc_7_axuser_4_reg_we(uc2rb_desc_7_axuser_4_reg_we),
                                               .uc2rb_desc_7_axuser_5_reg_we(uc2rb_desc_7_axuser_5_reg_we),
                                               .uc2rb_desc_7_axuser_6_reg_we(uc2rb_desc_7_axuser_6_reg_we),
                                               .uc2rb_desc_7_axuser_7_reg_we(uc2rb_desc_7_axuser_7_reg_we),
                                               .uc2rb_desc_7_axuser_8_reg_we(uc2rb_desc_7_axuser_8_reg_we),
                                               .uc2rb_desc_7_axuser_9_reg_we(uc2rb_desc_7_axuser_9_reg_we),
                                               .uc2rb_desc_7_axuser_10_reg_we(uc2rb_desc_7_axuser_10_reg_we),
                                               .uc2rb_desc_7_axuser_11_reg_we(uc2rb_desc_7_axuser_11_reg_we),
                                               .uc2rb_desc_7_axuser_12_reg_we(uc2rb_desc_7_axuser_12_reg_we),
                                               .uc2rb_desc_7_axuser_13_reg_we(uc2rb_desc_7_axuser_13_reg_we),
                                               .uc2rb_desc_7_axuser_14_reg_we(uc2rb_desc_7_axuser_14_reg_we),
                                               .uc2rb_desc_7_axuser_15_reg_we(uc2rb_desc_7_axuser_15_reg_we),
                                               .uc2rb_desc_7_wuser_0_reg_we(uc2rb_desc_7_wuser_0_reg_we),
                                               .uc2rb_desc_7_wuser_1_reg_we(uc2rb_desc_7_wuser_1_reg_we),
                                               .uc2rb_desc_7_wuser_2_reg_we(uc2rb_desc_7_wuser_2_reg_we),
                                               .uc2rb_desc_7_wuser_3_reg_we(uc2rb_desc_7_wuser_3_reg_we),
                                               .uc2rb_desc_7_wuser_4_reg_we(uc2rb_desc_7_wuser_4_reg_we),
                                               .uc2rb_desc_7_wuser_5_reg_we(uc2rb_desc_7_wuser_5_reg_we),
                                               .uc2rb_desc_7_wuser_6_reg_we(uc2rb_desc_7_wuser_6_reg_we),
                                               .uc2rb_desc_7_wuser_7_reg_we(uc2rb_desc_7_wuser_7_reg_we),
                                               .uc2rb_desc_7_wuser_8_reg_we(uc2rb_desc_7_wuser_8_reg_we),
                                               .uc2rb_desc_7_wuser_9_reg_we(uc2rb_desc_7_wuser_9_reg_we),
                                               .uc2rb_desc_7_wuser_10_reg_we(uc2rb_desc_7_wuser_10_reg_we),
                                               .uc2rb_desc_7_wuser_11_reg_we(uc2rb_desc_7_wuser_11_reg_we),
                                               .uc2rb_desc_7_wuser_12_reg_we(uc2rb_desc_7_wuser_12_reg_we),
                                               .uc2rb_desc_7_wuser_13_reg_we(uc2rb_desc_7_wuser_13_reg_we),
                                               .uc2rb_desc_7_wuser_14_reg_we(uc2rb_desc_7_wuser_14_reg_we),
                                               .uc2rb_desc_7_wuser_15_reg_we(uc2rb_desc_7_wuser_15_reg_we),
                                               .uc2rb_desc_8_txn_type_reg_we(uc2rb_desc_8_txn_type_reg_we),
                                               .uc2rb_desc_8_size_reg_we(uc2rb_desc_8_size_reg_we),
                                               .uc2rb_desc_8_data_offset_reg_we(uc2rb_desc_8_data_offset_reg_we),
                                               .uc2rb_desc_8_axsize_reg_we(uc2rb_desc_8_axsize_reg_we),
                                               .uc2rb_desc_8_attr_reg_we(uc2rb_desc_8_attr_reg_we),
                                               .uc2rb_desc_8_axaddr_0_reg_we(uc2rb_desc_8_axaddr_0_reg_we),
                                               .uc2rb_desc_8_axaddr_1_reg_we(uc2rb_desc_8_axaddr_1_reg_we),
                                               .uc2rb_desc_8_axaddr_2_reg_we(uc2rb_desc_8_axaddr_2_reg_we),
                                               .uc2rb_desc_8_axaddr_3_reg_we(uc2rb_desc_8_axaddr_3_reg_we),
                                               .uc2rb_desc_8_axid_0_reg_we(uc2rb_desc_8_axid_0_reg_we),
                                               .uc2rb_desc_8_axid_1_reg_we(uc2rb_desc_8_axid_1_reg_we),
                                               .uc2rb_desc_8_axid_2_reg_we(uc2rb_desc_8_axid_2_reg_we),
                                               .uc2rb_desc_8_axid_3_reg_we(uc2rb_desc_8_axid_3_reg_we),
                                               .uc2rb_desc_8_axuser_0_reg_we(uc2rb_desc_8_axuser_0_reg_we),
                                               .uc2rb_desc_8_axuser_1_reg_we(uc2rb_desc_8_axuser_1_reg_we),
                                               .uc2rb_desc_8_axuser_2_reg_we(uc2rb_desc_8_axuser_2_reg_we),
                                               .uc2rb_desc_8_axuser_3_reg_we(uc2rb_desc_8_axuser_3_reg_we),
                                               .uc2rb_desc_8_axuser_4_reg_we(uc2rb_desc_8_axuser_4_reg_we),
                                               .uc2rb_desc_8_axuser_5_reg_we(uc2rb_desc_8_axuser_5_reg_we),
                                               .uc2rb_desc_8_axuser_6_reg_we(uc2rb_desc_8_axuser_6_reg_we),
                                               .uc2rb_desc_8_axuser_7_reg_we(uc2rb_desc_8_axuser_7_reg_we),
                                               .uc2rb_desc_8_axuser_8_reg_we(uc2rb_desc_8_axuser_8_reg_we),
                                               .uc2rb_desc_8_axuser_9_reg_we(uc2rb_desc_8_axuser_9_reg_we),
                                               .uc2rb_desc_8_axuser_10_reg_we(uc2rb_desc_8_axuser_10_reg_we),
                                               .uc2rb_desc_8_axuser_11_reg_we(uc2rb_desc_8_axuser_11_reg_we),
                                               .uc2rb_desc_8_axuser_12_reg_we(uc2rb_desc_8_axuser_12_reg_we),
                                               .uc2rb_desc_8_axuser_13_reg_we(uc2rb_desc_8_axuser_13_reg_we),
                                               .uc2rb_desc_8_axuser_14_reg_we(uc2rb_desc_8_axuser_14_reg_we),
                                               .uc2rb_desc_8_axuser_15_reg_we(uc2rb_desc_8_axuser_15_reg_we),
                                               .uc2rb_desc_8_wuser_0_reg_we(uc2rb_desc_8_wuser_0_reg_we),
                                               .uc2rb_desc_8_wuser_1_reg_we(uc2rb_desc_8_wuser_1_reg_we),
                                               .uc2rb_desc_8_wuser_2_reg_we(uc2rb_desc_8_wuser_2_reg_we),
                                               .uc2rb_desc_8_wuser_3_reg_we(uc2rb_desc_8_wuser_3_reg_we),
                                               .uc2rb_desc_8_wuser_4_reg_we(uc2rb_desc_8_wuser_4_reg_we),
                                               .uc2rb_desc_8_wuser_5_reg_we(uc2rb_desc_8_wuser_5_reg_we),
                                               .uc2rb_desc_8_wuser_6_reg_we(uc2rb_desc_8_wuser_6_reg_we),
                                               .uc2rb_desc_8_wuser_7_reg_we(uc2rb_desc_8_wuser_7_reg_we),
                                               .uc2rb_desc_8_wuser_8_reg_we(uc2rb_desc_8_wuser_8_reg_we),
                                               .uc2rb_desc_8_wuser_9_reg_we(uc2rb_desc_8_wuser_9_reg_we),
                                               .uc2rb_desc_8_wuser_10_reg_we(uc2rb_desc_8_wuser_10_reg_we),
                                               .uc2rb_desc_8_wuser_11_reg_we(uc2rb_desc_8_wuser_11_reg_we),
                                               .uc2rb_desc_8_wuser_12_reg_we(uc2rb_desc_8_wuser_12_reg_we),
                                               .uc2rb_desc_8_wuser_13_reg_we(uc2rb_desc_8_wuser_13_reg_we),
                                               .uc2rb_desc_8_wuser_14_reg_we(uc2rb_desc_8_wuser_14_reg_we),
                                               .uc2rb_desc_8_wuser_15_reg_we(uc2rb_desc_8_wuser_15_reg_we),
                                               .uc2rb_desc_9_txn_type_reg_we(uc2rb_desc_9_txn_type_reg_we),
                                               .uc2rb_desc_9_size_reg_we(uc2rb_desc_9_size_reg_we),
                                               .uc2rb_desc_9_data_offset_reg_we(uc2rb_desc_9_data_offset_reg_we),
                                               .uc2rb_desc_9_axsize_reg_we(uc2rb_desc_9_axsize_reg_we),
                                               .uc2rb_desc_9_attr_reg_we(uc2rb_desc_9_attr_reg_we),
                                               .uc2rb_desc_9_axaddr_0_reg_we(uc2rb_desc_9_axaddr_0_reg_we),
                                               .uc2rb_desc_9_axaddr_1_reg_we(uc2rb_desc_9_axaddr_1_reg_we),
                                               .uc2rb_desc_9_axaddr_2_reg_we(uc2rb_desc_9_axaddr_2_reg_we),
                                               .uc2rb_desc_9_axaddr_3_reg_we(uc2rb_desc_9_axaddr_3_reg_we),
                                               .uc2rb_desc_9_axid_0_reg_we(uc2rb_desc_9_axid_0_reg_we),
                                               .uc2rb_desc_9_axid_1_reg_we(uc2rb_desc_9_axid_1_reg_we),
                                               .uc2rb_desc_9_axid_2_reg_we(uc2rb_desc_9_axid_2_reg_we),
                                               .uc2rb_desc_9_axid_3_reg_we(uc2rb_desc_9_axid_3_reg_we),
                                               .uc2rb_desc_9_axuser_0_reg_we(uc2rb_desc_9_axuser_0_reg_we),
                                               .uc2rb_desc_9_axuser_1_reg_we(uc2rb_desc_9_axuser_1_reg_we),
                                               .uc2rb_desc_9_axuser_2_reg_we(uc2rb_desc_9_axuser_2_reg_we),
                                               .uc2rb_desc_9_axuser_3_reg_we(uc2rb_desc_9_axuser_3_reg_we),
                                               .uc2rb_desc_9_axuser_4_reg_we(uc2rb_desc_9_axuser_4_reg_we),
                                               .uc2rb_desc_9_axuser_5_reg_we(uc2rb_desc_9_axuser_5_reg_we),
                                               .uc2rb_desc_9_axuser_6_reg_we(uc2rb_desc_9_axuser_6_reg_we),
                                               .uc2rb_desc_9_axuser_7_reg_we(uc2rb_desc_9_axuser_7_reg_we),
                                               .uc2rb_desc_9_axuser_8_reg_we(uc2rb_desc_9_axuser_8_reg_we),
                                               .uc2rb_desc_9_axuser_9_reg_we(uc2rb_desc_9_axuser_9_reg_we),
                                               .uc2rb_desc_9_axuser_10_reg_we(uc2rb_desc_9_axuser_10_reg_we),
                                               .uc2rb_desc_9_axuser_11_reg_we(uc2rb_desc_9_axuser_11_reg_we),
                                               .uc2rb_desc_9_axuser_12_reg_we(uc2rb_desc_9_axuser_12_reg_we),
                                               .uc2rb_desc_9_axuser_13_reg_we(uc2rb_desc_9_axuser_13_reg_we),
                                               .uc2rb_desc_9_axuser_14_reg_we(uc2rb_desc_9_axuser_14_reg_we),
                                               .uc2rb_desc_9_axuser_15_reg_we(uc2rb_desc_9_axuser_15_reg_we),
                                               .uc2rb_desc_9_wuser_0_reg_we(uc2rb_desc_9_wuser_0_reg_we),
                                               .uc2rb_desc_9_wuser_1_reg_we(uc2rb_desc_9_wuser_1_reg_we),
                                               .uc2rb_desc_9_wuser_2_reg_we(uc2rb_desc_9_wuser_2_reg_we),
                                               .uc2rb_desc_9_wuser_3_reg_we(uc2rb_desc_9_wuser_3_reg_we),
                                               .uc2rb_desc_9_wuser_4_reg_we(uc2rb_desc_9_wuser_4_reg_we),
                                               .uc2rb_desc_9_wuser_5_reg_we(uc2rb_desc_9_wuser_5_reg_we),
                                               .uc2rb_desc_9_wuser_6_reg_we(uc2rb_desc_9_wuser_6_reg_we),
                                               .uc2rb_desc_9_wuser_7_reg_we(uc2rb_desc_9_wuser_7_reg_we),
                                               .uc2rb_desc_9_wuser_8_reg_we(uc2rb_desc_9_wuser_8_reg_we),
                                               .uc2rb_desc_9_wuser_9_reg_we(uc2rb_desc_9_wuser_9_reg_we),
                                               .uc2rb_desc_9_wuser_10_reg_we(uc2rb_desc_9_wuser_10_reg_we),
                                               .uc2rb_desc_9_wuser_11_reg_we(uc2rb_desc_9_wuser_11_reg_we),
                                               .uc2rb_desc_9_wuser_12_reg_we(uc2rb_desc_9_wuser_12_reg_we),
                                               .uc2rb_desc_9_wuser_13_reg_we(uc2rb_desc_9_wuser_13_reg_we),
                                               .uc2rb_desc_9_wuser_14_reg_we(uc2rb_desc_9_wuser_14_reg_we),
                                               .uc2rb_desc_9_wuser_15_reg_we(uc2rb_desc_9_wuser_15_reg_we),
                                               .uc2rb_desc_10_txn_type_reg_we(uc2rb_desc_10_txn_type_reg_we),
                                               .uc2rb_desc_10_size_reg_we(uc2rb_desc_10_size_reg_we),
                                               .uc2rb_desc_10_data_offset_reg_we(uc2rb_desc_10_data_offset_reg_we),
                                               .uc2rb_desc_10_axsize_reg_we(uc2rb_desc_10_axsize_reg_we),
                                               .uc2rb_desc_10_attr_reg_we(uc2rb_desc_10_attr_reg_we),
                                               .uc2rb_desc_10_axaddr_0_reg_we(uc2rb_desc_10_axaddr_0_reg_we),
                                               .uc2rb_desc_10_axaddr_1_reg_we(uc2rb_desc_10_axaddr_1_reg_we),
                                               .uc2rb_desc_10_axaddr_2_reg_we(uc2rb_desc_10_axaddr_2_reg_we),
                                               .uc2rb_desc_10_axaddr_3_reg_we(uc2rb_desc_10_axaddr_3_reg_we),
                                               .uc2rb_desc_10_axid_0_reg_we(uc2rb_desc_10_axid_0_reg_we),
                                               .uc2rb_desc_10_axid_1_reg_we(uc2rb_desc_10_axid_1_reg_we),
                                               .uc2rb_desc_10_axid_2_reg_we(uc2rb_desc_10_axid_2_reg_we),
                                               .uc2rb_desc_10_axid_3_reg_we(uc2rb_desc_10_axid_3_reg_we),
                                               .uc2rb_desc_10_axuser_0_reg_we(uc2rb_desc_10_axuser_0_reg_we),
                                               .uc2rb_desc_10_axuser_1_reg_we(uc2rb_desc_10_axuser_1_reg_we),
                                               .uc2rb_desc_10_axuser_2_reg_we(uc2rb_desc_10_axuser_2_reg_we),
                                               .uc2rb_desc_10_axuser_3_reg_we(uc2rb_desc_10_axuser_3_reg_we),
                                               .uc2rb_desc_10_axuser_4_reg_we(uc2rb_desc_10_axuser_4_reg_we),
                                               .uc2rb_desc_10_axuser_5_reg_we(uc2rb_desc_10_axuser_5_reg_we),
                                               .uc2rb_desc_10_axuser_6_reg_we(uc2rb_desc_10_axuser_6_reg_we),
                                               .uc2rb_desc_10_axuser_7_reg_we(uc2rb_desc_10_axuser_7_reg_we),
                                               .uc2rb_desc_10_axuser_8_reg_we(uc2rb_desc_10_axuser_8_reg_we),
                                               .uc2rb_desc_10_axuser_9_reg_we(uc2rb_desc_10_axuser_9_reg_we),
                                               .uc2rb_desc_10_axuser_10_reg_we(uc2rb_desc_10_axuser_10_reg_we),
                                               .uc2rb_desc_10_axuser_11_reg_we(uc2rb_desc_10_axuser_11_reg_we),
                                               .uc2rb_desc_10_axuser_12_reg_we(uc2rb_desc_10_axuser_12_reg_we),
                                               .uc2rb_desc_10_axuser_13_reg_we(uc2rb_desc_10_axuser_13_reg_we),
                                               .uc2rb_desc_10_axuser_14_reg_we(uc2rb_desc_10_axuser_14_reg_we),
                                               .uc2rb_desc_10_axuser_15_reg_we(uc2rb_desc_10_axuser_15_reg_we),
                                               .uc2rb_desc_10_wuser_0_reg_we(uc2rb_desc_10_wuser_0_reg_we),
                                               .uc2rb_desc_10_wuser_1_reg_we(uc2rb_desc_10_wuser_1_reg_we),
                                               .uc2rb_desc_10_wuser_2_reg_we(uc2rb_desc_10_wuser_2_reg_we),
                                               .uc2rb_desc_10_wuser_3_reg_we(uc2rb_desc_10_wuser_3_reg_we),
                                               .uc2rb_desc_10_wuser_4_reg_we(uc2rb_desc_10_wuser_4_reg_we),
                                               .uc2rb_desc_10_wuser_5_reg_we(uc2rb_desc_10_wuser_5_reg_we),
                                               .uc2rb_desc_10_wuser_6_reg_we(uc2rb_desc_10_wuser_6_reg_we),
                                               .uc2rb_desc_10_wuser_7_reg_we(uc2rb_desc_10_wuser_7_reg_we),
                                               .uc2rb_desc_10_wuser_8_reg_we(uc2rb_desc_10_wuser_8_reg_we),
                                               .uc2rb_desc_10_wuser_9_reg_we(uc2rb_desc_10_wuser_9_reg_we),
                                               .uc2rb_desc_10_wuser_10_reg_we(uc2rb_desc_10_wuser_10_reg_we),
                                               .uc2rb_desc_10_wuser_11_reg_we(uc2rb_desc_10_wuser_11_reg_we),
                                               .uc2rb_desc_10_wuser_12_reg_we(uc2rb_desc_10_wuser_12_reg_we),
                                               .uc2rb_desc_10_wuser_13_reg_we(uc2rb_desc_10_wuser_13_reg_we),
                                               .uc2rb_desc_10_wuser_14_reg_we(uc2rb_desc_10_wuser_14_reg_we),
                                               .uc2rb_desc_10_wuser_15_reg_we(uc2rb_desc_10_wuser_15_reg_we),
                                               .uc2rb_desc_11_txn_type_reg_we(uc2rb_desc_11_txn_type_reg_we),
                                               .uc2rb_desc_11_size_reg_we(uc2rb_desc_11_size_reg_we),
                                               .uc2rb_desc_11_data_offset_reg_we(uc2rb_desc_11_data_offset_reg_we),
                                               .uc2rb_desc_11_axsize_reg_we(uc2rb_desc_11_axsize_reg_we),
                                               .uc2rb_desc_11_attr_reg_we(uc2rb_desc_11_attr_reg_we),
                                               .uc2rb_desc_11_axaddr_0_reg_we(uc2rb_desc_11_axaddr_0_reg_we),
                                               .uc2rb_desc_11_axaddr_1_reg_we(uc2rb_desc_11_axaddr_1_reg_we),
                                               .uc2rb_desc_11_axaddr_2_reg_we(uc2rb_desc_11_axaddr_2_reg_we),
                                               .uc2rb_desc_11_axaddr_3_reg_we(uc2rb_desc_11_axaddr_3_reg_we),
                                               .uc2rb_desc_11_axid_0_reg_we(uc2rb_desc_11_axid_0_reg_we),
                                               .uc2rb_desc_11_axid_1_reg_we(uc2rb_desc_11_axid_1_reg_we),
                                               .uc2rb_desc_11_axid_2_reg_we(uc2rb_desc_11_axid_2_reg_we),
                                               .uc2rb_desc_11_axid_3_reg_we(uc2rb_desc_11_axid_3_reg_we),
                                               .uc2rb_desc_11_axuser_0_reg_we(uc2rb_desc_11_axuser_0_reg_we),
                                               .uc2rb_desc_11_axuser_1_reg_we(uc2rb_desc_11_axuser_1_reg_we),
                                               .uc2rb_desc_11_axuser_2_reg_we(uc2rb_desc_11_axuser_2_reg_we),
                                               .uc2rb_desc_11_axuser_3_reg_we(uc2rb_desc_11_axuser_3_reg_we),
                                               .uc2rb_desc_11_axuser_4_reg_we(uc2rb_desc_11_axuser_4_reg_we),
                                               .uc2rb_desc_11_axuser_5_reg_we(uc2rb_desc_11_axuser_5_reg_we),
                                               .uc2rb_desc_11_axuser_6_reg_we(uc2rb_desc_11_axuser_6_reg_we),
                                               .uc2rb_desc_11_axuser_7_reg_we(uc2rb_desc_11_axuser_7_reg_we),
                                               .uc2rb_desc_11_axuser_8_reg_we(uc2rb_desc_11_axuser_8_reg_we),
                                               .uc2rb_desc_11_axuser_9_reg_we(uc2rb_desc_11_axuser_9_reg_we),
                                               .uc2rb_desc_11_axuser_10_reg_we(uc2rb_desc_11_axuser_10_reg_we),
                                               .uc2rb_desc_11_axuser_11_reg_we(uc2rb_desc_11_axuser_11_reg_we),
                                               .uc2rb_desc_11_axuser_12_reg_we(uc2rb_desc_11_axuser_12_reg_we),
                                               .uc2rb_desc_11_axuser_13_reg_we(uc2rb_desc_11_axuser_13_reg_we),
                                               .uc2rb_desc_11_axuser_14_reg_we(uc2rb_desc_11_axuser_14_reg_we),
                                               .uc2rb_desc_11_axuser_15_reg_we(uc2rb_desc_11_axuser_15_reg_we),
                                               .uc2rb_desc_11_wuser_0_reg_we(uc2rb_desc_11_wuser_0_reg_we),
                                               .uc2rb_desc_11_wuser_1_reg_we(uc2rb_desc_11_wuser_1_reg_we),
                                               .uc2rb_desc_11_wuser_2_reg_we(uc2rb_desc_11_wuser_2_reg_we),
                                               .uc2rb_desc_11_wuser_3_reg_we(uc2rb_desc_11_wuser_3_reg_we),
                                               .uc2rb_desc_11_wuser_4_reg_we(uc2rb_desc_11_wuser_4_reg_we),
                                               .uc2rb_desc_11_wuser_5_reg_we(uc2rb_desc_11_wuser_5_reg_we),
                                               .uc2rb_desc_11_wuser_6_reg_we(uc2rb_desc_11_wuser_6_reg_we),
                                               .uc2rb_desc_11_wuser_7_reg_we(uc2rb_desc_11_wuser_7_reg_we),
                                               .uc2rb_desc_11_wuser_8_reg_we(uc2rb_desc_11_wuser_8_reg_we),
                                               .uc2rb_desc_11_wuser_9_reg_we(uc2rb_desc_11_wuser_9_reg_we),
                                               .uc2rb_desc_11_wuser_10_reg_we(uc2rb_desc_11_wuser_10_reg_we),
                                               .uc2rb_desc_11_wuser_11_reg_we(uc2rb_desc_11_wuser_11_reg_we),
                                               .uc2rb_desc_11_wuser_12_reg_we(uc2rb_desc_11_wuser_12_reg_we),
                                               .uc2rb_desc_11_wuser_13_reg_we(uc2rb_desc_11_wuser_13_reg_we),
                                               .uc2rb_desc_11_wuser_14_reg_we(uc2rb_desc_11_wuser_14_reg_we),
                                               .uc2rb_desc_11_wuser_15_reg_we(uc2rb_desc_11_wuser_15_reg_we),
                                               .uc2rb_desc_12_txn_type_reg_we(uc2rb_desc_12_txn_type_reg_we),
                                               .uc2rb_desc_12_size_reg_we(uc2rb_desc_12_size_reg_we),
                                               .uc2rb_desc_12_data_offset_reg_we(uc2rb_desc_12_data_offset_reg_we),
                                               .uc2rb_desc_12_axsize_reg_we(uc2rb_desc_12_axsize_reg_we),
                                               .uc2rb_desc_12_attr_reg_we(uc2rb_desc_12_attr_reg_we),
                                               .uc2rb_desc_12_axaddr_0_reg_we(uc2rb_desc_12_axaddr_0_reg_we),
                                               .uc2rb_desc_12_axaddr_1_reg_we(uc2rb_desc_12_axaddr_1_reg_we),
                                               .uc2rb_desc_12_axaddr_2_reg_we(uc2rb_desc_12_axaddr_2_reg_we),
                                               .uc2rb_desc_12_axaddr_3_reg_we(uc2rb_desc_12_axaddr_3_reg_we),
                                               .uc2rb_desc_12_axid_0_reg_we(uc2rb_desc_12_axid_0_reg_we),
                                               .uc2rb_desc_12_axid_1_reg_we(uc2rb_desc_12_axid_1_reg_we),
                                               .uc2rb_desc_12_axid_2_reg_we(uc2rb_desc_12_axid_2_reg_we),
                                               .uc2rb_desc_12_axid_3_reg_we(uc2rb_desc_12_axid_3_reg_we),
                                               .uc2rb_desc_12_axuser_0_reg_we(uc2rb_desc_12_axuser_0_reg_we),
                                               .uc2rb_desc_12_axuser_1_reg_we(uc2rb_desc_12_axuser_1_reg_we),
                                               .uc2rb_desc_12_axuser_2_reg_we(uc2rb_desc_12_axuser_2_reg_we),
                                               .uc2rb_desc_12_axuser_3_reg_we(uc2rb_desc_12_axuser_3_reg_we),
                                               .uc2rb_desc_12_axuser_4_reg_we(uc2rb_desc_12_axuser_4_reg_we),
                                               .uc2rb_desc_12_axuser_5_reg_we(uc2rb_desc_12_axuser_5_reg_we),
                                               .uc2rb_desc_12_axuser_6_reg_we(uc2rb_desc_12_axuser_6_reg_we),
                                               .uc2rb_desc_12_axuser_7_reg_we(uc2rb_desc_12_axuser_7_reg_we),
                                               .uc2rb_desc_12_axuser_8_reg_we(uc2rb_desc_12_axuser_8_reg_we),
                                               .uc2rb_desc_12_axuser_9_reg_we(uc2rb_desc_12_axuser_9_reg_we),
                                               .uc2rb_desc_12_axuser_10_reg_we(uc2rb_desc_12_axuser_10_reg_we),
                                               .uc2rb_desc_12_axuser_11_reg_we(uc2rb_desc_12_axuser_11_reg_we),
                                               .uc2rb_desc_12_axuser_12_reg_we(uc2rb_desc_12_axuser_12_reg_we),
                                               .uc2rb_desc_12_axuser_13_reg_we(uc2rb_desc_12_axuser_13_reg_we),
                                               .uc2rb_desc_12_axuser_14_reg_we(uc2rb_desc_12_axuser_14_reg_we),
                                               .uc2rb_desc_12_axuser_15_reg_we(uc2rb_desc_12_axuser_15_reg_we),
                                               .uc2rb_desc_12_wuser_0_reg_we(uc2rb_desc_12_wuser_0_reg_we),
                                               .uc2rb_desc_12_wuser_1_reg_we(uc2rb_desc_12_wuser_1_reg_we),
                                               .uc2rb_desc_12_wuser_2_reg_we(uc2rb_desc_12_wuser_2_reg_we),
                                               .uc2rb_desc_12_wuser_3_reg_we(uc2rb_desc_12_wuser_3_reg_we),
                                               .uc2rb_desc_12_wuser_4_reg_we(uc2rb_desc_12_wuser_4_reg_we),
                                               .uc2rb_desc_12_wuser_5_reg_we(uc2rb_desc_12_wuser_5_reg_we),
                                               .uc2rb_desc_12_wuser_6_reg_we(uc2rb_desc_12_wuser_6_reg_we),
                                               .uc2rb_desc_12_wuser_7_reg_we(uc2rb_desc_12_wuser_7_reg_we),
                                               .uc2rb_desc_12_wuser_8_reg_we(uc2rb_desc_12_wuser_8_reg_we),
                                               .uc2rb_desc_12_wuser_9_reg_we(uc2rb_desc_12_wuser_9_reg_we),
                                               .uc2rb_desc_12_wuser_10_reg_we(uc2rb_desc_12_wuser_10_reg_we),
                                               .uc2rb_desc_12_wuser_11_reg_we(uc2rb_desc_12_wuser_11_reg_we),
                                               .uc2rb_desc_12_wuser_12_reg_we(uc2rb_desc_12_wuser_12_reg_we),
                                               .uc2rb_desc_12_wuser_13_reg_we(uc2rb_desc_12_wuser_13_reg_we),
                                               .uc2rb_desc_12_wuser_14_reg_we(uc2rb_desc_12_wuser_14_reg_we),
                                               .uc2rb_desc_12_wuser_15_reg_we(uc2rb_desc_12_wuser_15_reg_we),
                                               .uc2rb_desc_13_txn_type_reg_we(uc2rb_desc_13_txn_type_reg_we),
                                               .uc2rb_desc_13_size_reg_we(uc2rb_desc_13_size_reg_we),
                                               .uc2rb_desc_13_data_offset_reg_we(uc2rb_desc_13_data_offset_reg_we),
                                               .uc2rb_desc_13_axsize_reg_we(uc2rb_desc_13_axsize_reg_we),
                                               .uc2rb_desc_13_attr_reg_we(uc2rb_desc_13_attr_reg_we),
                                               .uc2rb_desc_13_axaddr_0_reg_we(uc2rb_desc_13_axaddr_0_reg_we),
                                               .uc2rb_desc_13_axaddr_1_reg_we(uc2rb_desc_13_axaddr_1_reg_we),
                                               .uc2rb_desc_13_axaddr_2_reg_we(uc2rb_desc_13_axaddr_2_reg_we),
                                               .uc2rb_desc_13_axaddr_3_reg_we(uc2rb_desc_13_axaddr_3_reg_we),
                                               .uc2rb_desc_13_axid_0_reg_we(uc2rb_desc_13_axid_0_reg_we),
                                               .uc2rb_desc_13_axid_1_reg_we(uc2rb_desc_13_axid_1_reg_we),
                                               .uc2rb_desc_13_axid_2_reg_we(uc2rb_desc_13_axid_2_reg_we),
                                               .uc2rb_desc_13_axid_3_reg_we(uc2rb_desc_13_axid_3_reg_we),
                                               .uc2rb_desc_13_axuser_0_reg_we(uc2rb_desc_13_axuser_0_reg_we),
                                               .uc2rb_desc_13_axuser_1_reg_we(uc2rb_desc_13_axuser_1_reg_we),
                                               .uc2rb_desc_13_axuser_2_reg_we(uc2rb_desc_13_axuser_2_reg_we),
                                               .uc2rb_desc_13_axuser_3_reg_we(uc2rb_desc_13_axuser_3_reg_we),
                                               .uc2rb_desc_13_axuser_4_reg_we(uc2rb_desc_13_axuser_4_reg_we),
                                               .uc2rb_desc_13_axuser_5_reg_we(uc2rb_desc_13_axuser_5_reg_we),
                                               .uc2rb_desc_13_axuser_6_reg_we(uc2rb_desc_13_axuser_6_reg_we),
                                               .uc2rb_desc_13_axuser_7_reg_we(uc2rb_desc_13_axuser_7_reg_we),
                                               .uc2rb_desc_13_axuser_8_reg_we(uc2rb_desc_13_axuser_8_reg_we),
                                               .uc2rb_desc_13_axuser_9_reg_we(uc2rb_desc_13_axuser_9_reg_we),
                                               .uc2rb_desc_13_axuser_10_reg_we(uc2rb_desc_13_axuser_10_reg_we),
                                               .uc2rb_desc_13_axuser_11_reg_we(uc2rb_desc_13_axuser_11_reg_we),
                                               .uc2rb_desc_13_axuser_12_reg_we(uc2rb_desc_13_axuser_12_reg_we),
                                               .uc2rb_desc_13_axuser_13_reg_we(uc2rb_desc_13_axuser_13_reg_we),
                                               .uc2rb_desc_13_axuser_14_reg_we(uc2rb_desc_13_axuser_14_reg_we),
                                               .uc2rb_desc_13_axuser_15_reg_we(uc2rb_desc_13_axuser_15_reg_we),
                                               .uc2rb_desc_13_wuser_0_reg_we(uc2rb_desc_13_wuser_0_reg_we),
                                               .uc2rb_desc_13_wuser_1_reg_we(uc2rb_desc_13_wuser_1_reg_we),
                                               .uc2rb_desc_13_wuser_2_reg_we(uc2rb_desc_13_wuser_2_reg_we),
                                               .uc2rb_desc_13_wuser_3_reg_we(uc2rb_desc_13_wuser_3_reg_we),
                                               .uc2rb_desc_13_wuser_4_reg_we(uc2rb_desc_13_wuser_4_reg_we),
                                               .uc2rb_desc_13_wuser_5_reg_we(uc2rb_desc_13_wuser_5_reg_we),
                                               .uc2rb_desc_13_wuser_6_reg_we(uc2rb_desc_13_wuser_6_reg_we),
                                               .uc2rb_desc_13_wuser_7_reg_we(uc2rb_desc_13_wuser_7_reg_we),
                                               .uc2rb_desc_13_wuser_8_reg_we(uc2rb_desc_13_wuser_8_reg_we),
                                               .uc2rb_desc_13_wuser_9_reg_we(uc2rb_desc_13_wuser_9_reg_we),
                                               .uc2rb_desc_13_wuser_10_reg_we(uc2rb_desc_13_wuser_10_reg_we),
                                               .uc2rb_desc_13_wuser_11_reg_we(uc2rb_desc_13_wuser_11_reg_we),
                                               .uc2rb_desc_13_wuser_12_reg_we(uc2rb_desc_13_wuser_12_reg_we),
                                               .uc2rb_desc_13_wuser_13_reg_we(uc2rb_desc_13_wuser_13_reg_we),
                                               .uc2rb_desc_13_wuser_14_reg_we(uc2rb_desc_13_wuser_14_reg_we),
                                               .uc2rb_desc_13_wuser_15_reg_we(uc2rb_desc_13_wuser_15_reg_we),
                                               .uc2rb_desc_14_txn_type_reg_we(uc2rb_desc_14_txn_type_reg_we),
                                               .uc2rb_desc_14_size_reg_we(uc2rb_desc_14_size_reg_we),
                                               .uc2rb_desc_14_data_offset_reg_we(uc2rb_desc_14_data_offset_reg_we),
                                               .uc2rb_desc_14_axsize_reg_we(uc2rb_desc_14_axsize_reg_we),
                                               .uc2rb_desc_14_attr_reg_we(uc2rb_desc_14_attr_reg_we),
                                               .uc2rb_desc_14_axaddr_0_reg_we(uc2rb_desc_14_axaddr_0_reg_we),
                                               .uc2rb_desc_14_axaddr_1_reg_we(uc2rb_desc_14_axaddr_1_reg_we),
                                               .uc2rb_desc_14_axaddr_2_reg_we(uc2rb_desc_14_axaddr_2_reg_we),
                                               .uc2rb_desc_14_axaddr_3_reg_we(uc2rb_desc_14_axaddr_3_reg_we),
                                               .uc2rb_desc_14_axid_0_reg_we(uc2rb_desc_14_axid_0_reg_we),
                                               .uc2rb_desc_14_axid_1_reg_we(uc2rb_desc_14_axid_1_reg_we),
                                               .uc2rb_desc_14_axid_2_reg_we(uc2rb_desc_14_axid_2_reg_we),
                                               .uc2rb_desc_14_axid_3_reg_we(uc2rb_desc_14_axid_3_reg_we),
                                               .uc2rb_desc_14_axuser_0_reg_we(uc2rb_desc_14_axuser_0_reg_we),
                                               .uc2rb_desc_14_axuser_1_reg_we(uc2rb_desc_14_axuser_1_reg_we),
                                               .uc2rb_desc_14_axuser_2_reg_we(uc2rb_desc_14_axuser_2_reg_we),
                                               .uc2rb_desc_14_axuser_3_reg_we(uc2rb_desc_14_axuser_3_reg_we),
                                               .uc2rb_desc_14_axuser_4_reg_we(uc2rb_desc_14_axuser_4_reg_we),
                                               .uc2rb_desc_14_axuser_5_reg_we(uc2rb_desc_14_axuser_5_reg_we),
                                               .uc2rb_desc_14_axuser_6_reg_we(uc2rb_desc_14_axuser_6_reg_we),
                                               .uc2rb_desc_14_axuser_7_reg_we(uc2rb_desc_14_axuser_7_reg_we),
                                               .uc2rb_desc_14_axuser_8_reg_we(uc2rb_desc_14_axuser_8_reg_we),
                                               .uc2rb_desc_14_axuser_9_reg_we(uc2rb_desc_14_axuser_9_reg_we),
                                               .uc2rb_desc_14_axuser_10_reg_we(uc2rb_desc_14_axuser_10_reg_we),
                                               .uc2rb_desc_14_axuser_11_reg_we(uc2rb_desc_14_axuser_11_reg_we),
                                               .uc2rb_desc_14_axuser_12_reg_we(uc2rb_desc_14_axuser_12_reg_we),
                                               .uc2rb_desc_14_axuser_13_reg_we(uc2rb_desc_14_axuser_13_reg_we),
                                               .uc2rb_desc_14_axuser_14_reg_we(uc2rb_desc_14_axuser_14_reg_we),
                                               .uc2rb_desc_14_axuser_15_reg_we(uc2rb_desc_14_axuser_15_reg_we),
                                               .uc2rb_desc_14_wuser_0_reg_we(uc2rb_desc_14_wuser_0_reg_we),
                                               .uc2rb_desc_14_wuser_1_reg_we(uc2rb_desc_14_wuser_1_reg_we),
                                               .uc2rb_desc_14_wuser_2_reg_we(uc2rb_desc_14_wuser_2_reg_we),
                                               .uc2rb_desc_14_wuser_3_reg_we(uc2rb_desc_14_wuser_3_reg_we),
                                               .uc2rb_desc_14_wuser_4_reg_we(uc2rb_desc_14_wuser_4_reg_we),
                                               .uc2rb_desc_14_wuser_5_reg_we(uc2rb_desc_14_wuser_5_reg_we),
                                               .uc2rb_desc_14_wuser_6_reg_we(uc2rb_desc_14_wuser_6_reg_we),
                                               .uc2rb_desc_14_wuser_7_reg_we(uc2rb_desc_14_wuser_7_reg_we),
                                               .uc2rb_desc_14_wuser_8_reg_we(uc2rb_desc_14_wuser_8_reg_we),
                                               .uc2rb_desc_14_wuser_9_reg_we(uc2rb_desc_14_wuser_9_reg_we),
                                               .uc2rb_desc_14_wuser_10_reg_we(uc2rb_desc_14_wuser_10_reg_we),
                                               .uc2rb_desc_14_wuser_11_reg_we(uc2rb_desc_14_wuser_11_reg_we),
                                               .uc2rb_desc_14_wuser_12_reg_we(uc2rb_desc_14_wuser_12_reg_we),
                                               .uc2rb_desc_14_wuser_13_reg_we(uc2rb_desc_14_wuser_13_reg_we),
                                               .uc2rb_desc_14_wuser_14_reg_we(uc2rb_desc_14_wuser_14_reg_we),
                                               .uc2rb_desc_14_wuser_15_reg_we(uc2rb_desc_14_wuser_15_reg_we),
                                               .uc2rb_desc_15_txn_type_reg_we(uc2rb_desc_15_txn_type_reg_we),
                                               .uc2rb_desc_15_size_reg_we(uc2rb_desc_15_size_reg_we),
                                               .uc2rb_desc_15_data_offset_reg_we(uc2rb_desc_15_data_offset_reg_we),
                                               .uc2rb_desc_15_axsize_reg_we(uc2rb_desc_15_axsize_reg_we),
                                               .uc2rb_desc_15_attr_reg_we(uc2rb_desc_15_attr_reg_we),
                                               .uc2rb_desc_15_axaddr_0_reg_we(uc2rb_desc_15_axaddr_0_reg_we),
                                               .uc2rb_desc_15_axaddr_1_reg_we(uc2rb_desc_15_axaddr_1_reg_we),
                                               .uc2rb_desc_15_axaddr_2_reg_we(uc2rb_desc_15_axaddr_2_reg_we),
                                               .uc2rb_desc_15_axaddr_3_reg_we(uc2rb_desc_15_axaddr_3_reg_we),
                                               .uc2rb_desc_15_axid_0_reg_we(uc2rb_desc_15_axid_0_reg_we),
                                               .uc2rb_desc_15_axid_1_reg_we(uc2rb_desc_15_axid_1_reg_we),
                                               .uc2rb_desc_15_axid_2_reg_we(uc2rb_desc_15_axid_2_reg_we),
                                               .uc2rb_desc_15_axid_3_reg_we(uc2rb_desc_15_axid_3_reg_we),
                                               .uc2rb_desc_15_axuser_0_reg_we(uc2rb_desc_15_axuser_0_reg_we),
                                               .uc2rb_desc_15_axuser_1_reg_we(uc2rb_desc_15_axuser_1_reg_we),
                                               .uc2rb_desc_15_axuser_2_reg_we(uc2rb_desc_15_axuser_2_reg_we),
                                               .uc2rb_desc_15_axuser_3_reg_we(uc2rb_desc_15_axuser_3_reg_we),
                                               .uc2rb_desc_15_axuser_4_reg_we(uc2rb_desc_15_axuser_4_reg_we),
                                               .uc2rb_desc_15_axuser_5_reg_we(uc2rb_desc_15_axuser_5_reg_we),
                                               .uc2rb_desc_15_axuser_6_reg_we(uc2rb_desc_15_axuser_6_reg_we),
                                               .uc2rb_desc_15_axuser_7_reg_we(uc2rb_desc_15_axuser_7_reg_we),
                                               .uc2rb_desc_15_axuser_8_reg_we(uc2rb_desc_15_axuser_8_reg_we),
                                               .uc2rb_desc_15_axuser_9_reg_we(uc2rb_desc_15_axuser_9_reg_we),
                                               .uc2rb_desc_15_axuser_10_reg_we(uc2rb_desc_15_axuser_10_reg_we),
                                               .uc2rb_desc_15_axuser_11_reg_we(uc2rb_desc_15_axuser_11_reg_we),
                                               .uc2rb_desc_15_axuser_12_reg_we(uc2rb_desc_15_axuser_12_reg_we),
                                               .uc2rb_desc_15_axuser_13_reg_we(uc2rb_desc_15_axuser_13_reg_we),
                                               .uc2rb_desc_15_axuser_14_reg_we(uc2rb_desc_15_axuser_14_reg_we),
                                               .uc2rb_desc_15_axuser_15_reg_we(uc2rb_desc_15_axuser_15_reg_we),
                                               .uc2rb_desc_15_wuser_0_reg_we(uc2rb_desc_15_wuser_0_reg_we),
                                               .uc2rb_desc_15_wuser_1_reg_we(uc2rb_desc_15_wuser_1_reg_we),
                                               .uc2rb_desc_15_wuser_2_reg_we(uc2rb_desc_15_wuser_2_reg_we),
                                               .uc2rb_desc_15_wuser_3_reg_we(uc2rb_desc_15_wuser_3_reg_we),
                                               .uc2rb_desc_15_wuser_4_reg_we(uc2rb_desc_15_wuser_4_reg_we),
                                               .uc2rb_desc_15_wuser_5_reg_we(uc2rb_desc_15_wuser_5_reg_we),
                                               .uc2rb_desc_15_wuser_6_reg_we(uc2rb_desc_15_wuser_6_reg_we),
                                               .uc2rb_desc_15_wuser_7_reg_we(uc2rb_desc_15_wuser_7_reg_we),
                                               .uc2rb_desc_15_wuser_8_reg_we(uc2rb_desc_15_wuser_8_reg_we),
                                               .uc2rb_desc_15_wuser_9_reg_we(uc2rb_desc_15_wuser_9_reg_we),
                                               .uc2rb_desc_15_wuser_10_reg_we(uc2rb_desc_15_wuser_10_reg_we),
                                               .uc2rb_desc_15_wuser_11_reg_we(uc2rb_desc_15_wuser_11_reg_we),
                                               .uc2rb_desc_15_wuser_12_reg_we(uc2rb_desc_15_wuser_12_reg_we),
                                               .uc2rb_desc_15_wuser_13_reg_we(uc2rb_desc_15_wuser_13_reg_we),
                                               .uc2rb_desc_15_wuser_14_reg_we(uc2rb_desc_15_wuser_14_reg_we),
                                               .uc2rb_desc_15_wuser_15_reg_we(uc2rb_desc_15_wuser_15_reg_we),
                                               .uc2rb_rd_addr   (uc2rb_rd_addr),
                                               .uc2rb_wr_we     (uc2rb_wr_we),
                                               .uc2rb_wr_bwe    (uc2rb_wr_bwe),
                                               .uc2rb_wr_addr   (uc2rb_wr_addr),
                                               .uc2rb_wr_data   (uc2rb_wr_data),
                                               .uc2rb_wr_wstrb  (uc2rb_wr_wstrb),
                                               .uc2hm_trig      (uc2hm_trig),
                                               // Inputs
                                               .axi_aclk        (axi_aclk),
                                               .axi_aresetn     (rst_n),

                                               .version_reg     (version_reg),
                                               .bridge_type_reg (bridge_type_reg),
                                               .mode_select_reg (mode_select_reg),
                                               .reset_reg       (reset_reg),
                                               .axi_bridge_config_reg(axi_bridge_config_reg),
                                               .axi_max_desc_reg(axi_max_desc_reg),
                                               .intr_status_reg (intr_status_reg),
                                               .intr_error_status_reg(intr_error_status_reg),
                                               .intr_error_clear_reg(intr_error_clear_reg),
                                               .intr_error_enable_reg(intr_error_enable_reg),
                                               .addr_in_0_reg   (addr_in_0_reg),
                                               .addr_in_1_reg   (addr_in_1_reg),
                                               .addr_in_2_reg   (addr_in_2_reg),
                                               .addr_in_3_reg   (addr_in_3_reg),
                                               .trans_mask_0_reg(trans_mask_0_reg),
                                               .trans_mask_1_reg(trans_mask_1_reg),
                                               .trans_mask_2_reg(trans_mask_2_reg),
                                               .trans_mask_3_reg(trans_mask_3_reg),
                                               .trans_addr_0_reg(trans_addr_0_reg),
                                               .trans_addr_1_reg(trans_addr_1_reg),
                                               .trans_addr_2_reg(trans_addr_2_reg),
                                               .trans_addr_3_reg(trans_addr_3_reg),
                                               .ownership_reg   (ownership_reg),
                                               .ownership_flip_reg(ownership_flip_reg),
                                               .status_resp_reg (status_resp_reg),
                                               .intr_txn_avail_status_reg(intr_txn_avail_status_reg),
                                               .intr_txn_avail_clear_reg(intr_txn_avail_clear_reg),
                                               .intr_txn_avail_enable_reg(intr_txn_avail_enable_reg),
                                               .intr_comp_status_reg(intr_comp_status_reg),
                                               .intr_comp_clear_reg(intr_comp_clear_reg),
                                               .intr_comp_enable_reg(intr_comp_enable_reg),
                                               .status_resp_comp_reg(status_resp_comp_reg),
                                               .status_busy_reg (status_busy_reg),
                                               .resp_fifo_free_level_reg(resp_fifo_free_level_reg),
                                               .resp_order_reg(resp_order_reg),
                                               .desc_0_txn_type_reg(desc_0_txn_type_reg),
                                               .desc_0_size_reg (desc_0_size_reg),
                                               .desc_0_data_offset_reg(desc_0_data_offset_reg),
                                               .desc_0_data_host_addr_0_reg(desc_0_data_host_addr_0_reg),
                                               .desc_0_data_host_addr_1_reg(desc_0_data_host_addr_1_reg),
                                               .desc_0_data_host_addr_2_reg(desc_0_data_host_addr_2_reg),
                                               .desc_0_data_host_addr_3_reg(desc_0_data_host_addr_3_reg),
                                               .desc_0_wstrb_host_addr_0_reg(desc_0_wstrb_host_addr_0_reg),
                                               .desc_0_wstrb_host_addr_1_reg(desc_0_wstrb_host_addr_1_reg),
                                               .desc_0_wstrb_host_addr_2_reg(desc_0_wstrb_host_addr_2_reg),
                                               .desc_0_wstrb_host_addr_3_reg(desc_0_wstrb_host_addr_3_reg),
                                               .desc_0_axsize_reg(desc_0_axsize_reg),
                                               .desc_0_attr_reg (desc_0_attr_reg),
                                               .desc_0_axaddr_0_reg(desc_0_axaddr_0_reg),
                                               .desc_0_axaddr_1_reg(desc_0_axaddr_1_reg),
                                               .desc_0_axaddr_2_reg(desc_0_axaddr_2_reg),
                                               .desc_0_axaddr_3_reg(desc_0_axaddr_3_reg),
                                               .desc_0_axid_0_reg(desc_0_axid_0_reg),
                                               .desc_0_axid_1_reg(desc_0_axid_1_reg),
                                               .desc_0_axid_2_reg(desc_0_axid_2_reg),
                                               .desc_0_axid_3_reg(desc_0_axid_3_reg),
                                               .desc_0_axuser_0_reg(desc_0_axuser_0_reg),
                                               .desc_0_axuser_1_reg(desc_0_axuser_1_reg),
                                               .desc_0_axuser_2_reg(desc_0_axuser_2_reg),
                                               .desc_0_axuser_3_reg(desc_0_axuser_3_reg),
                                               .desc_0_axuser_4_reg(desc_0_axuser_4_reg),
                                               .desc_0_axuser_5_reg(desc_0_axuser_5_reg),
                                               .desc_0_axuser_6_reg(desc_0_axuser_6_reg),
                                               .desc_0_axuser_7_reg(desc_0_axuser_7_reg),
                                               .desc_0_axuser_8_reg(desc_0_axuser_8_reg),
                                               .desc_0_axuser_9_reg(desc_0_axuser_9_reg),
                                               .desc_0_axuser_10_reg(desc_0_axuser_10_reg),
                                               .desc_0_axuser_11_reg(desc_0_axuser_11_reg),
                                               .desc_0_axuser_12_reg(desc_0_axuser_12_reg),
                                               .desc_0_axuser_13_reg(desc_0_axuser_13_reg),
                                               .desc_0_axuser_14_reg(desc_0_axuser_14_reg),
                                               .desc_0_axuser_15_reg(desc_0_axuser_15_reg),
                                               .desc_0_xuser_0_reg(desc_0_xuser_0_reg),
                                               .desc_0_xuser_1_reg(desc_0_xuser_1_reg),
                                               .desc_0_xuser_2_reg(desc_0_xuser_2_reg),
                                               .desc_0_xuser_3_reg(desc_0_xuser_3_reg),
                                               .desc_0_xuser_4_reg(desc_0_xuser_4_reg),
                                               .desc_0_xuser_5_reg(desc_0_xuser_5_reg),
                                               .desc_0_xuser_6_reg(desc_0_xuser_6_reg),
                                               .desc_0_xuser_7_reg(desc_0_xuser_7_reg),
                                               .desc_0_xuser_8_reg(desc_0_xuser_8_reg),
                                               .desc_0_xuser_9_reg(desc_0_xuser_9_reg),
                                               .desc_0_xuser_10_reg(desc_0_xuser_10_reg),
                                               .desc_0_xuser_11_reg(desc_0_xuser_11_reg),
                                               .desc_0_xuser_12_reg(desc_0_xuser_12_reg),
                                               .desc_0_xuser_13_reg(desc_0_xuser_13_reg),
                                               .desc_0_xuser_14_reg(desc_0_xuser_14_reg),
                                               .desc_0_xuser_15_reg(desc_0_xuser_15_reg),
                                               .desc_0_wuser_0_reg(desc_0_wuser_0_reg),
                                               .desc_0_wuser_1_reg(desc_0_wuser_1_reg),
                                               .desc_0_wuser_2_reg(desc_0_wuser_2_reg),
                                               .desc_0_wuser_3_reg(desc_0_wuser_3_reg),
                                               .desc_0_wuser_4_reg(desc_0_wuser_4_reg),
                                               .desc_0_wuser_5_reg(desc_0_wuser_5_reg),
                                               .desc_0_wuser_6_reg(desc_0_wuser_6_reg),
                                               .desc_0_wuser_7_reg(desc_0_wuser_7_reg),
                                               .desc_0_wuser_8_reg(desc_0_wuser_8_reg),
                                               .desc_0_wuser_9_reg(desc_0_wuser_9_reg),
                                               .desc_0_wuser_10_reg(desc_0_wuser_10_reg),
                                               .desc_0_wuser_11_reg(desc_0_wuser_11_reg),
                                               .desc_0_wuser_12_reg(desc_0_wuser_12_reg),
                                               .desc_0_wuser_13_reg(desc_0_wuser_13_reg),
                                               .desc_0_wuser_14_reg(desc_0_wuser_14_reg),
                                               .desc_0_wuser_15_reg(desc_0_wuser_15_reg),
                                               .desc_1_txn_type_reg(desc_1_txn_type_reg),
                                               .desc_1_size_reg (desc_1_size_reg),
                                               .desc_1_data_offset_reg(desc_1_data_offset_reg),
                                               .desc_1_data_host_addr_0_reg(desc_1_data_host_addr_0_reg),
                                               .desc_1_data_host_addr_1_reg(desc_1_data_host_addr_1_reg),
                                               .desc_1_data_host_addr_2_reg(desc_1_data_host_addr_2_reg),
                                               .desc_1_data_host_addr_3_reg(desc_1_data_host_addr_3_reg),
                                               .desc_1_wstrb_host_addr_0_reg(desc_1_wstrb_host_addr_0_reg),
                                               .desc_1_wstrb_host_addr_1_reg(desc_1_wstrb_host_addr_1_reg),
                                               .desc_1_wstrb_host_addr_2_reg(desc_1_wstrb_host_addr_2_reg),
                                               .desc_1_wstrb_host_addr_3_reg(desc_1_wstrb_host_addr_3_reg),
                                               .desc_1_axsize_reg(desc_1_axsize_reg),
                                               .desc_1_attr_reg (desc_1_attr_reg),
                                               .desc_1_axaddr_0_reg(desc_1_axaddr_0_reg),
                                               .desc_1_axaddr_1_reg(desc_1_axaddr_1_reg),
                                               .desc_1_axaddr_2_reg(desc_1_axaddr_2_reg),
                                               .desc_1_axaddr_3_reg(desc_1_axaddr_3_reg),
                                               .desc_1_axid_0_reg(desc_1_axid_0_reg),
                                               .desc_1_axid_1_reg(desc_1_axid_1_reg),
                                               .desc_1_axid_2_reg(desc_1_axid_2_reg),
                                               .desc_1_axid_3_reg(desc_1_axid_3_reg),
                                               .desc_1_axuser_0_reg(desc_1_axuser_0_reg),
                                               .desc_1_axuser_1_reg(desc_1_axuser_1_reg),
                                               .desc_1_axuser_2_reg(desc_1_axuser_2_reg),
                                               .desc_1_axuser_3_reg(desc_1_axuser_3_reg),
                                               .desc_1_axuser_4_reg(desc_1_axuser_4_reg),
                                               .desc_1_axuser_5_reg(desc_1_axuser_5_reg),
                                               .desc_1_axuser_6_reg(desc_1_axuser_6_reg),
                                               .desc_1_axuser_7_reg(desc_1_axuser_7_reg),
                                               .desc_1_axuser_8_reg(desc_1_axuser_8_reg),
                                               .desc_1_axuser_9_reg(desc_1_axuser_9_reg),
                                               .desc_1_axuser_10_reg(desc_1_axuser_10_reg),
                                               .desc_1_axuser_11_reg(desc_1_axuser_11_reg),
                                               .desc_1_axuser_12_reg(desc_1_axuser_12_reg),
                                               .desc_1_axuser_13_reg(desc_1_axuser_13_reg),
                                               .desc_1_axuser_14_reg(desc_1_axuser_14_reg),
                                               .desc_1_axuser_15_reg(desc_1_axuser_15_reg),
                                               .desc_1_xuser_0_reg(desc_1_xuser_0_reg),
                                               .desc_1_xuser_1_reg(desc_1_xuser_1_reg),
                                               .desc_1_xuser_2_reg(desc_1_xuser_2_reg),
                                               .desc_1_xuser_3_reg(desc_1_xuser_3_reg),
                                               .desc_1_xuser_4_reg(desc_1_xuser_4_reg),
                                               .desc_1_xuser_5_reg(desc_1_xuser_5_reg),
                                               .desc_1_xuser_6_reg(desc_1_xuser_6_reg),
                                               .desc_1_xuser_7_reg(desc_1_xuser_7_reg),
                                               .desc_1_xuser_8_reg(desc_1_xuser_8_reg),
                                               .desc_1_xuser_9_reg(desc_1_xuser_9_reg),
                                               .desc_1_xuser_10_reg(desc_1_xuser_10_reg),
                                               .desc_1_xuser_11_reg(desc_1_xuser_11_reg),
                                               .desc_1_xuser_12_reg(desc_1_xuser_12_reg),
                                               .desc_1_xuser_13_reg(desc_1_xuser_13_reg),
                                               .desc_1_xuser_14_reg(desc_1_xuser_14_reg),
                                               .desc_1_xuser_15_reg(desc_1_xuser_15_reg),
                                               .desc_1_wuser_0_reg(desc_1_wuser_0_reg),
                                               .desc_1_wuser_1_reg(desc_1_wuser_1_reg),
                                               .desc_1_wuser_2_reg(desc_1_wuser_2_reg),
                                               .desc_1_wuser_3_reg(desc_1_wuser_3_reg),
                                               .desc_1_wuser_4_reg(desc_1_wuser_4_reg),
                                               .desc_1_wuser_5_reg(desc_1_wuser_5_reg),
                                               .desc_1_wuser_6_reg(desc_1_wuser_6_reg),
                                               .desc_1_wuser_7_reg(desc_1_wuser_7_reg),
                                               .desc_1_wuser_8_reg(desc_1_wuser_8_reg),
                                               .desc_1_wuser_9_reg(desc_1_wuser_9_reg),
                                               .desc_1_wuser_10_reg(desc_1_wuser_10_reg),
                                               .desc_1_wuser_11_reg(desc_1_wuser_11_reg),
                                               .desc_1_wuser_12_reg(desc_1_wuser_12_reg),
                                               .desc_1_wuser_13_reg(desc_1_wuser_13_reg),
                                               .desc_1_wuser_14_reg(desc_1_wuser_14_reg),
                                               .desc_1_wuser_15_reg(desc_1_wuser_15_reg),
                                               .desc_2_txn_type_reg(desc_2_txn_type_reg),
                                               .desc_2_size_reg (desc_2_size_reg),
                                               .desc_2_data_offset_reg(desc_2_data_offset_reg),
                                               .desc_2_data_host_addr_0_reg(desc_2_data_host_addr_0_reg),
                                               .desc_2_data_host_addr_1_reg(desc_2_data_host_addr_1_reg),
                                               .desc_2_data_host_addr_2_reg(desc_2_data_host_addr_2_reg),
                                               .desc_2_data_host_addr_3_reg(desc_2_data_host_addr_3_reg),
                                               .desc_2_wstrb_host_addr_0_reg(desc_2_wstrb_host_addr_0_reg),
                                               .desc_2_wstrb_host_addr_1_reg(desc_2_wstrb_host_addr_1_reg),
                                               .desc_2_wstrb_host_addr_2_reg(desc_2_wstrb_host_addr_2_reg),
                                               .desc_2_wstrb_host_addr_3_reg(desc_2_wstrb_host_addr_3_reg),
                                               .desc_2_axsize_reg(desc_2_axsize_reg),
                                               .desc_2_attr_reg (desc_2_attr_reg),
                                               .desc_2_axaddr_0_reg(desc_2_axaddr_0_reg),
                                               .desc_2_axaddr_1_reg(desc_2_axaddr_1_reg),
                                               .desc_2_axaddr_2_reg(desc_2_axaddr_2_reg),
                                               .desc_2_axaddr_3_reg(desc_2_axaddr_3_reg),
                                               .desc_2_axid_0_reg(desc_2_axid_0_reg),
                                               .desc_2_axid_1_reg(desc_2_axid_1_reg),
                                               .desc_2_axid_2_reg(desc_2_axid_2_reg),
                                               .desc_2_axid_3_reg(desc_2_axid_3_reg),
                                               .desc_2_axuser_0_reg(desc_2_axuser_0_reg),
                                               .desc_2_axuser_1_reg(desc_2_axuser_1_reg),
                                               .desc_2_axuser_2_reg(desc_2_axuser_2_reg),
                                               .desc_2_axuser_3_reg(desc_2_axuser_3_reg),
                                               .desc_2_axuser_4_reg(desc_2_axuser_4_reg),
                                               .desc_2_axuser_5_reg(desc_2_axuser_5_reg),
                                               .desc_2_axuser_6_reg(desc_2_axuser_6_reg),
                                               .desc_2_axuser_7_reg(desc_2_axuser_7_reg),
                                               .desc_2_axuser_8_reg(desc_2_axuser_8_reg),
                                               .desc_2_axuser_9_reg(desc_2_axuser_9_reg),
                                               .desc_2_axuser_10_reg(desc_2_axuser_10_reg),
                                               .desc_2_axuser_11_reg(desc_2_axuser_11_reg),
                                               .desc_2_axuser_12_reg(desc_2_axuser_12_reg),
                                               .desc_2_axuser_13_reg(desc_2_axuser_13_reg),
                                               .desc_2_axuser_14_reg(desc_2_axuser_14_reg),
                                               .desc_2_axuser_15_reg(desc_2_axuser_15_reg),
                                               .desc_2_xuser_0_reg(desc_2_xuser_0_reg),
                                               .desc_2_xuser_1_reg(desc_2_xuser_1_reg),
                                               .desc_2_xuser_2_reg(desc_2_xuser_2_reg),
                                               .desc_2_xuser_3_reg(desc_2_xuser_3_reg),
                                               .desc_2_xuser_4_reg(desc_2_xuser_4_reg),
                                               .desc_2_xuser_5_reg(desc_2_xuser_5_reg),
                                               .desc_2_xuser_6_reg(desc_2_xuser_6_reg),
                                               .desc_2_xuser_7_reg(desc_2_xuser_7_reg),
                                               .desc_2_xuser_8_reg(desc_2_xuser_8_reg),
                                               .desc_2_xuser_9_reg(desc_2_xuser_9_reg),
                                               .desc_2_xuser_10_reg(desc_2_xuser_10_reg),
                                               .desc_2_xuser_11_reg(desc_2_xuser_11_reg),
                                               .desc_2_xuser_12_reg(desc_2_xuser_12_reg),
                                               .desc_2_xuser_13_reg(desc_2_xuser_13_reg),
                                               .desc_2_xuser_14_reg(desc_2_xuser_14_reg),
                                               .desc_2_xuser_15_reg(desc_2_xuser_15_reg),
                                               .desc_2_wuser_0_reg(desc_2_wuser_0_reg),
                                               .desc_2_wuser_1_reg(desc_2_wuser_1_reg),
                                               .desc_2_wuser_2_reg(desc_2_wuser_2_reg),
                                               .desc_2_wuser_3_reg(desc_2_wuser_3_reg),
                                               .desc_2_wuser_4_reg(desc_2_wuser_4_reg),
                                               .desc_2_wuser_5_reg(desc_2_wuser_5_reg),
                                               .desc_2_wuser_6_reg(desc_2_wuser_6_reg),
                                               .desc_2_wuser_7_reg(desc_2_wuser_7_reg),
                                               .desc_2_wuser_8_reg(desc_2_wuser_8_reg),
                                               .desc_2_wuser_9_reg(desc_2_wuser_9_reg),
                                               .desc_2_wuser_10_reg(desc_2_wuser_10_reg),
                                               .desc_2_wuser_11_reg(desc_2_wuser_11_reg),
                                               .desc_2_wuser_12_reg(desc_2_wuser_12_reg),
                                               .desc_2_wuser_13_reg(desc_2_wuser_13_reg),
                                               .desc_2_wuser_14_reg(desc_2_wuser_14_reg),
                                               .desc_2_wuser_15_reg(desc_2_wuser_15_reg),
                                               .desc_3_txn_type_reg(desc_3_txn_type_reg),
                                               .desc_3_size_reg (desc_3_size_reg),
                                               .desc_3_data_offset_reg(desc_3_data_offset_reg),
                                               .desc_3_data_host_addr_0_reg(desc_3_data_host_addr_0_reg),
                                               .desc_3_data_host_addr_1_reg(desc_3_data_host_addr_1_reg),
                                               .desc_3_data_host_addr_2_reg(desc_3_data_host_addr_2_reg),
                                               .desc_3_data_host_addr_3_reg(desc_3_data_host_addr_3_reg),
                                               .desc_3_wstrb_host_addr_0_reg(desc_3_wstrb_host_addr_0_reg),
                                               .desc_3_wstrb_host_addr_1_reg(desc_3_wstrb_host_addr_1_reg),
                                               .desc_3_wstrb_host_addr_2_reg(desc_3_wstrb_host_addr_2_reg),
                                               .desc_3_wstrb_host_addr_3_reg(desc_3_wstrb_host_addr_3_reg),
                                               .desc_3_axsize_reg(desc_3_axsize_reg),
                                               .desc_3_attr_reg (desc_3_attr_reg),
                                               .desc_3_axaddr_0_reg(desc_3_axaddr_0_reg),
                                               .desc_3_axaddr_1_reg(desc_3_axaddr_1_reg),
                                               .desc_3_axaddr_2_reg(desc_3_axaddr_2_reg),
                                               .desc_3_axaddr_3_reg(desc_3_axaddr_3_reg),
                                               .desc_3_axid_0_reg(desc_3_axid_0_reg),
                                               .desc_3_axid_1_reg(desc_3_axid_1_reg),
                                               .desc_3_axid_2_reg(desc_3_axid_2_reg),
                                               .desc_3_axid_3_reg(desc_3_axid_3_reg),
                                               .desc_3_axuser_0_reg(desc_3_axuser_0_reg),
                                               .desc_3_axuser_1_reg(desc_3_axuser_1_reg),
                                               .desc_3_axuser_2_reg(desc_3_axuser_2_reg),
                                               .desc_3_axuser_3_reg(desc_3_axuser_3_reg),
                                               .desc_3_axuser_4_reg(desc_3_axuser_4_reg),
                                               .desc_3_axuser_5_reg(desc_3_axuser_5_reg),
                                               .desc_3_axuser_6_reg(desc_3_axuser_6_reg),
                                               .desc_3_axuser_7_reg(desc_3_axuser_7_reg),
                                               .desc_3_axuser_8_reg(desc_3_axuser_8_reg),
                                               .desc_3_axuser_9_reg(desc_3_axuser_9_reg),
                                               .desc_3_axuser_10_reg(desc_3_axuser_10_reg),
                                               .desc_3_axuser_11_reg(desc_3_axuser_11_reg),
                                               .desc_3_axuser_12_reg(desc_3_axuser_12_reg),
                                               .desc_3_axuser_13_reg(desc_3_axuser_13_reg),
                                               .desc_3_axuser_14_reg(desc_3_axuser_14_reg),
                                               .desc_3_axuser_15_reg(desc_3_axuser_15_reg),
                                               .desc_3_xuser_0_reg(desc_3_xuser_0_reg),
                                               .desc_3_xuser_1_reg(desc_3_xuser_1_reg),
                                               .desc_3_xuser_2_reg(desc_3_xuser_2_reg),
                                               .desc_3_xuser_3_reg(desc_3_xuser_3_reg),
                                               .desc_3_xuser_4_reg(desc_3_xuser_4_reg),
                                               .desc_3_xuser_5_reg(desc_3_xuser_5_reg),
                                               .desc_3_xuser_6_reg(desc_3_xuser_6_reg),
                                               .desc_3_xuser_7_reg(desc_3_xuser_7_reg),
                                               .desc_3_xuser_8_reg(desc_3_xuser_8_reg),
                                               .desc_3_xuser_9_reg(desc_3_xuser_9_reg),
                                               .desc_3_xuser_10_reg(desc_3_xuser_10_reg),
                                               .desc_3_xuser_11_reg(desc_3_xuser_11_reg),
                                               .desc_3_xuser_12_reg(desc_3_xuser_12_reg),
                                               .desc_3_xuser_13_reg(desc_3_xuser_13_reg),
                                               .desc_3_xuser_14_reg(desc_3_xuser_14_reg),
                                               .desc_3_xuser_15_reg(desc_3_xuser_15_reg),
                                               .desc_3_wuser_0_reg(desc_3_wuser_0_reg),
                                               .desc_3_wuser_1_reg(desc_3_wuser_1_reg),
                                               .desc_3_wuser_2_reg(desc_3_wuser_2_reg),
                                               .desc_3_wuser_3_reg(desc_3_wuser_3_reg),
                                               .desc_3_wuser_4_reg(desc_3_wuser_4_reg),
                                               .desc_3_wuser_5_reg(desc_3_wuser_5_reg),
                                               .desc_3_wuser_6_reg(desc_3_wuser_6_reg),
                                               .desc_3_wuser_7_reg(desc_3_wuser_7_reg),
                                               .desc_3_wuser_8_reg(desc_3_wuser_8_reg),
                                               .desc_3_wuser_9_reg(desc_3_wuser_9_reg),
                                               .desc_3_wuser_10_reg(desc_3_wuser_10_reg),
                                               .desc_3_wuser_11_reg(desc_3_wuser_11_reg),
                                               .desc_3_wuser_12_reg(desc_3_wuser_12_reg),
                                               .desc_3_wuser_13_reg(desc_3_wuser_13_reg),
                                               .desc_3_wuser_14_reg(desc_3_wuser_14_reg),
                                               .desc_3_wuser_15_reg(desc_3_wuser_15_reg),
                                               .desc_4_txn_type_reg(desc_4_txn_type_reg),
                                               .desc_4_size_reg (desc_4_size_reg),
                                               .desc_4_data_offset_reg(desc_4_data_offset_reg),
                                               .desc_4_data_host_addr_0_reg(desc_4_data_host_addr_0_reg),
                                               .desc_4_data_host_addr_1_reg(desc_4_data_host_addr_1_reg),
                                               .desc_4_data_host_addr_2_reg(desc_4_data_host_addr_2_reg),
                                               .desc_4_data_host_addr_3_reg(desc_4_data_host_addr_3_reg),
                                               .desc_4_wstrb_host_addr_0_reg(desc_4_wstrb_host_addr_0_reg),
                                               .desc_4_wstrb_host_addr_1_reg(desc_4_wstrb_host_addr_1_reg),
                                               .desc_4_wstrb_host_addr_2_reg(desc_4_wstrb_host_addr_2_reg),
                                               .desc_4_wstrb_host_addr_3_reg(desc_4_wstrb_host_addr_3_reg),
                                               .desc_4_axsize_reg(desc_4_axsize_reg),
                                               .desc_4_attr_reg (desc_4_attr_reg),
                                               .desc_4_axaddr_0_reg(desc_4_axaddr_0_reg),
                                               .desc_4_axaddr_1_reg(desc_4_axaddr_1_reg),
                                               .desc_4_axaddr_2_reg(desc_4_axaddr_2_reg),
                                               .desc_4_axaddr_3_reg(desc_4_axaddr_3_reg),
                                               .desc_4_axid_0_reg(desc_4_axid_0_reg),
                                               .desc_4_axid_1_reg(desc_4_axid_1_reg),
                                               .desc_4_axid_2_reg(desc_4_axid_2_reg),
                                               .desc_4_axid_3_reg(desc_4_axid_3_reg),
                                               .desc_4_axuser_0_reg(desc_4_axuser_0_reg),
                                               .desc_4_axuser_1_reg(desc_4_axuser_1_reg),
                                               .desc_4_axuser_2_reg(desc_4_axuser_2_reg),
                                               .desc_4_axuser_3_reg(desc_4_axuser_3_reg),
                                               .desc_4_axuser_4_reg(desc_4_axuser_4_reg),
                                               .desc_4_axuser_5_reg(desc_4_axuser_5_reg),
                                               .desc_4_axuser_6_reg(desc_4_axuser_6_reg),
                                               .desc_4_axuser_7_reg(desc_4_axuser_7_reg),
                                               .desc_4_axuser_8_reg(desc_4_axuser_8_reg),
                                               .desc_4_axuser_9_reg(desc_4_axuser_9_reg),
                                               .desc_4_axuser_10_reg(desc_4_axuser_10_reg),
                                               .desc_4_axuser_11_reg(desc_4_axuser_11_reg),
                                               .desc_4_axuser_12_reg(desc_4_axuser_12_reg),
                                               .desc_4_axuser_13_reg(desc_4_axuser_13_reg),
                                               .desc_4_axuser_14_reg(desc_4_axuser_14_reg),
                                               .desc_4_axuser_15_reg(desc_4_axuser_15_reg),
                                               .desc_4_xuser_0_reg(desc_4_xuser_0_reg),
                                               .desc_4_xuser_1_reg(desc_4_xuser_1_reg),
                                               .desc_4_xuser_2_reg(desc_4_xuser_2_reg),
                                               .desc_4_xuser_3_reg(desc_4_xuser_3_reg),
                                               .desc_4_xuser_4_reg(desc_4_xuser_4_reg),
                                               .desc_4_xuser_5_reg(desc_4_xuser_5_reg),
                                               .desc_4_xuser_6_reg(desc_4_xuser_6_reg),
                                               .desc_4_xuser_7_reg(desc_4_xuser_7_reg),
                                               .desc_4_xuser_8_reg(desc_4_xuser_8_reg),
                                               .desc_4_xuser_9_reg(desc_4_xuser_9_reg),
                                               .desc_4_xuser_10_reg(desc_4_xuser_10_reg),
                                               .desc_4_xuser_11_reg(desc_4_xuser_11_reg),
                                               .desc_4_xuser_12_reg(desc_4_xuser_12_reg),
                                               .desc_4_xuser_13_reg(desc_4_xuser_13_reg),
                                               .desc_4_xuser_14_reg(desc_4_xuser_14_reg),
                                               .desc_4_xuser_15_reg(desc_4_xuser_15_reg),
                                               .desc_4_wuser_0_reg(desc_4_wuser_0_reg),
                                               .desc_4_wuser_1_reg(desc_4_wuser_1_reg),
                                               .desc_4_wuser_2_reg(desc_4_wuser_2_reg),
                                               .desc_4_wuser_3_reg(desc_4_wuser_3_reg),
                                               .desc_4_wuser_4_reg(desc_4_wuser_4_reg),
                                               .desc_4_wuser_5_reg(desc_4_wuser_5_reg),
                                               .desc_4_wuser_6_reg(desc_4_wuser_6_reg),
                                               .desc_4_wuser_7_reg(desc_4_wuser_7_reg),
                                               .desc_4_wuser_8_reg(desc_4_wuser_8_reg),
                                               .desc_4_wuser_9_reg(desc_4_wuser_9_reg),
                                               .desc_4_wuser_10_reg(desc_4_wuser_10_reg),
                                               .desc_4_wuser_11_reg(desc_4_wuser_11_reg),
                                               .desc_4_wuser_12_reg(desc_4_wuser_12_reg),
                                               .desc_4_wuser_13_reg(desc_4_wuser_13_reg),
                                               .desc_4_wuser_14_reg(desc_4_wuser_14_reg),
                                               .desc_4_wuser_15_reg(desc_4_wuser_15_reg),
                                               .desc_5_txn_type_reg(desc_5_txn_type_reg),
                                               .desc_5_size_reg (desc_5_size_reg),
                                               .desc_5_data_offset_reg(desc_5_data_offset_reg),
                                               .desc_5_data_host_addr_0_reg(desc_5_data_host_addr_0_reg),
                                               .desc_5_data_host_addr_1_reg(desc_5_data_host_addr_1_reg),
                                               .desc_5_data_host_addr_2_reg(desc_5_data_host_addr_2_reg),
                                               .desc_5_data_host_addr_3_reg(desc_5_data_host_addr_3_reg),
                                               .desc_5_wstrb_host_addr_0_reg(desc_5_wstrb_host_addr_0_reg),
                                               .desc_5_wstrb_host_addr_1_reg(desc_5_wstrb_host_addr_1_reg),
                                               .desc_5_wstrb_host_addr_2_reg(desc_5_wstrb_host_addr_2_reg),
                                               .desc_5_wstrb_host_addr_3_reg(desc_5_wstrb_host_addr_3_reg),
                                               .desc_5_axsize_reg(desc_5_axsize_reg),
                                               .desc_5_attr_reg (desc_5_attr_reg),
                                               .desc_5_axaddr_0_reg(desc_5_axaddr_0_reg),
                                               .desc_5_axaddr_1_reg(desc_5_axaddr_1_reg),
                                               .desc_5_axaddr_2_reg(desc_5_axaddr_2_reg),
                                               .desc_5_axaddr_3_reg(desc_5_axaddr_3_reg),
                                               .desc_5_axid_0_reg(desc_5_axid_0_reg),
                                               .desc_5_axid_1_reg(desc_5_axid_1_reg),
                                               .desc_5_axid_2_reg(desc_5_axid_2_reg),
                                               .desc_5_axid_3_reg(desc_5_axid_3_reg),
                                               .desc_5_axuser_0_reg(desc_5_axuser_0_reg),
                                               .desc_5_axuser_1_reg(desc_5_axuser_1_reg),
                                               .desc_5_axuser_2_reg(desc_5_axuser_2_reg),
                                               .desc_5_axuser_3_reg(desc_5_axuser_3_reg),
                                               .desc_5_axuser_4_reg(desc_5_axuser_4_reg),
                                               .desc_5_axuser_5_reg(desc_5_axuser_5_reg),
                                               .desc_5_axuser_6_reg(desc_5_axuser_6_reg),
                                               .desc_5_axuser_7_reg(desc_5_axuser_7_reg),
                                               .desc_5_axuser_8_reg(desc_5_axuser_8_reg),
                                               .desc_5_axuser_9_reg(desc_5_axuser_9_reg),
                                               .desc_5_axuser_10_reg(desc_5_axuser_10_reg),
                                               .desc_5_axuser_11_reg(desc_5_axuser_11_reg),
                                               .desc_5_axuser_12_reg(desc_5_axuser_12_reg),
                                               .desc_5_axuser_13_reg(desc_5_axuser_13_reg),
                                               .desc_5_axuser_14_reg(desc_5_axuser_14_reg),
                                               .desc_5_axuser_15_reg(desc_5_axuser_15_reg),
                                               .desc_5_xuser_0_reg(desc_5_xuser_0_reg),
                                               .desc_5_xuser_1_reg(desc_5_xuser_1_reg),
                                               .desc_5_xuser_2_reg(desc_5_xuser_2_reg),
                                               .desc_5_xuser_3_reg(desc_5_xuser_3_reg),
                                               .desc_5_xuser_4_reg(desc_5_xuser_4_reg),
                                               .desc_5_xuser_5_reg(desc_5_xuser_5_reg),
                                               .desc_5_xuser_6_reg(desc_5_xuser_6_reg),
                                               .desc_5_xuser_7_reg(desc_5_xuser_7_reg),
                                               .desc_5_xuser_8_reg(desc_5_xuser_8_reg),
                                               .desc_5_xuser_9_reg(desc_5_xuser_9_reg),
                                               .desc_5_xuser_10_reg(desc_5_xuser_10_reg),
                                               .desc_5_xuser_11_reg(desc_5_xuser_11_reg),
                                               .desc_5_xuser_12_reg(desc_5_xuser_12_reg),
                                               .desc_5_xuser_13_reg(desc_5_xuser_13_reg),
                                               .desc_5_xuser_14_reg(desc_5_xuser_14_reg),
                                               .desc_5_xuser_15_reg(desc_5_xuser_15_reg),
                                               .desc_5_wuser_0_reg(desc_5_wuser_0_reg),
                                               .desc_5_wuser_1_reg(desc_5_wuser_1_reg),
                                               .desc_5_wuser_2_reg(desc_5_wuser_2_reg),
                                               .desc_5_wuser_3_reg(desc_5_wuser_3_reg),
                                               .desc_5_wuser_4_reg(desc_5_wuser_4_reg),
                                               .desc_5_wuser_5_reg(desc_5_wuser_5_reg),
                                               .desc_5_wuser_6_reg(desc_5_wuser_6_reg),
                                               .desc_5_wuser_7_reg(desc_5_wuser_7_reg),
                                               .desc_5_wuser_8_reg(desc_5_wuser_8_reg),
                                               .desc_5_wuser_9_reg(desc_5_wuser_9_reg),
                                               .desc_5_wuser_10_reg(desc_5_wuser_10_reg),
                                               .desc_5_wuser_11_reg(desc_5_wuser_11_reg),
                                               .desc_5_wuser_12_reg(desc_5_wuser_12_reg),
                                               .desc_5_wuser_13_reg(desc_5_wuser_13_reg),
                                               .desc_5_wuser_14_reg(desc_5_wuser_14_reg),
                                               .desc_5_wuser_15_reg(desc_5_wuser_15_reg),
                                               .desc_6_txn_type_reg(desc_6_txn_type_reg),
                                               .desc_6_size_reg (desc_6_size_reg),
                                               .desc_6_data_offset_reg(desc_6_data_offset_reg),
                                               .desc_6_data_host_addr_0_reg(desc_6_data_host_addr_0_reg),
                                               .desc_6_data_host_addr_1_reg(desc_6_data_host_addr_1_reg),
                                               .desc_6_data_host_addr_2_reg(desc_6_data_host_addr_2_reg),
                                               .desc_6_data_host_addr_3_reg(desc_6_data_host_addr_3_reg),
                                               .desc_6_wstrb_host_addr_0_reg(desc_6_wstrb_host_addr_0_reg),
                                               .desc_6_wstrb_host_addr_1_reg(desc_6_wstrb_host_addr_1_reg),
                                               .desc_6_wstrb_host_addr_2_reg(desc_6_wstrb_host_addr_2_reg),
                                               .desc_6_wstrb_host_addr_3_reg(desc_6_wstrb_host_addr_3_reg),
                                               .desc_6_axsize_reg(desc_6_axsize_reg),
                                               .desc_6_attr_reg (desc_6_attr_reg),
                                               .desc_6_axaddr_0_reg(desc_6_axaddr_0_reg),
                                               .desc_6_axaddr_1_reg(desc_6_axaddr_1_reg),
                                               .desc_6_axaddr_2_reg(desc_6_axaddr_2_reg),
                                               .desc_6_axaddr_3_reg(desc_6_axaddr_3_reg),
                                               .desc_6_axid_0_reg(desc_6_axid_0_reg),
                                               .desc_6_axid_1_reg(desc_6_axid_1_reg),
                                               .desc_6_axid_2_reg(desc_6_axid_2_reg),
                                               .desc_6_axid_3_reg(desc_6_axid_3_reg),
                                               .desc_6_axuser_0_reg(desc_6_axuser_0_reg),
                                               .desc_6_axuser_1_reg(desc_6_axuser_1_reg),
                                               .desc_6_axuser_2_reg(desc_6_axuser_2_reg),
                                               .desc_6_axuser_3_reg(desc_6_axuser_3_reg),
                                               .desc_6_axuser_4_reg(desc_6_axuser_4_reg),
                                               .desc_6_axuser_5_reg(desc_6_axuser_5_reg),
                                               .desc_6_axuser_6_reg(desc_6_axuser_6_reg),
                                               .desc_6_axuser_7_reg(desc_6_axuser_7_reg),
                                               .desc_6_axuser_8_reg(desc_6_axuser_8_reg),
                                               .desc_6_axuser_9_reg(desc_6_axuser_9_reg),
                                               .desc_6_axuser_10_reg(desc_6_axuser_10_reg),
                                               .desc_6_axuser_11_reg(desc_6_axuser_11_reg),
                                               .desc_6_axuser_12_reg(desc_6_axuser_12_reg),
                                               .desc_6_axuser_13_reg(desc_6_axuser_13_reg),
                                               .desc_6_axuser_14_reg(desc_6_axuser_14_reg),
                                               .desc_6_axuser_15_reg(desc_6_axuser_15_reg),
                                               .desc_6_xuser_0_reg(desc_6_xuser_0_reg),
                                               .desc_6_xuser_1_reg(desc_6_xuser_1_reg),
                                               .desc_6_xuser_2_reg(desc_6_xuser_2_reg),
                                               .desc_6_xuser_3_reg(desc_6_xuser_3_reg),
                                               .desc_6_xuser_4_reg(desc_6_xuser_4_reg),
                                               .desc_6_xuser_5_reg(desc_6_xuser_5_reg),
                                               .desc_6_xuser_6_reg(desc_6_xuser_6_reg),
                                               .desc_6_xuser_7_reg(desc_6_xuser_7_reg),
                                               .desc_6_xuser_8_reg(desc_6_xuser_8_reg),
                                               .desc_6_xuser_9_reg(desc_6_xuser_9_reg),
                                               .desc_6_xuser_10_reg(desc_6_xuser_10_reg),
                                               .desc_6_xuser_11_reg(desc_6_xuser_11_reg),
                                               .desc_6_xuser_12_reg(desc_6_xuser_12_reg),
                                               .desc_6_xuser_13_reg(desc_6_xuser_13_reg),
                                               .desc_6_xuser_14_reg(desc_6_xuser_14_reg),
                                               .desc_6_xuser_15_reg(desc_6_xuser_15_reg),
                                               .desc_6_wuser_0_reg(desc_6_wuser_0_reg),
                                               .desc_6_wuser_1_reg(desc_6_wuser_1_reg),
                                               .desc_6_wuser_2_reg(desc_6_wuser_2_reg),
                                               .desc_6_wuser_3_reg(desc_6_wuser_3_reg),
                                               .desc_6_wuser_4_reg(desc_6_wuser_4_reg),
                                               .desc_6_wuser_5_reg(desc_6_wuser_5_reg),
                                               .desc_6_wuser_6_reg(desc_6_wuser_6_reg),
                                               .desc_6_wuser_7_reg(desc_6_wuser_7_reg),
                                               .desc_6_wuser_8_reg(desc_6_wuser_8_reg),
                                               .desc_6_wuser_9_reg(desc_6_wuser_9_reg),
                                               .desc_6_wuser_10_reg(desc_6_wuser_10_reg),
                                               .desc_6_wuser_11_reg(desc_6_wuser_11_reg),
                                               .desc_6_wuser_12_reg(desc_6_wuser_12_reg),
                                               .desc_6_wuser_13_reg(desc_6_wuser_13_reg),
                                               .desc_6_wuser_14_reg(desc_6_wuser_14_reg),
                                               .desc_6_wuser_15_reg(desc_6_wuser_15_reg),
                                               .desc_7_txn_type_reg(desc_7_txn_type_reg),
                                               .desc_7_size_reg (desc_7_size_reg),
                                               .desc_7_data_offset_reg(desc_7_data_offset_reg),
                                               .desc_7_data_host_addr_0_reg(desc_7_data_host_addr_0_reg),
                                               .desc_7_data_host_addr_1_reg(desc_7_data_host_addr_1_reg),
                                               .desc_7_data_host_addr_2_reg(desc_7_data_host_addr_2_reg),
                                               .desc_7_data_host_addr_3_reg(desc_7_data_host_addr_3_reg),
                                               .desc_7_wstrb_host_addr_0_reg(desc_7_wstrb_host_addr_0_reg),
                                               .desc_7_wstrb_host_addr_1_reg(desc_7_wstrb_host_addr_1_reg),
                                               .desc_7_wstrb_host_addr_2_reg(desc_7_wstrb_host_addr_2_reg),
                                               .desc_7_wstrb_host_addr_3_reg(desc_7_wstrb_host_addr_3_reg),
                                               .desc_7_axsize_reg(desc_7_axsize_reg),
                                               .desc_7_attr_reg (desc_7_attr_reg),
                                               .desc_7_axaddr_0_reg(desc_7_axaddr_0_reg),
                                               .desc_7_axaddr_1_reg(desc_7_axaddr_1_reg),
                                               .desc_7_axaddr_2_reg(desc_7_axaddr_2_reg),
                                               .desc_7_axaddr_3_reg(desc_7_axaddr_3_reg),
                                               .desc_7_axid_0_reg(desc_7_axid_0_reg),
                                               .desc_7_axid_1_reg(desc_7_axid_1_reg),
                                               .desc_7_axid_2_reg(desc_7_axid_2_reg),
                                               .desc_7_axid_3_reg(desc_7_axid_3_reg),
                                               .desc_7_axuser_0_reg(desc_7_axuser_0_reg),
                                               .desc_7_axuser_1_reg(desc_7_axuser_1_reg),
                                               .desc_7_axuser_2_reg(desc_7_axuser_2_reg),
                                               .desc_7_axuser_3_reg(desc_7_axuser_3_reg),
                                               .desc_7_axuser_4_reg(desc_7_axuser_4_reg),
                                               .desc_7_axuser_5_reg(desc_7_axuser_5_reg),
                                               .desc_7_axuser_6_reg(desc_7_axuser_6_reg),
                                               .desc_7_axuser_7_reg(desc_7_axuser_7_reg),
                                               .desc_7_axuser_8_reg(desc_7_axuser_8_reg),
                                               .desc_7_axuser_9_reg(desc_7_axuser_9_reg),
                                               .desc_7_axuser_10_reg(desc_7_axuser_10_reg),
                                               .desc_7_axuser_11_reg(desc_7_axuser_11_reg),
                                               .desc_7_axuser_12_reg(desc_7_axuser_12_reg),
                                               .desc_7_axuser_13_reg(desc_7_axuser_13_reg),
                                               .desc_7_axuser_14_reg(desc_7_axuser_14_reg),
                                               .desc_7_axuser_15_reg(desc_7_axuser_15_reg),
                                               .desc_7_xuser_0_reg(desc_7_xuser_0_reg),
                                               .desc_7_xuser_1_reg(desc_7_xuser_1_reg),
                                               .desc_7_xuser_2_reg(desc_7_xuser_2_reg),
                                               .desc_7_xuser_3_reg(desc_7_xuser_3_reg),
                                               .desc_7_xuser_4_reg(desc_7_xuser_4_reg),
                                               .desc_7_xuser_5_reg(desc_7_xuser_5_reg),
                                               .desc_7_xuser_6_reg(desc_7_xuser_6_reg),
                                               .desc_7_xuser_7_reg(desc_7_xuser_7_reg),
                                               .desc_7_xuser_8_reg(desc_7_xuser_8_reg),
                                               .desc_7_xuser_9_reg(desc_7_xuser_9_reg),
                                               .desc_7_xuser_10_reg(desc_7_xuser_10_reg),
                                               .desc_7_xuser_11_reg(desc_7_xuser_11_reg),
                                               .desc_7_xuser_12_reg(desc_7_xuser_12_reg),
                                               .desc_7_xuser_13_reg(desc_7_xuser_13_reg),
                                               .desc_7_xuser_14_reg(desc_7_xuser_14_reg),
                                               .desc_7_xuser_15_reg(desc_7_xuser_15_reg),
                                               .desc_7_wuser_0_reg(desc_7_wuser_0_reg),
                                               .desc_7_wuser_1_reg(desc_7_wuser_1_reg),
                                               .desc_7_wuser_2_reg(desc_7_wuser_2_reg),
                                               .desc_7_wuser_3_reg(desc_7_wuser_3_reg),
                                               .desc_7_wuser_4_reg(desc_7_wuser_4_reg),
                                               .desc_7_wuser_5_reg(desc_7_wuser_5_reg),
                                               .desc_7_wuser_6_reg(desc_7_wuser_6_reg),
                                               .desc_7_wuser_7_reg(desc_7_wuser_7_reg),
                                               .desc_7_wuser_8_reg(desc_7_wuser_8_reg),
                                               .desc_7_wuser_9_reg(desc_7_wuser_9_reg),
                                               .desc_7_wuser_10_reg(desc_7_wuser_10_reg),
                                               .desc_7_wuser_11_reg(desc_7_wuser_11_reg),
                                               .desc_7_wuser_12_reg(desc_7_wuser_12_reg),
                                               .desc_7_wuser_13_reg(desc_7_wuser_13_reg),
                                               .desc_7_wuser_14_reg(desc_7_wuser_14_reg),
                                               .desc_7_wuser_15_reg(desc_7_wuser_15_reg),
                                               .desc_8_txn_type_reg(desc_8_txn_type_reg),
                                               .desc_8_size_reg (desc_8_size_reg),
                                               .desc_8_data_offset_reg(desc_8_data_offset_reg),
                                               .desc_8_data_host_addr_0_reg(desc_8_data_host_addr_0_reg),
                                               .desc_8_data_host_addr_1_reg(desc_8_data_host_addr_1_reg),
                                               .desc_8_data_host_addr_2_reg(desc_8_data_host_addr_2_reg),
                                               .desc_8_data_host_addr_3_reg(desc_8_data_host_addr_3_reg),
                                               .desc_8_wstrb_host_addr_0_reg(desc_8_wstrb_host_addr_0_reg),
                                               .desc_8_wstrb_host_addr_1_reg(desc_8_wstrb_host_addr_1_reg),
                                               .desc_8_wstrb_host_addr_2_reg(desc_8_wstrb_host_addr_2_reg),
                                               .desc_8_wstrb_host_addr_3_reg(desc_8_wstrb_host_addr_3_reg),
                                               .desc_8_axsize_reg(desc_8_axsize_reg),
                                               .desc_8_attr_reg (desc_8_attr_reg),
                                               .desc_8_axaddr_0_reg(desc_8_axaddr_0_reg),
                                               .desc_8_axaddr_1_reg(desc_8_axaddr_1_reg),
                                               .desc_8_axaddr_2_reg(desc_8_axaddr_2_reg),
                                               .desc_8_axaddr_3_reg(desc_8_axaddr_3_reg),
                                               .desc_8_axid_0_reg(desc_8_axid_0_reg),
                                               .desc_8_axid_1_reg(desc_8_axid_1_reg),
                                               .desc_8_axid_2_reg(desc_8_axid_2_reg),
                                               .desc_8_axid_3_reg(desc_8_axid_3_reg),
                                               .desc_8_axuser_0_reg(desc_8_axuser_0_reg),
                                               .desc_8_axuser_1_reg(desc_8_axuser_1_reg),
                                               .desc_8_axuser_2_reg(desc_8_axuser_2_reg),
                                               .desc_8_axuser_3_reg(desc_8_axuser_3_reg),
                                               .desc_8_axuser_4_reg(desc_8_axuser_4_reg),
                                               .desc_8_axuser_5_reg(desc_8_axuser_5_reg),
                                               .desc_8_axuser_6_reg(desc_8_axuser_6_reg),
                                               .desc_8_axuser_7_reg(desc_8_axuser_7_reg),
                                               .desc_8_axuser_8_reg(desc_8_axuser_8_reg),
                                               .desc_8_axuser_9_reg(desc_8_axuser_9_reg),
                                               .desc_8_axuser_10_reg(desc_8_axuser_10_reg),
                                               .desc_8_axuser_11_reg(desc_8_axuser_11_reg),
                                               .desc_8_axuser_12_reg(desc_8_axuser_12_reg),
                                               .desc_8_axuser_13_reg(desc_8_axuser_13_reg),
                                               .desc_8_axuser_14_reg(desc_8_axuser_14_reg),
                                               .desc_8_axuser_15_reg(desc_8_axuser_15_reg),
                                               .desc_8_xuser_0_reg(desc_8_xuser_0_reg),
                                               .desc_8_xuser_1_reg(desc_8_xuser_1_reg),
                                               .desc_8_xuser_2_reg(desc_8_xuser_2_reg),
                                               .desc_8_xuser_3_reg(desc_8_xuser_3_reg),
                                               .desc_8_xuser_4_reg(desc_8_xuser_4_reg),
                                               .desc_8_xuser_5_reg(desc_8_xuser_5_reg),
                                               .desc_8_xuser_6_reg(desc_8_xuser_6_reg),
                                               .desc_8_xuser_7_reg(desc_8_xuser_7_reg),
                                               .desc_8_xuser_8_reg(desc_8_xuser_8_reg),
                                               .desc_8_xuser_9_reg(desc_8_xuser_9_reg),
                                               .desc_8_xuser_10_reg(desc_8_xuser_10_reg),
                                               .desc_8_xuser_11_reg(desc_8_xuser_11_reg),
                                               .desc_8_xuser_12_reg(desc_8_xuser_12_reg),
                                               .desc_8_xuser_13_reg(desc_8_xuser_13_reg),
                                               .desc_8_xuser_14_reg(desc_8_xuser_14_reg),
                                               .desc_8_xuser_15_reg(desc_8_xuser_15_reg),
                                               .desc_8_wuser_0_reg(desc_8_wuser_0_reg),
                                               .desc_8_wuser_1_reg(desc_8_wuser_1_reg),
                                               .desc_8_wuser_2_reg(desc_8_wuser_2_reg),
                                               .desc_8_wuser_3_reg(desc_8_wuser_3_reg),
                                               .desc_8_wuser_4_reg(desc_8_wuser_4_reg),
                                               .desc_8_wuser_5_reg(desc_8_wuser_5_reg),
                                               .desc_8_wuser_6_reg(desc_8_wuser_6_reg),
                                               .desc_8_wuser_7_reg(desc_8_wuser_7_reg),
                                               .desc_8_wuser_8_reg(desc_8_wuser_8_reg),
                                               .desc_8_wuser_9_reg(desc_8_wuser_9_reg),
                                               .desc_8_wuser_10_reg(desc_8_wuser_10_reg),
                                               .desc_8_wuser_11_reg(desc_8_wuser_11_reg),
                                               .desc_8_wuser_12_reg(desc_8_wuser_12_reg),
                                               .desc_8_wuser_13_reg(desc_8_wuser_13_reg),
                                               .desc_8_wuser_14_reg(desc_8_wuser_14_reg),
                                               .desc_8_wuser_15_reg(desc_8_wuser_15_reg),
                                               .desc_9_txn_type_reg(desc_9_txn_type_reg),
                                               .desc_9_size_reg (desc_9_size_reg),
                                               .desc_9_data_offset_reg(desc_9_data_offset_reg),
                                               .desc_9_data_host_addr_0_reg(desc_9_data_host_addr_0_reg),
                                               .desc_9_data_host_addr_1_reg(desc_9_data_host_addr_1_reg),
                                               .desc_9_data_host_addr_2_reg(desc_9_data_host_addr_2_reg),
                                               .desc_9_data_host_addr_3_reg(desc_9_data_host_addr_3_reg),
                                               .desc_9_wstrb_host_addr_0_reg(desc_9_wstrb_host_addr_0_reg),
                                               .desc_9_wstrb_host_addr_1_reg(desc_9_wstrb_host_addr_1_reg),
                                               .desc_9_wstrb_host_addr_2_reg(desc_9_wstrb_host_addr_2_reg),
                                               .desc_9_wstrb_host_addr_3_reg(desc_9_wstrb_host_addr_3_reg),
                                               .desc_9_axsize_reg(desc_9_axsize_reg),
                                               .desc_9_attr_reg (desc_9_attr_reg),
                                               .desc_9_axaddr_0_reg(desc_9_axaddr_0_reg),
                                               .desc_9_axaddr_1_reg(desc_9_axaddr_1_reg),
                                               .desc_9_axaddr_2_reg(desc_9_axaddr_2_reg),
                                               .desc_9_axaddr_3_reg(desc_9_axaddr_3_reg),
                                               .desc_9_axid_0_reg(desc_9_axid_0_reg),
                                               .desc_9_axid_1_reg(desc_9_axid_1_reg),
                                               .desc_9_axid_2_reg(desc_9_axid_2_reg),
                                               .desc_9_axid_3_reg(desc_9_axid_3_reg),
                                               .desc_9_axuser_0_reg(desc_9_axuser_0_reg),
                                               .desc_9_axuser_1_reg(desc_9_axuser_1_reg),
                                               .desc_9_axuser_2_reg(desc_9_axuser_2_reg),
                                               .desc_9_axuser_3_reg(desc_9_axuser_3_reg),
                                               .desc_9_axuser_4_reg(desc_9_axuser_4_reg),
                                               .desc_9_axuser_5_reg(desc_9_axuser_5_reg),
                                               .desc_9_axuser_6_reg(desc_9_axuser_6_reg),
                                               .desc_9_axuser_7_reg(desc_9_axuser_7_reg),
                                               .desc_9_axuser_8_reg(desc_9_axuser_8_reg),
                                               .desc_9_axuser_9_reg(desc_9_axuser_9_reg),
                                               .desc_9_axuser_10_reg(desc_9_axuser_10_reg),
                                               .desc_9_axuser_11_reg(desc_9_axuser_11_reg),
                                               .desc_9_axuser_12_reg(desc_9_axuser_12_reg),
                                               .desc_9_axuser_13_reg(desc_9_axuser_13_reg),
                                               .desc_9_axuser_14_reg(desc_9_axuser_14_reg),
                                               .desc_9_axuser_15_reg(desc_9_axuser_15_reg),
                                               .desc_9_xuser_0_reg(desc_9_xuser_0_reg),
                                               .desc_9_xuser_1_reg(desc_9_xuser_1_reg),
                                               .desc_9_xuser_2_reg(desc_9_xuser_2_reg),
                                               .desc_9_xuser_3_reg(desc_9_xuser_3_reg),
                                               .desc_9_xuser_4_reg(desc_9_xuser_4_reg),
                                               .desc_9_xuser_5_reg(desc_9_xuser_5_reg),
                                               .desc_9_xuser_6_reg(desc_9_xuser_6_reg),
                                               .desc_9_xuser_7_reg(desc_9_xuser_7_reg),
                                               .desc_9_xuser_8_reg(desc_9_xuser_8_reg),
                                               .desc_9_xuser_9_reg(desc_9_xuser_9_reg),
                                               .desc_9_xuser_10_reg(desc_9_xuser_10_reg),
                                               .desc_9_xuser_11_reg(desc_9_xuser_11_reg),
                                               .desc_9_xuser_12_reg(desc_9_xuser_12_reg),
                                               .desc_9_xuser_13_reg(desc_9_xuser_13_reg),
                                               .desc_9_xuser_14_reg(desc_9_xuser_14_reg),
                                               .desc_9_xuser_15_reg(desc_9_xuser_15_reg),
                                               .desc_9_wuser_0_reg(desc_9_wuser_0_reg),
                                               .desc_9_wuser_1_reg(desc_9_wuser_1_reg),
                                               .desc_9_wuser_2_reg(desc_9_wuser_2_reg),
                                               .desc_9_wuser_3_reg(desc_9_wuser_3_reg),
                                               .desc_9_wuser_4_reg(desc_9_wuser_4_reg),
                                               .desc_9_wuser_5_reg(desc_9_wuser_5_reg),
                                               .desc_9_wuser_6_reg(desc_9_wuser_6_reg),
                                               .desc_9_wuser_7_reg(desc_9_wuser_7_reg),
                                               .desc_9_wuser_8_reg(desc_9_wuser_8_reg),
                                               .desc_9_wuser_9_reg(desc_9_wuser_9_reg),
                                               .desc_9_wuser_10_reg(desc_9_wuser_10_reg),
                                               .desc_9_wuser_11_reg(desc_9_wuser_11_reg),
                                               .desc_9_wuser_12_reg(desc_9_wuser_12_reg),
                                               .desc_9_wuser_13_reg(desc_9_wuser_13_reg),
                                               .desc_9_wuser_14_reg(desc_9_wuser_14_reg),
                                               .desc_9_wuser_15_reg(desc_9_wuser_15_reg),
                                               .desc_10_txn_type_reg(desc_10_txn_type_reg),
                                               .desc_10_size_reg(desc_10_size_reg),
                                               .desc_10_data_offset_reg(desc_10_data_offset_reg),
                                               .desc_10_data_host_addr_0_reg(desc_10_data_host_addr_0_reg),
                                               .desc_10_data_host_addr_1_reg(desc_10_data_host_addr_1_reg),
                                               .desc_10_data_host_addr_2_reg(desc_10_data_host_addr_2_reg),
                                               .desc_10_data_host_addr_3_reg(desc_10_data_host_addr_3_reg),
                                               .desc_10_wstrb_host_addr_0_reg(desc_10_wstrb_host_addr_0_reg),
                                               .desc_10_wstrb_host_addr_1_reg(desc_10_wstrb_host_addr_1_reg),
                                               .desc_10_wstrb_host_addr_2_reg(desc_10_wstrb_host_addr_2_reg),
                                               .desc_10_wstrb_host_addr_3_reg(desc_10_wstrb_host_addr_3_reg),
                                               .desc_10_axsize_reg(desc_10_axsize_reg),
                                               .desc_10_attr_reg(desc_10_attr_reg),
                                               .desc_10_axaddr_0_reg(desc_10_axaddr_0_reg),
                                               .desc_10_axaddr_1_reg(desc_10_axaddr_1_reg),
                                               .desc_10_axaddr_2_reg(desc_10_axaddr_2_reg),
                                               .desc_10_axaddr_3_reg(desc_10_axaddr_3_reg),
                                               .desc_10_axid_0_reg(desc_10_axid_0_reg),
                                               .desc_10_axid_1_reg(desc_10_axid_1_reg),
                                               .desc_10_axid_2_reg(desc_10_axid_2_reg),
                                               .desc_10_axid_3_reg(desc_10_axid_3_reg),
                                               .desc_10_axuser_0_reg(desc_10_axuser_0_reg),
                                               .desc_10_axuser_1_reg(desc_10_axuser_1_reg),
                                               .desc_10_axuser_2_reg(desc_10_axuser_2_reg),
                                               .desc_10_axuser_3_reg(desc_10_axuser_3_reg),
                                               .desc_10_axuser_4_reg(desc_10_axuser_4_reg),
                                               .desc_10_axuser_5_reg(desc_10_axuser_5_reg),
                                               .desc_10_axuser_6_reg(desc_10_axuser_6_reg),
                                               .desc_10_axuser_7_reg(desc_10_axuser_7_reg),
                                               .desc_10_axuser_8_reg(desc_10_axuser_8_reg),
                                               .desc_10_axuser_9_reg(desc_10_axuser_9_reg),
                                               .desc_10_axuser_10_reg(desc_10_axuser_10_reg),
                                               .desc_10_axuser_11_reg(desc_10_axuser_11_reg),
                                               .desc_10_axuser_12_reg(desc_10_axuser_12_reg),
                                               .desc_10_axuser_13_reg(desc_10_axuser_13_reg),
                                               .desc_10_axuser_14_reg(desc_10_axuser_14_reg),
                                               .desc_10_axuser_15_reg(desc_10_axuser_15_reg),
                                               .desc_10_xuser_0_reg(desc_10_xuser_0_reg),
                                               .desc_10_xuser_1_reg(desc_10_xuser_1_reg),
                                               .desc_10_xuser_2_reg(desc_10_xuser_2_reg),
                                               .desc_10_xuser_3_reg(desc_10_xuser_3_reg),
                                               .desc_10_xuser_4_reg(desc_10_xuser_4_reg),
                                               .desc_10_xuser_5_reg(desc_10_xuser_5_reg),
                                               .desc_10_xuser_6_reg(desc_10_xuser_6_reg),
                                               .desc_10_xuser_7_reg(desc_10_xuser_7_reg),
                                               .desc_10_xuser_8_reg(desc_10_xuser_8_reg),
                                               .desc_10_xuser_9_reg(desc_10_xuser_9_reg),
                                               .desc_10_xuser_10_reg(desc_10_xuser_10_reg),
                                               .desc_10_xuser_11_reg(desc_10_xuser_11_reg),
                                               .desc_10_xuser_12_reg(desc_10_xuser_12_reg),
                                               .desc_10_xuser_13_reg(desc_10_xuser_13_reg),
                                               .desc_10_xuser_14_reg(desc_10_xuser_14_reg),
                                               .desc_10_xuser_15_reg(desc_10_xuser_15_reg),
                                               .desc_10_wuser_0_reg(desc_10_wuser_0_reg),
                                               .desc_10_wuser_1_reg(desc_10_wuser_1_reg),
                                               .desc_10_wuser_2_reg(desc_10_wuser_2_reg),
                                               .desc_10_wuser_3_reg(desc_10_wuser_3_reg),
                                               .desc_10_wuser_4_reg(desc_10_wuser_4_reg),
                                               .desc_10_wuser_5_reg(desc_10_wuser_5_reg),
                                               .desc_10_wuser_6_reg(desc_10_wuser_6_reg),
                                               .desc_10_wuser_7_reg(desc_10_wuser_7_reg),
                                               .desc_10_wuser_8_reg(desc_10_wuser_8_reg),
                                               .desc_10_wuser_9_reg(desc_10_wuser_9_reg),
                                               .desc_10_wuser_10_reg(desc_10_wuser_10_reg),
                                               .desc_10_wuser_11_reg(desc_10_wuser_11_reg),
                                               .desc_10_wuser_12_reg(desc_10_wuser_12_reg),
                                               .desc_10_wuser_13_reg(desc_10_wuser_13_reg),
                                               .desc_10_wuser_14_reg(desc_10_wuser_14_reg),
                                               .desc_10_wuser_15_reg(desc_10_wuser_15_reg),
                                               .desc_11_txn_type_reg(desc_11_txn_type_reg),
                                               .desc_11_size_reg(desc_11_size_reg),
                                               .desc_11_data_offset_reg(desc_11_data_offset_reg),
                                               .desc_11_data_host_addr_0_reg(desc_11_data_host_addr_0_reg),
                                               .desc_11_data_host_addr_1_reg(desc_11_data_host_addr_1_reg),
                                               .desc_11_data_host_addr_2_reg(desc_11_data_host_addr_2_reg),
                                               .desc_11_data_host_addr_3_reg(desc_11_data_host_addr_3_reg),
                                               .desc_11_wstrb_host_addr_0_reg(desc_11_wstrb_host_addr_0_reg),
                                               .desc_11_wstrb_host_addr_1_reg(desc_11_wstrb_host_addr_1_reg),
                                               .desc_11_wstrb_host_addr_2_reg(desc_11_wstrb_host_addr_2_reg),
                                               .desc_11_wstrb_host_addr_3_reg(desc_11_wstrb_host_addr_3_reg),
                                               .desc_11_axsize_reg(desc_11_axsize_reg),
                                               .desc_11_attr_reg(desc_11_attr_reg),
                                               .desc_11_axaddr_0_reg(desc_11_axaddr_0_reg),
                                               .desc_11_axaddr_1_reg(desc_11_axaddr_1_reg),
                                               .desc_11_axaddr_2_reg(desc_11_axaddr_2_reg),
                                               .desc_11_axaddr_3_reg(desc_11_axaddr_3_reg),
                                               .desc_11_axid_0_reg(desc_11_axid_0_reg),
                                               .desc_11_axid_1_reg(desc_11_axid_1_reg),
                                               .desc_11_axid_2_reg(desc_11_axid_2_reg),
                                               .desc_11_axid_3_reg(desc_11_axid_3_reg),
                                               .desc_11_axuser_0_reg(desc_11_axuser_0_reg),
                                               .desc_11_axuser_1_reg(desc_11_axuser_1_reg),
                                               .desc_11_axuser_2_reg(desc_11_axuser_2_reg),
                                               .desc_11_axuser_3_reg(desc_11_axuser_3_reg),
                                               .desc_11_axuser_4_reg(desc_11_axuser_4_reg),
                                               .desc_11_axuser_5_reg(desc_11_axuser_5_reg),
                                               .desc_11_axuser_6_reg(desc_11_axuser_6_reg),
                                               .desc_11_axuser_7_reg(desc_11_axuser_7_reg),
                                               .desc_11_axuser_8_reg(desc_11_axuser_8_reg),
                                               .desc_11_axuser_9_reg(desc_11_axuser_9_reg),
                                               .desc_11_axuser_10_reg(desc_11_axuser_10_reg),
                                               .desc_11_axuser_11_reg(desc_11_axuser_11_reg),
                                               .desc_11_axuser_12_reg(desc_11_axuser_12_reg),
                                               .desc_11_axuser_13_reg(desc_11_axuser_13_reg),
                                               .desc_11_axuser_14_reg(desc_11_axuser_14_reg),
                                               .desc_11_axuser_15_reg(desc_11_axuser_15_reg),
                                               .desc_11_xuser_0_reg(desc_11_xuser_0_reg),
                                               .desc_11_xuser_1_reg(desc_11_xuser_1_reg),
                                               .desc_11_xuser_2_reg(desc_11_xuser_2_reg),
                                               .desc_11_xuser_3_reg(desc_11_xuser_3_reg),
                                               .desc_11_xuser_4_reg(desc_11_xuser_4_reg),
                                               .desc_11_xuser_5_reg(desc_11_xuser_5_reg),
                                               .desc_11_xuser_6_reg(desc_11_xuser_6_reg),
                                               .desc_11_xuser_7_reg(desc_11_xuser_7_reg),
                                               .desc_11_xuser_8_reg(desc_11_xuser_8_reg),
                                               .desc_11_xuser_9_reg(desc_11_xuser_9_reg),
                                               .desc_11_xuser_10_reg(desc_11_xuser_10_reg),
                                               .desc_11_xuser_11_reg(desc_11_xuser_11_reg),
                                               .desc_11_xuser_12_reg(desc_11_xuser_12_reg),
                                               .desc_11_xuser_13_reg(desc_11_xuser_13_reg),
                                               .desc_11_xuser_14_reg(desc_11_xuser_14_reg),
                                               .desc_11_xuser_15_reg(desc_11_xuser_15_reg),
                                               .desc_11_wuser_0_reg(desc_11_wuser_0_reg),
                                               .desc_11_wuser_1_reg(desc_11_wuser_1_reg),
                                               .desc_11_wuser_2_reg(desc_11_wuser_2_reg),
                                               .desc_11_wuser_3_reg(desc_11_wuser_3_reg),
                                               .desc_11_wuser_4_reg(desc_11_wuser_4_reg),
                                               .desc_11_wuser_5_reg(desc_11_wuser_5_reg),
                                               .desc_11_wuser_6_reg(desc_11_wuser_6_reg),
                                               .desc_11_wuser_7_reg(desc_11_wuser_7_reg),
                                               .desc_11_wuser_8_reg(desc_11_wuser_8_reg),
                                               .desc_11_wuser_9_reg(desc_11_wuser_9_reg),
                                               .desc_11_wuser_10_reg(desc_11_wuser_10_reg),
                                               .desc_11_wuser_11_reg(desc_11_wuser_11_reg),
                                               .desc_11_wuser_12_reg(desc_11_wuser_12_reg),
                                               .desc_11_wuser_13_reg(desc_11_wuser_13_reg),
                                               .desc_11_wuser_14_reg(desc_11_wuser_14_reg),
                                               .desc_11_wuser_15_reg(desc_11_wuser_15_reg),
                                               .desc_12_txn_type_reg(desc_12_txn_type_reg),
                                               .desc_12_size_reg(desc_12_size_reg),
                                               .desc_12_data_offset_reg(desc_12_data_offset_reg),
                                               .desc_12_data_host_addr_0_reg(desc_12_data_host_addr_0_reg),
                                               .desc_12_data_host_addr_1_reg(desc_12_data_host_addr_1_reg),
                                               .desc_12_data_host_addr_2_reg(desc_12_data_host_addr_2_reg),
                                               .desc_12_data_host_addr_3_reg(desc_12_data_host_addr_3_reg),
                                               .desc_12_wstrb_host_addr_0_reg(desc_12_wstrb_host_addr_0_reg),
                                               .desc_12_wstrb_host_addr_1_reg(desc_12_wstrb_host_addr_1_reg),
                                               .desc_12_wstrb_host_addr_2_reg(desc_12_wstrb_host_addr_2_reg),
                                               .desc_12_wstrb_host_addr_3_reg(desc_12_wstrb_host_addr_3_reg),
                                               .desc_12_axsize_reg(desc_12_axsize_reg),
                                               .desc_12_attr_reg(desc_12_attr_reg),
                                               .desc_12_axaddr_0_reg(desc_12_axaddr_0_reg),
                                               .desc_12_axaddr_1_reg(desc_12_axaddr_1_reg),
                                               .desc_12_axaddr_2_reg(desc_12_axaddr_2_reg),
                                               .desc_12_axaddr_3_reg(desc_12_axaddr_3_reg),
                                               .desc_12_axid_0_reg(desc_12_axid_0_reg),
                                               .desc_12_axid_1_reg(desc_12_axid_1_reg),
                                               .desc_12_axid_2_reg(desc_12_axid_2_reg),
                                               .desc_12_axid_3_reg(desc_12_axid_3_reg),
                                               .desc_12_axuser_0_reg(desc_12_axuser_0_reg),
                                               .desc_12_axuser_1_reg(desc_12_axuser_1_reg),
                                               .desc_12_axuser_2_reg(desc_12_axuser_2_reg),
                                               .desc_12_axuser_3_reg(desc_12_axuser_3_reg),
                                               .desc_12_axuser_4_reg(desc_12_axuser_4_reg),
                                               .desc_12_axuser_5_reg(desc_12_axuser_5_reg),
                                               .desc_12_axuser_6_reg(desc_12_axuser_6_reg),
                                               .desc_12_axuser_7_reg(desc_12_axuser_7_reg),
                                               .desc_12_axuser_8_reg(desc_12_axuser_8_reg),
                                               .desc_12_axuser_9_reg(desc_12_axuser_9_reg),
                                               .desc_12_axuser_10_reg(desc_12_axuser_10_reg),
                                               .desc_12_axuser_11_reg(desc_12_axuser_11_reg),
                                               .desc_12_axuser_12_reg(desc_12_axuser_12_reg),
                                               .desc_12_axuser_13_reg(desc_12_axuser_13_reg),
                                               .desc_12_axuser_14_reg(desc_12_axuser_14_reg),
                                               .desc_12_axuser_15_reg(desc_12_axuser_15_reg),
                                               .desc_12_xuser_0_reg(desc_12_xuser_0_reg),
                                               .desc_12_xuser_1_reg(desc_12_xuser_1_reg),
                                               .desc_12_xuser_2_reg(desc_12_xuser_2_reg),
                                               .desc_12_xuser_3_reg(desc_12_xuser_3_reg),
                                               .desc_12_xuser_4_reg(desc_12_xuser_4_reg),
                                               .desc_12_xuser_5_reg(desc_12_xuser_5_reg),
                                               .desc_12_xuser_6_reg(desc_12_xuser_6_reg),
                                               .desc_12_xuser_7_reg(desc_12_xuser_7_reg),
                                               .desc_12_xuser_8_reg(desc_12_xuser_8_reg),
                                               .desc_12_xuser_9_reg(desc_12_xuser_9_reg),
                                               .desc_12_xuser_10_reg(desc_12_xuser_10_reg),
                                               .desc_12_xuser_11_reg(desc_12_xuser_11_reg),
                                               .desc_12_xuser_12_reg(desc_12_xuser_12_reg),
                                               .desc_12_xuser_13_reg(desc_12_xuser_13_reg),
                                               .desc_12_xuser_14_reg(desc_12_xuser_14_reg),
                                               .desc_12_xuser_15_reg(desc_12_xuser_15_reg),
                                               .desc_12_wuser_0_reg(desc_12_wuser_0_reg),
                                               .desc_12_wuser_1_reg(desc_12_wuser_1_reg),
                                               .desc_12_wuser_2_reg(desc_12_wuser_2_reg),
                                               .desc_12_wuser_3_reg(desc_12_wuser_3_reg),
                                               .desc_12_wuser_4_reg(desc_12_wuser_4_reg),
                                               .desc_12_wuser_5_reg(desc_12_wuser_5_reg),
                                               .desc_12_wuser_6_reg(desc_12_wuser_6_reg),
                                               .desc_12_wuser_7_reg(desc_12_wuser_7_reg),
                                               .desc_12_wuser_8_reg(desc_12_wuser_8_reg),
                                               .desc_12_wuser_9_reg(desc_12_wuser_9_reg),
                                               .desc_12_wuser_10_reg(desc_12_wuser_10_reg),
                                               .desc_12_wuser_11_reg(desc_12_wuser_11_reg),
                                               .desc_12_wuser_12_reg(desc_12_wuser_12_reg),
                                               .desc_12_wuser_13_reg(desc_12_wuser_13_reg),
                                               .desc_12_wuser_14_reg(desc_12_wuser_14_reg),
                                               .desc_12_wuser_15_reg(desc_12_wuser_15_reg),
                                               .desc_13_txn_type_reg(desc_13_txn_type_reg),
                                               .desc_13_size_reg(desc_13_size_reg),
                                               .desc_13_data_offset_reg(desc_13_data_offset_reg),
                                               .desc_13_data_host_addr_0_reg(desc_13_data_host_addr_0_reg),
                                               .desc_13_data_host_addr_1_reg(desc_13_data_host_addr_1_reg),
                                               .desc_13_data_host_addr_2_reg(desc_13_data_host_addr_2_reg),
                                               .desc_13_data_host_addr_3_reg(desc_13_data_host_addr_3_reg),
                                               .desc_13_wstrb_host_addr_0_reg(desc_13_wstrb_host_addr_0_reg),
                                               .desc_13_wstrb_host_addr_1_reg(desc_13_wstrb_host_addr_1_reg),
                                               .desc_13_wstrb_host_addr_2_reg(desc_13_wstrb_host_addr_2_reg),
                                               .desc_13_wstrb_host_addr_3_reg(desc_13_wstrb_host_addr_3_reg),
                                               .desc_13_axsize_reg(desc_13_axsize_reg),
                                               .desc_13_attr_reg(desc_13_attr_reg),
                                               .desc_13_axaddr_0_reg(desc_13_axaddr_0_reg),
                                               .desc_13_axaddr_1_reg(desc_13_axaddr_1_reg),
                                               .desc_13_axaddr_2_reg(desc_13_axaddr_2_reg),
                                               .desc_13_axaddr_3_reg(desc_13_axaddr_3_reg),
                                               .desc_13_axid_0_reg(desc_13_axid_0_reg),
                                               .desc_13_axid_1_reg(desc_13_axid_1_reg),
                                               .desc_13_axid_2_reg(desc_13_axid_2_reg),
                                               .desc_13_axid_3_reg(desc_13_axid_3_reg),
                                               .desc_13_axuser_0_reg(desc_13_axuser_0_reg),
                                               .desc_13_axuser_1_reg(desc_13_axuser_1_reg),
                                               .desc_13_axuser_2_reg(desc_13_axuser_2_reg),
                                               .desc_13_axuser_3_reg(desc_13_axuser_3_reg),
                                               .desc_13_axuser_4_reg(desc_13_axuser_4_reg),
                                               .desc_13_axuser_5_reg(desc_13_axuser_5_reg),
                                               .desc_13_axuser_6_reg(desc_13_axuser_6_reg),
                                               .desc_13_axuser_7_reg(desc_13_axuser_7_reg),
                                               .desc_13_axuser_8_reg(desc_13_axuser_8_reg),
                                               .desc_13_axuser_9_reg(desc_13_axuser_9_reg),
                                               .desc_13_axuser_10_reg(desc_13_axuser_10_reg),
                                               .desc_13_axuser_11_reg(desc_13_axuser_11_reg),
                                               .desc_13_axuser_12_reg(desc_13_axuser_12_reg),
                                               .desc_13_axuser_13_reg(desc_13_axuser_13_reg),
                                               .desc_13_axuser_14_reg(desc_13_axuser_14_reg),
                                               .desc_13_axuser_15_reg(desc_13_axuser_15_reg),
                                               .desc_13_xuser_0_reg(desc_13_xuser_0_reg),
                                               .desc_13_xuser_1_reg(desc_13_xuser_1_reg),
                                               .desc_13_xuser_2_reg(desc_13_xuser_2_reg),
                                               .desc_13_xuser_3_reg(desc_13_xuser_3_reg),
                                               .desc_13_xuser_4_reg(desc_13_xuser_4_reg),
                                               .desc_13_xuser_5_reg(desc_13_xuser_5_reg),
                                               .desc_13_xuser_6_reg(desc_13_xuser_6_reg),
                                               .desc_13_xuser_7_reg(desc_13_xuser_7_reg),
                                               .desc_13_xuser_8_reg(desc_13_xuser_8_reg),
                                               .desc_13_xuser_9_reg(desc_13_xuser_9_reg),
                                               .desc_13_xuser_10_reg(desc_13_xuser_10_reg),
                                               .desc_13_xuser_11_reg(desc_13_xuser_11_reg),
                                               .desc_13_xuser_12_reg(desc_13_xuser_12_reg),
                                               .desc_13_xuser_13_reg(desc_13_xuser_13_reg),
                                               .desc_13_xuser_14_reg(desc_13_xuser_14_reg),
                                               .desc_13_xuser_15_reg(desc_13_xuser_15_reg),
                                               .desc_13_wuser_0_reg(desc_13_wuser_0_reg),
                                               .desc_13_wuser_1_reg(desc_13_wuser_1_reg),
                                               .desc_13_wuser_2_reg(desc_13_wuser_2_reg),
                                               .desc_13_wuser_3_reg(desc_13_wuser_3_reg),
                                               .desc_13_wuser_4_reg(desc_13_wuser_4_reg),
                                               .desc_13_wuser_5_reg(desc_13_wuser_5_reg),
                                               .desc_13_wuser_6_reg(desc_13_wuser_6_reg),
                                               .desc_13_wuser_7_reg(desc_13_wuser_7_reg),
                                               .desc_13_wuser_8_reg(desc_13_wuser_8_reg),
                                               .desc_13_wuser_9_reg(desc_13_wuser_9_reg),
                                               .desc_13_wuser_10_reg(desc_13_wuser_10_reg),
                                               .desc_13_wuser_11_reg(desc_13_wuser_11_reg),
                                               .desc_13_wuser_12_reg(desc_13_wuser_12_reg),
                                               .desc_13_wuser_13_reg(desc_13_wuser_13_reg),
                                               .desc_13_wuser_14_reg(desc_13_wuser_14_reg),
                                               .desc_13_wuser_15_reg(desc_13_wuser_15_reg),
                                               .desc_14_txn_type_reg(desc_14_txn_type_reg),
                                               .desc_14_size_reg(desc_14_size_reg),
                                               .desc_14_data_offset_reg(desc_14_data_offset_reg),
                                               .desc_14_data_host_addr_0_reg(desc_14_data_host_addr_0_reg),
                                               .desc_14_data_host_addr_1_reg(desc_14_data_host_addr_1_reg),
                                               .desc_14_data_host_addr_2_reg(desc_14_data_host_addr_2_reg),
                                               .desc_14_data_host_addr_3_reg(desc_14_data_host_addr_3_reg),
                                               .desc_14_wstrb_host_addr_0_reg(desc_14_wstrb_host_addr_0_reg),
                                               .desc_14_wstrb_host_addr_1_reg(desc_14_wstrb_host_addr_1_reg),
                                               .desc_14_wstrb_host_addr_2_reg(desc_14_wstrb_host_addr_2_reg),
                                               .desc_14_wstrb_host_addr_3_reg(desc_14_wstrb_host_addr_3_reg),
                                               .desc_14_axsize_reg(desc_14_axsize_reg),
                                               .desc_14_attr_reg(desc_14_attr_reg),
                                               .desc_14_axaddr_0_reg(desc_14_axaddr_0_reg),
                                               .desc_14_axaddr_1_reg(desc_14_axaddr_1_reg),
                                               .desc_14_axaddr_2_reg(desc_14_axaddr_2_reg),
                                               .desc_14_axaddr_3_reg(desc_14_axaddr_3_reg),
                                               .desc_14_axid_0_reg(desc_14_axid_0_reg),
                                               .desc_14_axid_1_reg(desc_14_axid_1_reg),
                                               .desc_14_axid_2_reg(desc_14_axid_2_reg),
                                               .desc_14_axid_3_reg(desc_14_axid_3_reg),
                                               .desc_14_axuser_0_reg(desc_14_axuser_0_reg),
                                               .desc_14_axuser_1_reg(desc_14_axuser_1_reg),
                                               .desc_14_axuser_2_reg(desc_14_axuser_2_reg),
                                               .desc_14_axuser_3_reg(desc_14_axuser_3_reg),
                                               .desc_14_axuser_4_reg(desc_14_axuser_4_reg),
                                               .desc_14_axuser_5_reg(desc_14_axuser_5_reg),
                                               .desc_14_axuser_6_reg(desc_14_axuser_6_reg),
                                               .desc_14_axuser_7_reg(desc_14_axuser_7_reg),
                                               .desc_14_axuser_8_reg(desc_14_axuser_8_reg),
                                               .desc_14_axuser_9_reg(desc_14_axuser_9_reg),
                                               .desc_14_axuser_10_reg(desc_14_axuser_10_reg),
                                               .desc_14_axuser_11_reg(desc_14_axuser_11_reg),
                                               .desc_14_axuser_12_reg(desc_14_axuser_12_reg),
                                               .desc_14_axuser_13_reg(desc_14_axuser_13_reg),
                                               .desc_14_axuser_14_reg(desc_14_axuser_14_reg),
                                               .desc_14_axuser_15_reg(desc_14_axuser_15_reg),
                                               .desc_14_xuser_0_reg(desc_14_xuser_0_reg),
                                               .desc_14_xuser_1_reg(desc_14_xuser_1_reg),
                                               .desc_14_xuser_2_reg(desc_14_xuser_2_reg),
                                               .desc_14_xuser_3_reg(desc_14_xuser_3_reg),
                                               .desc_14_xuser_4_reg(desc_14_xuser_4_reg),
                                               .desc_14_xuser_5_reg(desc_14_xuser_5_reg),
                                               .desc_14_xuser_6_reg(desc_14_xuser_6_reg),
                                               .desc_14_xuser_7_reg(desc_14_xuser_7_reg),
                                               .desc_14_xuser_8_reg(desc_14_xuser_8_reg),
                                               .desc_14_xuser_9_reg(desc_14_xuser_9_reg),
                                               .desc_14_xuser_10_reg(desc_14_xuser_10_reg),
                                               .desc_14_xuser_11_reg(desc_14_xuser_11_reg),
                                               .desc_14_xuser_12_reg(desc_14_xuser_12_reg),
                                               .desc_14_xuser_13_reg(desc_14_xuser_13_reg),
                                               .desc_14_xuser_14_reg(desc_14_xuser_14_reg),
                                               .desc_14_xuser_15_reg(desc_14_xuser_15_reg),
                                               .desc_14_wuser_0_reg(desc_14_wuser_0_reg),
                                               .desc_14_wuser_1_reg(desc_14_wuser_1_reg),
                                               .desc_14_wuser_2_reg(desc_14_wuser_2_reg),
                                               .desc_14_wuser_3_reg(desc_14_wuser_3_reg),
                                               .desc_14_wuser_4_reg(desc_14_wuser_4_reg),
                                               .desc_14_wuser_5_reg(desc_14_wuser_5_reg),
                                               .desc_14_wuser_6_reg(desc_14_wuser_6_reg),
                                               .desc_14_wuser_7_reg(desc_14_wuser_7_reg),
                                               .desc_14_wuser_8_reg(desc_14_wuser_8_reg),
                                               .desc_14_wuser_9_reg(desc_14_wuser_9_reg),
                                               .desc_14_wuser_10_reg(desc_14_wuser_10_reg),
                                               .desc_14_wuser_11_reg(desc_14_wuser_11_reg),
                                               .desc_14_wuser_12_reg(desc_14_wuser_12_reg),
                                               .desc_14_wuser_13_reg(desc_14_wuser_13_reg),
                                               .desc_14_wuser_14_reg(desc_14_wuser_14_reg),
                                               .desc_14_wuser_15_reg(desc_14_wuser_15_reg),
                                               .desc_15_txn_type_reg(desc_15_txn_type_reg),
                                               .desc_15_size_reg(desc_15_size_reg),
                                               .desc_15_data_offset_reg(desc_15_data_offset_reg),
                                               .desc_15_data_host_addr_0_reg(desc_15_data_host_addr_0_reg),
                                               .desc_15_data_host_addr_1_reg(desc_15_data_host_addr_1_reg),
                                               .desc_15_data_host_addr_2_reg(desc_15_data_host_addr_2_reg),
                                               .desc_15_data_host_addr_3_reg(desc_15_data_host_addr_3_reg),
                                               .desc_15_wstrb_host_addr_0_reg(desc_15_wstrb_host_addr_0_reg),
                                               .desc_15_wstrb_host_addr_1_reg(desc_15_wstrb_host_addr_1_reg),
                                               .desc_15_wstrb_host_addr_2_reg(desc_15_wstrb_host_addr_2_reg),
                                               .desc_15_wstrb_host_addr_3_reg(desc_15_wstrb_host_addr_3_reg),
                                               .desc_15_axsize_reg(desc_15_axsize_reg),
                                               .desc_15_attr_reg(desc_15_attr_reg),
                                               .desc_15_axaddr_0_reg(desc_15_axaddr_0_reg),
                                               .desc_15_axaddr_1_reg(desc_15_axaddr_1_reg),
                                               .desc_15_axaddr_2_reg(desc_15_axaddr_2_reg),
                                               .desc_15_axaddr_3_reg(desc_15_axaddr_3_reg),
                                               .desc_15_axid_0_reg(desc_15_axid_0_reg),
                                               .desc_15_axid_1_reg(desc_15_axid_1_reg),
                                               .desc_15_axid_2_reg(desc_15_axid_2_reg),
                                               .desc_15_axid_3_reg(desc_15_axid_3_reg),
                                               .desc_15_axuser_0_reg(desc_15_axuser_0_reg),
                                               .desc_15_axuser_1_reg(desc_15_axuser_1_reg),
                                               .desc_15_axuser_2_reg(desc_15_axuser_2_reg),
                                               .desc_15_axuser_3_reg(desc_15_axuser_3_reg),
                                               .desc_15_axuser_4_reg(desc_15_axuser_4_reg),
                                               .desc_15_axuser_5_reg(desc_15_axuser_5_reg),
                                               .desc_15_axuser_6_reg(desc_15_axuser_6_reg),
                                               .desc_15_axuser_7_reg(desc_15_axuser_7_reg),
                                               .desc_15_axuser_8_reg(desc_15_axuser_8_reg),
                                               .desc_15_axuser_9_reg(desc_15_axuser_9_reg),
                                               .desc_15_axuser_10_reg(desc_15_axuser_10_reg),
                                               .desc_15_axuser_11_reg(desc_15_axuser_11_reg),
                                               .desc_15_axuser_12_reg(desc_15_axuser_12_reg),
                                               .desc_15_axuser_13_reg(desc_15_axuser_13_reg),
                                               .desc_15_axuser_14_reg(desc_15_axuser_14_reg),
                                               .desc_15_axuser_15_reg(desc_15_axuser_15_reg),
                                               .desc_15_xuser_0_reg(desc_15_xuser_0_reg),
                                               .desc_15_xuser_1_reg(desc_15_xuser_1_reg),
                                               .desc_15_xuser_2_reg(desc_15_xuser_2_reg),
                                               .desc_15_xuser_3_reg(desc_15_xuser_3_reg),
                                               .desc_15_xuser_4_reg(desc_15_xuser_4_reg),
                                               .desc_15_xuser_5_reg(desc_15_xuser_5_reg),
                                               .desc_15_xuser_6_reg(desc_15_xuser_6_reg),
                                               .desc_15_xuser_7_reg(desc_15_xuser_7_reg),
                                               .desc_15_xuser_8_reg(desc_15_xuser_8_reg),
                                               .desc_15_xuser_9_reg(desc_15_xuser_9_reg),
                                               .desc_15_xuser_10_reg(desc_15_xuser_10_reg),
                                               .desc_15_xuser_11_reg(desc_15_xuser_11_reg),
                                               .desc_15_xuser_12_reg(desc_15_xuser_12_reg),
                                               .desc_15_xuser_13_reg(desc_15_xuser_13_reg),
                                               .desc_15_xuser_14_reg(desc_15_xuser_14_reg),
                                               .desc_15_xuser_15_reg(desc_15_xuser_15_reg),
                                               .desc_15_wuser_0_reg(desc_15_wuser_0_reg),
                                               .desc_15_wuser_1_reg(desc_15_wuser_1_reg),
                                               .desc_15_wuser_2_reg(desc_15_wuser_2_reg),
                                               .desc_15_wuser_3_reg(desc_15_wuser_3_reg),
                                               .desc_15_wuser_4_reg(desc_15_wuser_4_reg),
                                               .desc_15_wuser_5_reg(desc_15_wuser_5_reg),
                                               .desc_15_wuser_6_reg(desc_15_wuser_6_reg),
                                               .desc_15_wuser_7_reg(desc_15_wuser_7_reg),
                                               .desc_15_wuser_8_reg(desc_15_wuser_8_reg),
                                               .desc_15_wuser_9_reg(desc_15_wuser_9_reg),
                                               .desc_15_wuser_10_reg(desc_15_wuser_10_reg),
                                               .desc_15_wuser_11_reg(desc_15_wuser_11_reg),
                                               .desc_15_wuser_12_reg(desc_15_wuser_12_reg),
                                               .desc_15_wuser_13_reg(desc_15_wuser_13_reg),
                                               .desc_15_wuser_14_reg(desc_15_wuser_14_reg),
                                               .desc_15_wuser_15_reg(desc_15_wuser_15_reg),
                                               .rb2uc_rd_data   (rb2uc_rd_data),
                                               .hm2uc_done      (hm2uc_done),

                                                 .s_axi_usr_awid       (s_axi_usr_awid    ),         
                                                 .s_axi_usr_awaddr     (s_axi_usr_awaddr  ),         
                                                 .s_axi_usr_awlen      (s_axi_usr_awlen   ),         
                                                 .s_axi_usr_awsize     (s_axi_usr_awsize  ),         
                                                 .s_axi_usr_awburst    (s_axi_usr_awburst ),         
                                                 .s_axi_usr_awlock     (s_axi_usr_awlock  ),         
                                                 .s_axi_usr_awcache    (s_axi_usr_awcache ),         
                                                 .s_axi_usr_awprot     (s_axi_usr_awprot  ),         
                                                 .s_axi_usr_awqos      (s_axi_usr_awqos   ),         
                                                 .s_axi_usr_awregion   (s_axi_usr_awregion),         
                                                 .s_axi_usr_awuser     (s_axi_usr_awuser  ),         
                                                 .s_axi_usr_awvalid    (s_axi_usr_awvalid ),         
                                                 .s_axi_usr_awready    (s_axi_usr_awready ),         
                                                 .s_axi_usr_wdata      (s_axi_usr_wdata   ),         
                                                 .s_axi_usr_wstrb      (s_axi_usr_wstrb   ), 
                                                 .s_axi_usr_wlast      (s_axi_usr_wlast   ),         
                                                 .s_axi_usr_wid        (s_axi_usr_wid     ),       
                                                 .s_axi_usr_wuser      (s_axi_usr_wuser   ),         
                                                 .s_axi_usr_wvalid     (s_axi_usr_wvalid  ),         
                                                 .s_axi_usr_wready     (s_axi_usr_wready  ),         
                                                 .s_axi_usr_bid        (s_axi_usr_bid     ), 
                                                 .s_axi_usr_bresp      (s_axi_usr_bresp   ),         
                                                 .s_axi_usr_buser      (s_axi_usr_buser   ),         
                                                 .s_axi_usr_bvalid     (s_axi_usr_bvalid  ),         
                                                 .s_axi_usr_bready     (s_axi_usr_bready  ),         
                                                 .s_axi_usr_arid       (s_axi_usr_arid    ), 
                                                 .s_axi_usr_araddr     (s_axi_usr_araddr  ),         
                                                 .s_axi_usr_arlen      (s_axi_usr_arlen   ),         
                                                 .s_axi_usr_arsize     (s_axi_usr_arsize  ),         
                                                 .s_axi_usr_arburst    (s_axi_usr_arburst ),         
                                                 .s_axi_usr_arlock     (s_axi_usr_arlock  ),         
                                                 .s_axi_usr_arcache    (s_axi_usr_arcache ),         
                                                 .s_axi_usr_arprot     (s_axi_usr_arprot  ),         
                                                 .s_axi_usr_arqos      (s_axi_usr_arqos   ),         
                                                 .s_axi_usr_arregion   (s_axi_usr_arregion),         
                                                 .s_axi_usr_aruser     (s_axi_usr_aruser  ),         
                                                 .s_axi_usr_arvalid    (s_axi_usr_arvalid ),         
                                                 .s_axi_usr_arready    (s_axi_usr_arready ),         
                                                 .s_axi_usr_rid        (s_axi_usr_rid     ), 
                                                 .s_axi_usr_rdata      (s_axi_usr_rdata   ),         
                                                 .s_axi_usr_rresp      (s_axi_usr_rresp   ),         
                                                 .s_axi_usr_rlast      (s_axi_usr_rlast   ),         
                                                 .s_axi_usr_ruser      (s_axi_usr_ruser   ),         
                                                 .s_axi_usr_rvalid     (s_axi_usr_rvalid  ),         
                                                 .s_axi_usr_rready     (s_axi_usr_rready  )  

       );
   
   regs_slave #(
                .EN_INTFS_AXI4          (EN_INTFS_AXI4       ),
                .EN_INTFS_AXI4LITE      (EN_INTFS_AXI4LITE   ),
                .EN_INTFS_AXI3          (EN_INTFS_AXI3       ),
                .S_AXI_ADDR_WIDTH       (S_AXI_ADDR_WIDTH    ),
                .S_AXI_DATA_WIDTH       (S_AXI_DATA_WIDTH    ),
                .RAM_SIZE               (RAM_SIZE            ),
                .S_AXI_USR_ADDR_WIDTH   (S_AXI_USR_ADDR_WIDTH), 
                .S_AXI_USR_ID_WIDTH     (S_AXI_USR_ID_WIDTH  ), 
                .S_AXI_USR_AWUSER_WIDTH (S_AXI_USR_AWUSER_WIDTH),
                .S_AXI_USR_WUSER_WIDTH  (S_AXI_USR_WUSER_WIDTH),
                .S_AXI_USR_BUSER_WIDTH  (S_AXI_USR_BUSER_WIDTH),
                .S_AXI_USR_ARUSER_WIDTH (S_AXI_USR_ARUSER_WIDTH),
                .S_AXI_USR_RUSER_WIDTH  (S_AXI_USR_RUSER_WIDTH),
                .S_AXI_USR_DATA_WIDTH   (S_AXI_USR_DATA_WIDTH),
                .MAX_DESC               (MAX_DESC            ),
		.LAST_BRIDGE		(LAST_BRIDGE),
		.EXTEND_WSTRB		(EXTEND_WSTRB),
	        .FORCE_RESP_ORDER     	(FORCE_RESP_ORDER)
                
     )
   

regs_slave_inst              (/*AUTOINST*/
                              // Outputs
                              .s_axi_awready    (s_axi_awready),
                              .s_axi_wready     (s_axi_wready),
                              .s_axi_bresp      (s_axi_bresp),
                              .s_axi_bvalid     (s_axi_bvalid),
                              .s_axi_arready    (s_axi_arready),
                              .s_axi_rdata      (s_axi_rdata),
                              .s_axi_rresp      (s_axi_rresp),
                              .s_axi_rvalid     (s_axi_rvalid),
                              .uc2rb_rd_addr    (uc2rb_rd_addr),
                              .uc2rb_wr_we      (uc2rb_wr_we),
                              .uc2rb_wr_bwe     (uc2rb_wr_bwe),
                              .uc2rb_wr_addr    (uc2rb_wr_addr),
                              .uc2rb_wr_data    (uc2rb_wr_data),
                              .uc2rb_wr_wstrb   (uc2rb_wr_wstrb),
                              .rb2hm_rd_data    (rb2hm_rd_data),
                              .rb2hm_rd_wstrb   (rb2hm_rd_wstrb),
                              .uc2hm_trig       (uc2hm_trig),
                              .version_reg      (version_reg),
                              .bridge_type_reg  (bridge_type_reg),
                              .mode_select_reg  (mode_select_reg),
                              .reset_reg        (reset_reg),
							  .h2c_intr_0_reg (h2c_intr_0_reg),
							  .h2c_intr_1_reg (h2c_intr_1_reg),
							  .h2c_intr_2_reg (h2c_intr_2_reg),
							  .h2c_intr_3_reg (h2c_intr_3_reg),
							  .h2c_gpio_0_reg (h2c_gpio_0_reg),
							  .h2c_gpio_1_reg (h2c_gpio_1_reg),
							  .h2c_gpio_2_reg (h2c_gpio_2_reg),
							  .h2c_gpio_3_reg (h2c_gpio_3_reg),
							  .h2c_gpio_4_reg (h2c_gpio_4_reg),
							  .h2c_gpio_5_reg (h2c_gpio_5_reg),
							  .h2c_gpio_6_reg (h2c_gpio_6_reg),
							  .h2c_gpio_7_reg (h2c_gpio_7_reg),
							  .c2h_intr_status_0_reg(c2h_intr_status_0_reg),
							  .c2h_intr_status_1_reg(c2h_intr_status_1_reg),
							  .intr_c2h_toggle_clear_0_reg(intr_c2h_toggle_clear_0_reg),
							  .intr_c2h_toggle_clear_1_reg(intr_c2h_toggle_clear_1_reg),
							  .intr_c2h_toggle_status_0_reg(intr_c2h_toggle_status_0_reg),
							  .intr_c2h_toggle_status_1_reg(intr_c2h_toggle_status_1_reg),
							  .intr_c2h_toggle_enable_0_reg(intr_c2h_toggle_enable_0_reg),
							  .intr_c2h_toggle_enable_1_reg(intr_c2h_toggle_enable_1_reg),
							  .c2h_gpio_0_reg(c2h_gpio_0_reg),
							  .c2h_gpio_1_reg(c2h_gpio_1_reg),
							  .c2h_gpio_2_reg(c2h_gpio_2_reg),
							  .c2h_gpio_3_reg(c2h_gpio_3_reg),
							  .c2h_gpio_4_reg(c2h_gpio_4_reg),
							  .c2h_gpio_5_reg(c2h_gpio_5_reg),
							  .c2h_gpio_6_reg(c2h_gpio_6_reg),
							  .c2h_gpio_7_reg(c2h_gpio_7_reg),
							  .c2h_gpio_8_reg(c2h_gpio_8_reg),
							  .c2h_gpio_9_reg(c2h_gpio_9_reg),
							  .c2h_gpio_10_reg(c2h_gpio_10_reg),
							  .c2h_gpio_11_reg(c2h_gpio_11_reg),
							  .c2h_gpio_12_reg(c2h_gpio_12_reg),
							  .c2h_gpio_13_reg(c2h_gpio_13_reg),
							  .c2h_gpio_14_reg(c2h_gpio_14_reg),
							  .c2h_gpio_15_reg(c2h_gpio_15_reg),
                              .axi_bridge_config_reg(axi_bridge_config_reg),
                              .axi_max_desc_reg (axi_max_desc_reg),
                              .intr_status_reg  (intr_status_reg),
                              .intr_error_status_reg(intr_error_status_reg),
                              .intr_error_clear_reg(intr_error_clear_reg),
                              .intr_error_enable_reg(intr_error_enable_reg),
                              .addr_in_0_reg    (addr_in_0_reg),
                              .addr_in_1_reg    (addr_in_1_reg),
                              .addr_in_2_reg    (addr_in_2_reg),
                              .addr_in_3_reg    (addr_in_3_reg),
                              .trans_mask_0_reg (trans_mask_0_reg),
                              .trans_mask_1_reg (trans_mask_1_reg),
                              .trans_mask_2_reg (trans_mask_2_reg),
                              .trans_mask_3_reg (trans_mask_3_reg),
                              .trans_addr_0_reg (trans_addr_0_reg),
                              .trans_addr_1_reg (trans_addr_1_reg),
                              .trans_addr_2_reg (trans_addr_2_reg),
                              .trans_addr_3_reg (trans_addr_3_reg),
                              .ownership_reg    (ownership_reg),
                              .ownership_flip_reg(ownership_flip_reg),
                              .status_resp_reg  (status_resp_reg),
                              .intr_txn_avail_status_reg(intr_txn_avail_status_reg),
                              .intr_txn_avail_clear_reg(intr_txn_avail_clear_reg),
                              .intr_txn_avail_enable_reg(intr_txn_avail_enable_reg),
                              .intr_comp_status_reg(intr_comp_status_reg),
                              .intr_comp_clear_reg(intr_comp_clear_reg),
                              .intr_comp_enable_reg(intr_comp_enable_reg),
                              .status_resp_comp_reg(status_resp_comp_reg),
                              .status_busy_reg  (status_busy_reg),
                              .resp_fifo_free_level_reg(resp_fifo_free_level_reg),
                              .resp_order_reg(resp_order_reg),
                              .desc_0_txn_type_reg(desc_0_txn_type_reg),
                              .desc_0_size_reg  (desc_0_size_reg),
                              .desc_0_data_offset_reg(desc_0_data_offset_reg),
                              .desc_0_data_host_addr_0_reg(desc_0_data_host_addr_0_reg),
                              .desc_0_data_host_addr_1_reg(desc_0_data_host_addr_1_reg),
                              .desc_0_data_host_addr_2_reg(desc_0_data_host_addr_2_reg),
                              .desc_0_data_host_addr_3_reg(desc_0_data_host_addr_3_reg),
                              .desc_0_wstrb_host_addr_0_reg(desc_0_wstrb_host_addr_0_reg),
                              .desc_0_wstrb_host_addr_1_reg(desc_0_wstrb_host_addr_1_reg),
                              .desc_0_wstrb_host_addr_2_reg(desc_0_wstrb_host_addr_2_reg),
                              .desc_0_wstrb_host_addr_3_reg(desc_0_wstrb_host_addr_3_reg),
                              .desc_0_axsize_reg(desc_0_axsize_reg),
                              .desc_0_attr_reg  (desc_0_attr_reg),
                              .desc_0_axaddr_0_reg(desc_0_axaddr_0_reg),
                              .desc_0_axaddr_1_reg(desc_0_axaddr_1_reg),
                              .desc_0_axaddr_2_reg(desc_0_axaddr_2_reg),
                              .desc_0_axaddr_3_reg(desc_0_axaddr_3_reg),
                              .desc_0_axid_0_reg(desc_0_axid_0_reg),
                              .desc_0_axid_1_reg(desc_0_axid_1_reg),
                              .desc_0_axid_2_reg(desc_0_axid_2_reg),
                              .desc_0_axid_3_reg(desc_0_axid_3_reg),
                              .desc_0_axuser_0_reg(desc_0_axuser_0_reg),
                              .desc_0_axuser_1_reg(desc_0_axuser_1_reg),
                              .desc_0_axuser_2_reg(desc_0_axuser_2_reg),
                              .desc_0_axuser_3_reg(desc_0_axuser_3_reg),
                              .desc_0_axuser_4_reg(desc_0_axuser_4_reg),
                              .desc_0_axuser_5_reg(desc_0_axuser_5_reg),
                              .desc_0_axuser_6_reg(desc_0_axuser_6_reg),
                              .desc_0_axuser_7_reg(desc_0_axuser_7_reg),
                              .desc_0_axuser_8_reg(desc_0_axuser_8_reg),
                              .desc_0_axuser_9_reg(desc_0_axuser_9_reg),
                              .desc_0_axuser_10_reg(desc_0_axuser_10_reg),
                              .desc_0_axuser_11_reg(desc_0_axuser_11_reg),
                              .desc_0_axuser_12_reg(desc_0_axuser_12_reg),
                              .desc_0_axuser_13_reg(desc_0_axuser_13_reg),
                              .desc_0_axuser_14_reg(desc_0_axuser_14_reg),
                              .desc_0_axuser_15_reg(desc_0_axuser_15_reg),
                              .desc_0_xuser_0_reg(desc_0_xuser_0_reg),
                              .desc_0_xuser_1_reg(desc_0_xuser_1_reg),
                              .desc_0_xuser_2_reg(desc_0_xuser_2_reg),
                              .desc_0_xuser_3_reg(desc_0_xuser_3_reg),
                              .desc_0_xuser_4_reg(desc_0_xuser_4_reg),
                              .desc_0_xuser_5_reg(desc_0_xuser_5_reg),
                              .desc_0_xuser_6_reg(desc_0_xuser_6_reg),
                              .desc_0_xuser_7_reg(desc_0_xuser_7_reg),
                              .desc_0_xuser_8_reg(desc_0_xuser_8_reg),
                              .desc_0_xuser_9_reg(desc_0_xuser_9_reg),
                              .desc_0_xuser_10_reg(desc_0_xuser_10_reg),
                              .desc_0_xuser_11_reg(desc_0_xuser_11_reg),
                              .desc_0_xuser_12_reg(desc_0_xuser_12_reg),
                              .desc_0_xuser_13_reg(desc_0_xuser_13_reg),
                              .desc_0_xuser_14_reg(desc_0_xuser_14_reg),
                              .desc_0_xuser_15_reg(desc_0_xuser_15_reg),
                              .desc_0_wuser_0_reg(desc_0_wuser_0_reg),
                              .desc_0_wuser_1_reg(desc_0_wuser_1_reg),
                              .desc_0_wuser_2_reg(desc_0_wuser_2_reg),
                              .desc_0_wuser_3_reg(desc_0_wuser_3_reg),
                              .desc_0_wuser_4_reg(desc_0_wuser_4_reg),
                              .desc_0_wuser_5_reg(desc_0_wuser_5_reg),
                              .desc_0_wuser_6_reg(desc_0_wuser_6_reg),
                              .desc_0_wuser_7_reg(desc_0_wuser_7_reg),
                              .desc_0_wuser_8_reg(desc_0_wuser_8_reg),
                              .desc_0_wuser_9_reg(desc_0_wuser_9_reg),
                              .desc_0_wuser_10_reg(desc_0_wuser_10_reg),
                              .desc_0_wuser_11_reg(desc_0_wuser_11_reg),
                              .desc_0_wuser_12_reg(desc_0_wuser_12_reg),
                              .desc_0_wuser_13_reg(desc_0_wuser_13_reg),
                              .desc_0_wuser_14_reg(desc_0_wuser_14_reg),
                              .desc_0_wuser_15_reg(desc_0_wuser_15_reg),
                              .desc_1_txn_type_reg(desc_1_txn_type_reg),
                              .desc_1_size_reg  (desc_1_size_reg),
                              .desc_1_data_offset_reg(desc_1_data_offset_reg),
                              .desc_1_data_host_addr_0_reg(desc_1_data_host_addr_0_reg),
                              .desc_1_data_host_addr_1_reg(desc_1_data_host_addr_1_reg),
                              .desc_1_data_host_addr_2_reg(desc_1_data_host_addr_2_reg),
                              .desc_1_data_host_addr_3_reg(desc_1_data_host_addr_3_reg),
                              .desc_1_wstrb_host_addr_0_reg(desc_1_wstrb_host_addr_0_reg),
                              .desc_1_wstrb_host_addr_1_reg(desc_1_wstrb_host_addr_1_reg),
                              .desc_1_wstrb_host_addr_2_reg(desc_1_wstrb_host_addr_2_reg),
                              .desc_1_wstrb_host_addr_3_reg(desc_1_wstrb_host_addr_3_reg),
                              .desc_1_axsize_reg(desc_1_axsize_reg),
                              .desc_1_attr_reg  (desc_1_attr_reg),
                              .desc_1_axaddr_0_reg(desc_1_axaddr_0_reg),
                              .desc_1_axaddr_1_reg(desc_1_axaddr_1_reg),
                              .desc_1_axaddr_2_reg(desc_1_axaddr_2_reg),
                              .desc_1_axaddr_3_reg(desc_1_axaddr_3_reg),
                              .desc_1_axid_0_reg(desc_1_axid_0_reg),
                              .desc_1_axid_1_reg(desc_1_axid_1_reg),
                              .desc_1_axid_2_reg(desc_1_axid_2_reg),
                              .desc_1_axid_3_reg(desc_1_axid_3_reg),
                              .desc_1_axuser_0_reg(desc_1_axuser_0_reg),
                              .desc_1_axuser_1_reg(desc_1_axuser_1_reg),
                              .desc_1_axuser_2_reg(desc_1_axuser_2_reg),
                              .desc_1_axuser_3_reg(desc_1_axuser_3_reg),
                              .desc_1_axuser_4_reg(desc_1_axuser_4_reg),
                              .desc_1_axuser_5_reg(desc_1_axuser_5_reg),
                              .desc_1_axuser_6_reg(desc_1_axuser_6_reg),
                              .desc_1_axuser_7_reg(desc_1_axuser_7_reg),
                              .desc_1_axuser_8_reg(desc_1_axuser_8_reg),
                              .desc_1_axuser_9_reg(desc_1_axuser_9_reg),
                              .desc_1_axuser_10_reg(desc_1_axuser_10_reg),
                              .desc_1_axuser_11_reg(desc_1_axuser_11_reg),
                              .desc_1_axuser_12_reg(desc_1_axuser_12_reg),
                              .desc_1_axuser_13_reg(desc_1_axuser_13_reg),
                              .desc_1_axuser_14_reg(desc_1_axuser_14_reg),
                              .desc_1_axuser_15_reg(desc_1_axuser_15_reg),
                              .desc_1_xuser_0_reg(desc_1_xuser_0_reg),
                              .desc_1_xuser_1_reg(desc_1_xuser_1_reg),
                              .desc_1_xuser_2_reg(desc_1_xuser_2_reg),
                              .desc_1_xuser_3_reg(desc_1_xuser_3_reg),
                              .desc_1_xuser_4_reg(desc_1_xuser_4_reg),
                              .desc_1_xuser_5_reg(desc_1_xuser_5_reg),
                              .desc_1_xuser_6_reg(desc_1_xuser_6_reg),
                              .desc_1_xuser_7_reg(desc_1_xuser_7_reg),
                              .desc_1_xuser_8_reg(desc_1_xuser_8_reg),
                              .desc_1_xuser_9_reg(desc_1_xuser_9_reg),
                              .desc_1_xuser_10_reg(desc_1_xuser_10_reg),
                              .desc_1_xuser_11_reg(desc_1_xuser_11_reg),
                              .desc_1_xuser_12_reg(desc_1_xuser_12_reg),
                              .desc_1_xuser_13_reg(desc_1_xuser_13_reg),
                              .desc_1_xuser_14_reg(desc_1_xuser_14_reg),
                              .desc_1_xuser_15_reg(desc_1_xuser_15_reg),
                              .desc_1_wuser_0_reg(desc_1_wuser_0_reg),
                              .desc_1_wuser_1_reg(desc_1_wuser_1_reg),
                              .desc_1_wuser_2_reg(desc_1_wuser_2_reg),
                              .desc_1_wuser_3_reg(desc_1_wuser_3_reg),
                              .desc_1_wuser_4_reg(desc_1_wuser_4_reg),
                              .desc_1_wuser_5_reg(desc_1_wuser_5_reg),
                              .desc_1_wuser_6_reg(desc_1_wuser_6_reg),
                              .desc_1_wuser_7_reg(desc_1_wuser_7_reg),
                              .desc_1_wuser_8_reg(desc_1_wuser_8_reg),
                              .desc_1_wuser_9_reg(desc_1_wuser_9_reg),
                              .desc_1_wuser_10_reg(desc_1_wuser_10_reg),
                              .desc_1_wuser_11_reg(desc_1_wuser_11_reg),
                              .desc_1_wuser_12_reg(desc_1_wuser_12_reg),
                              .desc_1_wuser_13_reg(desc_1_wuser_13_reg),
                              .desc_1_wuser_14_reg(desc_1_wuser_14_reg),
                              .desc_1_wuser_15_reg(desc_1_wuser_15_reg),
                              .desc_2_txn_type_reg(desc_2_txn_type_reg),
                              .desc_2_size_reg  (desc_2_size_reg),
                              .desc_2_data_offset_reg(desc_2_data_offset_reg),
                              .desc_2_data_host_addr_0_reg(desc_2_data_host_addr_0_reg),
                              .desc_2_data_host_addr_1_reg(desc_2_data_host_addr_1_reg),
                              .desc_2_data_host_addr_2_reg(desc_2_data_host_addr_2_reg),
                              .desc_2_data_host_addr_3_reg(desc_2_data_host_addr_3_reg),
                              .desc_2_wstrb_host_addr_0_reg(desc_2_wstrb_host_addr_0_reg),
                              .desc_2_wstrb_host_addr_1_reg(desc_2_wstrb_host_addr_1_reg),
                              .desc_2_wstrb_host_addr_2_reg(desc_2_wstrb_host_addr_2_reg),
                              .desc_2_wstrb_host_addr_3_reg(desc_2_wstrb_host_addr_3_reg),
                              .desc_2_axsize_reg(desc_2_axsize_reg),
                              .desc_2_attr_reg  (desc_2_attr_reg),
                              .desc_2_axaddr_0_reg(desc_2_axaddr_0_reg),
                              .desc_2_axaddr_1_reg(desc_2_axaddr_1_reg),
                              .desc_2_axaddr_2_reg(desc_2_axaddr_2_reg),
                              .desc_2_axaddr_3_reg(desc_2_axaddr_3_reg),
                              .desc_2_axid_0_reg(desc_2_axid_0_reg),
                              .desc_2_axid_1_reg(desc_2_axid_1_reg),
                              .desc_2_axid_2_reg(desc_2_axid_2_reg),
                              .desc_2_axid_3_reg(desc_2_axid_3_reg),
                              .desc_2_axuser_0_reg(desc_2_axuser_0_reg),
                              .desc_2_axuser_1_reg(desc_2_axuser_1_reg),
                              .desc_2_axuser_2_reg(desc_2_axuser_2_reg),
                              .desc_2_axuser_3_reg(desc_2_axuser_3_reg),
                              .desc_2_axuser_4_reg(desc_2_axuser_4_reg),
                              .desc_2_axuser_5_reg(desc_2_axuser_5_reg),
                              .desc_2_axuser_6_reg(desc_2_axuser_6_reg),
                              .desc_2_axuser_7_reg(desc_2_axuser_7_reg),
                              .desc_2_axuser_8_reg(desc_2_axuser_8_reg),
                              .desc_2_axuser_9_reg(desc_2_axuser_9_reg),
                              .desc_2_axuser_10_reg(desc_2_axuser_10_reg),
                              .desc_2_axuser_11_reg(desc_2_axuser_11_reg),
                              .desc_2_axuser_12_reg(desc_2_axuser_12_reg),
                              .desc_2_axuser_13_reg(desc_2_axuser_13_reg),
                              .desc_2_axuser_14_reg(desc_2_axuser_14_reg),
                              .desc_2_axuser_15_reg(desc_2_axuser_15_reg),
                              .desc_2_xuser_0_reg(desc_2_xuser_0_reg),
                              .desc_2_xuser_1_reg(desc_2_xuser_1_reg),
                              .desc_2_xuser_2_reg(desc_2_xuser_2_reg),
                              .desc_2_xuser_3_reg(desc_2_xuser_3_reg),
                              .desc_2_xuser_4_reg(desc_2_xuser_4_reg),
                              .desc_2_xuser_5_reg(desc_2_xuser_5_reg),
                              .desc_2_xuser_6_reg(desc_2_xuser_6_reg),
                              .desc_2_xuser_7_reg(desc_2_xuser_7_reg),
                              .desc_2_xuser_8_reg(desc_2_xuser_8_reg),
                              .desc_2_xuser_9_reg(desc_2_xuser_9_reg),
                              .desc_2_xuser_10_reg(desc_2_xuser_10_reg),
                              .desc_2_xuser_11_reg(desc_2_xuser_11_reg),
                              .desc_2_xuser_12_reg(desc_2_xuser_12_reg),
                              .desc_2_xuser_13_reg(desc_2_xuser_13_reg),
                              .desc_2_xuser_14_reg(desc_2_xuser_14_reg),
                              .desc_2_xuser_15_reg(desc_2_xuser_15_reg),
                              .desc_2_wuser_0_reg(desc_2_wuser_0_reg),
                              .desc_2_wuser_1_reg(desc_2_wuser_1_reg),
                              .desc_2_wuser_2_reg(desc_2_wuser_2_reg),
                              .desc_2_wuser_3_reg(desc_2_wuser_3_reg),
                              .desc_2_wuser_4_reg(desc_2_wuser_4_reg),
                              .desc_2_wuser_5_reg(desc_2_wuser_5_reg),
                              .desc_2_wuser_6_reg(desc_2_wuser_6_reg),
                              .desc_2_wuser_7_reg(desc_2_wuser_7_reg),
                              .desc_2_wuser_8_reg(desc_2_wuser_8_reg),
                              .desc_2_wuser_9_reg(desc_2_wuser_9_reg),
                              .desc_2_wuser_10_reg(desc_2_wuser_10_reg),
                              .desc_2_wuser_11_reg(desc_2_wuser_11_reg),
                              .desc_2_wuser_12_reg(desc_2_wuser_12_reg),
                              .desc_2_wuser_13_reg(desc_2_wuser_13_reg),
                              .desc_2_wuser_14_reg(desc_2_wuser_14_reg),
                              .desc_2_wuser_15_reg(desc_2_wuser_15_reg),
                              .desc_3_txn_type_reg(desc_3_txn_type_reg),
                              .desc_3_size_reg  (desc_3_size_reg),
                              .desc_3_data_offset_reg(desc_3_data_offset_reg),
                              .desc_3_data_host_addr_0_reg(desc_3_data_host_addr_0_reg),
                              .desc_3_data_host_addr_1_reg(desc_3_data_host_addr_1_reg),
                              .desc_3_data_host_addr_2_reg(desc_3_data_host_addr_2_reg),
                              .desc_3_data_host_addr_3_reg(desc_3_data_host_addr_3_reg),
                              .desc_3_wstrb_host_addr_0_reg(desc_3_wstrb_host_addr_0_reg),
                              .desc_3_wstrb_host_addr_1_reg(desc_3_wstrb_host_addr_1_reg),
                              .desc_3_wstrb_host_addr_2_reg(desc_3_wstrb_host_addr_2_reg),
                              .desc_3_wstrb_host_addr_3_reg(desc_3_wstrb_host_addr_3_reg),
                              .desc_3_axsize_reg(desc_3_axsize_reg),
                              .desc_3_attr_reg  (desc_3_attr_reg),
                              .desc_3_axaddr_0_reg(desc_3_axaddr_0_reg),
                              .desc_3_axaddr_1_reg(desc_3_axaddr_1_reg),
                              .desc_3_axaddr_2_reg(desc_3_axaddr_2_reg),
                              .desc_3_axaddr_3_reg(desc_3_axaddr_3_reg),
                              .desc_3_axid_0_reg(desc_3_axid_0_reg),
                              .desc_3_axid_1_reg(desc_3_axid_1_reg),
                              .desc_3_axid_2_reg(desc_3_axid_2_reg),
                              .desc_3_axid_3_reg(desc_3_axid_3_reg),
                              .desc_3_axuser_0_reg(desc_3_axuser_0_reg),
                              .desc_3_axuser_1_reg(desc_3_axuser_1_reg),
                              .desc_3_axuser_2_reg(desc_3_axuser_2_reg),
                              .desc_3_axuser_3_reg(desc_3_axuser_3_reg),
                              .desc_3_axuser_4_reg(desc_3_axuser_4_reg),
                              .desc_3_axuser_5_reg(desc_3_axuser_5_reg),
                              .desc_3_axuser_6_reg(desc_3_axuser_6_reg),
                              .desc_3_axuser_7_reg(desc_3_axuser_7_reg),
                              .desc_3_axuser_8_reg(desc_3_axuser_8_reg),
                              .desc_3_axuser_9_reg(desc_3_axuser_9_reg),
                              .desc_3_axuser_10_reg(desc_3_axuser_10_reg),
                              .desc_3_axuser_11_reg(desc_3_axuser_11_reg),
                              .desc_3_axuser_12_reg(desc_3_axuser_12_reg),
                              .desc_3_axuser_13_reg(desc_3_axuser_13_reg),
                              .desc_3_axuser_14_reg(desc_3_axuser_14_reg),
                              .desc_3_axuser_15_reg(desc_3_axuser_15_reg),
                              .desc_3_xuser_0_reg(desc_3_xuser_0_reg),
                              .desc_3_xuser_1_reg(desc_3_xuser_1_reg),
                              .desc_3_xuser_2_reg(desc_3_xuser_2_reg),
                              .desc_3_xuser_3_reg(desc_3_xuser_3_reg),
                              .desc_3_xuser_4_reg(desc_3_xuser_4_reg),
                              .desc_3_xuser_5_reg(desc_3_xuser_5_reg),
                              .desc_3_xuser_6_reg(desc_3_xuser_6_reg),
                              .desc_3_xuser_7_reg(desc_3_xuser_7_reg),
                              .desc_3_xuser_8_reg(desc_3_xuser_8_reg),
                              .desc_3_xuser_9_reg(desc_3_xuser_9_reg),
                              .desc_3_xuser_10_reg(desc_3_xuser_10_reg),
                              .desc_3_xuser_11_reg(desc_3_xuser_11_reg),
                              .desc_3_xuser_12_reg(desc_3_xuser_12_reg),
                              .desc_3_xuser_13_reg(desc_3_xuser_13_reg),
                              .desc_3_xuser_14_reg(desc_3_xuser_14_reg),
                              .desc_3_xuser_15_reg(desc_3_xuser_15_reg),
                              .desc_3_wuser_0_reg(desc_3_wuser_0_reg),
                              .desc_3_wuser_1_reg(desc_3_wuser_1_reg),
                              .desc_3_wuser_2_reg(desc_3_wuser_2_reg),
                              .desc_3_wuser_3_reg(desc_3_wuser_3_reg),
                              .desc_3_wuser_4_reg(desc_3_wuser_4_reg),
                              .desc_3_wuser_5_reg(desc_3_wuser_5_reg),
                              .desc_3_wuser_6_reg(desc_3_wuser_6_reg),
                              .desc_3_wuser_7_reg(desc_3_wuser_7_reg),
                              .desc_3_wuser_8_reg(desc_3_wuser_8_reg),
                              .desc_3_wuser_9_reg(desc_3_wuser_9_reg),
                              .desc_3_wuser_10_reg(desc_3_wuser_10_reg),
                              .desc_3_wuser_11_reg(desc_3_wuser_11_reg),
                              .desc_3_wuser_12_reg(desc_3_wuser_12_reg),
                              .desc_3_wuser_13_reg(desc_3_wuser_13_reg),
                              .desc_3_wuser_14_reg(desc_3_wuser_14_reg),
                              .desc_3_wuser_15_reg(desc_3_wuser_15_reg),
                              .desc_4_txn_type_reg(desc_4_txn_type_reg),
                              .desc_4_size_reg  (desc_4_size_reg),
                              .desc_4_data_offset_reg(desc_4_data_offset_reg),
                              .desc_4_data_host_addr_0_reg(desc_4_data_host_addr_0_reg),
                              .desc_4_data_host_addr_1_reg(desc_4_data_host_addr_1_reg),
                              .desc_4_data_host_addr_2_reg(desc_4_data_host_addr_2_reg),
                              .desc_4_data_host_addr_3_reg(desc_4_data_host_addr_3_reg),
                              .desc_4_wstrb_host_addr_0_reg(desc_4_wstrb_host_addr_0_reg),
                              .desc_4_wstrb_host_addr_1_reg(desc_4_wstrb_host_addr_1_reg),
                              .desc_4_wstrb_host_addr_2_reg(desc_4_wstrb_host_addr_2_reg),
                              .desc_4_wstrb_host_addr_3_reg(desc_4_wstrb_host_addr_3_reg),
                              .desc_4_axsize_reg(desc_4_axsize_reg),
                              .desc_4_attr_reg  (desc_4_attr_reg),
                              .desc_4_axaddr_0_reg(desc_4_axaddr_0_reg),
                              .desc_4_axaddr_1_reg(desc_4_axaddr_1_reg),
                              .desc_4_axaddr_2_reg(desc_4_axaddr_2_reg),
                              .desc_4_axaddr_3_reg(desc_4_axaddr_3_reg),
                              .desc_4_axid_0_reg(desc_4_axid_0_reg),
                              .desc_4_axid_1_reg(desc_4_axid_1_reg),
                              .desc_4_axid_2_reg(desc_4_axid_2_reg),
                              .desc_4_axid_3_reg(desc_4_axid_3_reg),
                              .desc_4_axuser_0_reg(desc_4_axuser_0_reg),
                              .desc_4_axuser_1_reg(desc_4_axuser_1_reg),
                              .desc_4_axuser_2_reg(desc_4_axuser_2_reg),
                              .desc_4_axuser_3_reg(desc_4_axuser_3_reg),
                              .desc_4_axuser_4_reg(desc_4_axuser_4_reg),
                              .desc_4_axuser_5_reg(desc_4_axuser_5_reg),
                              .desc_4_axuser_6_reg(desc_4_axuser_6_reg),
                              .desc_4_axuser_7_reg(desc_4_axuser_7_reg),
                              .desc_4_axuser_8_reg(desc_4_axuser_8_reg),
                              .desc_4_axuser_9_reg(desc_4_axuser_9_reg),
                              .desc_4_axuser_10_reg(desc_4_axuser_10_reg),
                              .desc_4_axuser_11_reg(desc_4_axuser_11_reg),
                              .desc_4_axuser_12_reg(desc_4_axuser_12_reg),
                              .desc_4_axuser_13_reg(desc_4_axuser_13_reg),
                              .desc_4_axuser_14_reg(desc_4_axuser_14_reg),
                              .desc_4_axuser_15_reg(desc_4_axuser_15_reg),
                              .desc_4_xuser_0_reg(desc_4_xuser_0_reg),
                              .desc_4_xuser_1_reg(desc_4_xuser_1_reg),
                              .desc_4_xuser_2_reg(desc_4_xuser_2_reg),
                              .desc_4_xuser_3_reg(desc_4_xuser_3_reg),
                              .desc_4_xuser_4_reg(desc_4_xuser_4_reg),
                              .desc_4_xuser_5_reg(desc_4_xuser_5_reg),
                              .desc_4_xuser_6_reg(desc_4_xuser_6_reg),
                              .desc_4_xuser_7_reg(desc_4_xuser_7_reg),
                              .desc_4_xuser_8_reg(desc_4_xuser_8_reg),
                              .desc_4_xuser_9_reg(desc_4_xuser_9_reg),
                              .desc_4_xuser_10_reg(desc_4_xuser_10_reg),
                              .desc_4_xuser_11_reg(desc_4_xuser_11_reg),
                              .desc_4_xuser_12_reg(desc_4_xuser_12_reg),
                              .desc_4_xuser_13_reg(desc_4_xuser_13_reg),
                              .desc_4_xuser_14_reg(desc_4_xuser_14_reg),
                              .desc_4_xuser_15_reg(desc_4_xuser_15_reg),
                              .desc_4_wuser_0_reg(desc_4_wuser_0_reg),
                              .desc_4_wuser_1_reg(desc_4_wuser_1_reg),
                              .desc_4_wuser_2_reg(desc_4_wuser_2_reg),
                              .desc_4_wuser_3_reg(desc_4_wuser_3_reg),
                              .desc_4_wuser_4_reg(desc_4_wuser_4_reg),
                              .desc_4_wuser_5_reg(desc_4_wuser_5_reg),
                              .desc_4_wuser_6_reg(desc_4_wuser_6_reg),
                              .desc_4_wuser_7_reg(desc_4_wuser_7_reg),
                              .desc_4_wuser_8_reg(desc_4_wuser_8_reg),
                              .desc_4_wuser_9_reg(desc_4_wuser_9_reg),
                              .desc_4_wuser_10_reg(desc_4_wuser_10_reg),
                              .desc_4_wuser_11_reg(desc_4_wuser_11_reg),
                              .desc_4_wuser_12_reg(desc_4_wuser_12_reg),
                              .desc_4_wuser_13_reg(desc_4_wuser_13_reg),
                              .desc_4_wuser_14_reg(desc_4_wuser_14_reg),
                              .desc_4_wuser_15_reg(desc_4_wuser_15_reg),
                              .desc_5_txn_type_reg(desc_5_txn_type_reg),
                              .desc_5_size_reg  (desc_5_size_reg),
                              .desc_5_data_offset_reg(desc_5_data_offset_reg),
                              .desc_5_data_host_addr_0_reg(desc_5_data_host_addr_0_reg),
                              .desc_5_data_host_addr_1_reg(desc_5_data_host_addr_1_reg),
                              .desc_5_data_host_addr_2_reg(desc_5_data_host_addr_2_reg),
                              .desc_5_data_host_addr_3_reg(desc_5_data_host_addr_3_reg),
                              .desc_5_wstrb_host_addr_0_reg(desc_5_wstrb_host_addr_0_reg),
                              .desc_5_wstrb_host_addr_1_reg(desc_5_wstrb_host_addr_1_reg),
                              .desc_5_wstrb_host_addr_2_reg(desc_5_wstrb_host_addr_2_reg),
                              .desc_5_wstrb_host_addr_3_reg(desc_5_wstrb_host_addr_3_reg),
                              .desc_5_axsize_reg(desc_5_axsize_reg),
                              .desc_5_attr_reg  (desc_5_attr_reg),
                              .desc_5_axaddr_0_reg(desc_5_axaddr_0_reg),
                              .desc_5_axaddr_1_reg(desc_5_axaddr_1_reg),
                              .desc_5_axaddr_2_reg(desc_5_axaddr_2_reg),
                              .desc_5_axaddr_3_reg(desc_5_axaddr_3_reg),
                              .desc_5_axid_0_reg(desc_5_axid_0_reg),
                              .desc_5_axid_1_reg(desc_5_axid_1_reg),
                              .desc_5_axid_2_reg(desc_5_axid_2_reg),
                              .desc_5_axid_3_reg(desc_5_axid_3_reg),
                              .desc_5_axuser_0_reg(desc_5_axuser_0_reg),
                              .desc_5_axuser_1_reg(desc_5_axuser_1_reg),
                              .desc_5_axuser_2_reg(desc_5_axuser_2_reg),
                              .desc_5_axuser_3_reg(desc_5_axuser_3_reg),
                              .desc_5_axuser_4_reg(desc_5_axuser_4_reg),
                              .desc_5_axuser_5_reg(desc_5_axuser_5_reg),
                              .desc_5_axuser_6_reg(desc_5_axuser_6_reg),
                              .desc_5_axuser_7_reg(desc_5_axuser_7_reg),
                              .desc_5_axuser_8_reg(desc_5_axuser_8_reg),
                              .desc_5_axuser_9_reg(desc_5_axuser_9_reg),
                              .desc_5_axuser_10_reg(desc_5_axuser_10_reg),
                              .desc_5_axuser_11_reg(desc_5_axuser_11_reg),
                              .desc_5_axuser_12_reg(desc_5_axuser_12_reg),
                              .desc_5_axuser_13_reg(desc_5_axuser_13_reg),
                              .desc_5_axuser_14_reg(desc_5_axuser_14_reg),
                              .desc_5_axuser_15_reg(desc_5_axuser_15_reg),
                              .desc_5_xuser_0_reg(desc_5_xuser_0_reg),
                              .desc_5_xuser_1_reg(desc_5_xuser_1_reg),
                              .desc_5_xuser_2_reg(desc_5_xuser_2_reg),
                              .desc_5_xuser_3_reg(desc_5_xuser_3_reg),
                              .desc_5_xuser_4_reg(desc_5_xuser_4_reg),
                              .desc_5_xuser_5_reg(desc_5_xuser_5_reg),
                              .desc_5_xuser_6_reg(desc_5_xuser_6_reg),
                              .desc_5_xuser_7_reg(desc_5_xuser_7_reg),
                              .desc_5_xuser_8_reg(desc_5_xuser_8_reg),
                              .desc_5_xuser_9_reg(desc_5_xuser_9_reg),
                              .desc_5_xuser_10_reg(desc_5_xuser_10_reg),
                              .desc_5_xuser_11_reg(desc_5_xuser_11_reg),
                              .desc_5_xuser_12_reg(desc_5_xuser_12_reg),
                              .desc_5_xuser_13_reg(desc_5_xuser_13_reg),
                              .desc_5_xuser_14_reg(desc_5_xuser_14_reg),
                              .desc_5_xuser_15_reg(desc_5_xuser_15_reg),
                              .desc_5_wuser_0_reg(desc_5_wuser_0_reg),
                              .desc_5_wuser_1_reg(desc_5_wuser_1_reg),
                              .desc_5_wuser_2_reg(desc_5_wuser_2_reg),
                              .desc_5_wuser_3_reg(desc_5_wuser_3_reg),
                              .desc_5_wuser_4_reg(desc_5_wuser_4_reg),
                              .desc_5_wuser_5_reg(desc_5_wuser_5_reg),
                              .desc_5_wuser_6_reg(desc_5_wuser_6_reg),
                              .desc_5_wuser_7_reg(desc_5_wuser_7_reg),
                              .desc_5_wuser_8_reg(desc_5_wuser_8_reg),
                              .desc_5_wuser_9_reg(desc_5_wuser_9_reg),
                              .desc_5_wuser_10_reg(desc_5_wuser_10_reg),
                              .desc_5_wuser_11_reg(desc_5_wuser_11_reg),
                              .desc_5_wuser_12_reg(desc_5_wuser_12_reg),
                              .desc_5_wuser_13_reg(desc_5_wuser_13_reg),
                              .desc_5_wuser_14_reg(desc_5_wuser_14_reg),
                              .desc_5_wuser_15_reg(desc_5_wuser_15_reg),
                              .desc_6_txn_type_reg(desc_6_txn_type_reg),
                              .desc_6_size_reg  (desc_6_size_reg),
                              .desc_6_data_offset_reg(desc_6_data_offset_reg),
                              .desc_6_data_host_addr_0_reg(desc_6_data_host_addr_0_reg),
                              .desc_6_data_host_addr_1_reg(desc_6_data_host_addr_1_reg),
                              .desc_6_data_host_addr_2_reg(desc_6_data_host_addr_2_reg),
                              .desc_6_data_host_addr_3_reg(desc_6_data_host_addr_3_reg),
                              .desc_6_wstrb_host_addr_0_reg(desc_6_wstrb_host_addr_0_reg),
                              .desc_6_wstrb_host_addr_1_reg(desc_6_wstrb_host_addr_1_reg),
                              .desc_6_wstrb_host_addr_2_reg(desc_6_wstrb_host_addr_2_reg),
                              .desc_6_wstrb_host_addr_3_reg(desc_6_wstrb_host_addr_3_reg),
                              .desc_6_axsize_reg(desc_6_axsize_reg),
                              .desc_6_attr_reg  (desc_6_attr_reg),
                              .desc_6_axaddr_0_reg(desc_6_axaddr_0_reg),
                              .desc_6_axaddr_1_reg(desc_6_axaddr_1_reg),
                              .desc_6_axaddr_2_reg(desc_6_axaddr_2_reg),
                              .desc_6_axaddr_3_reg(desc_6_axaddr_3_reg),
                              .desc_6_axid_0_reg(desc_6_axid_0_reg),
                              .desc_6_axid_1_reg(desc_6_axid_1_reg),
                              .desc_6_axid_2_reg(desc_6_axid_2_reg),
                              .desc_6_axid_3_reg(desc_6_axid_3_reg),
                              .desc_6_axuser_0_reg(desc_6_axuser_0_reg),
                              .desc_6_axuser_1_reg(desc_6_axuser_1_reg),
                              .desc_6_axuser_2_reg(desc_6_axuser_2_reg),
                              .desc_6_axuser_3_reg(desc_6_axuser_3_reg),
                              .desc_6_axuser_4_reg(desc_6_axuser_4_reg),
                              .desc_6_axuser_5_reg(desc_6_axuser_5_reg),
                              .desc_6_axuser_6_reg(desc_6_axuser_6_reg),
                              .desc_6_axuser_7_reg(desc_6_axuser_7_reg),
                              .desc_6_axuser_8_reg(desc_6_axuser_8_reg),
                              .desc_6_axuser_9_reg(desc_6_axuser_9_reg),
                              .desc_6_axuser_10_reg(desc_6_axuser_10_reg),
                              .desc_6_axuser_11_reg(desc_6_axuser_11_reg),
                              .desc_6_axuser_12_reg(desc_6_axuser_12_reg),
                              .desc_6_axuser_13_reg(desc_6_axuser_13_reg),
                              .desc_6_axuser_14_reg(desc_6_axuser_14_reg),
                              .desc_6_axuser_15_reg(desc_6_axuser_15_reg),
                              .desc_6_xuser_0_reg(desc_6_xuser_0_reg),
                              .desc_6_xuser_1_reg(desc_6_xuser_1_reg),
                              .desc_6_xuser_2_reg(desc_6_xuser_2_reg),
                              .desc_6_xuser_3_reg(desc_6_xuser_3_reg),
                              .desc_6_xuser_4_reg(desc_6_xuser_4_reg),
                              .desc_6_xuser_5_reg(desc_6_xuser_5_reg),
                              .desc_6_xuser_6_reg(desc_6_xuser_6_reg),
                              .desc_6_xuser_7_reg(desc_6_xuser_7_reg),
                              .desc_6_xuser_8_reg(desc_6_xuser_8_reg),
                              .desc_6_xuser_9_reg(desc_6_xuser_9_reg),
                              .desc_6_xuser_10_reg(desc_6_xuser_10_reg),
                              .desc_6_xuser_11_reg(desc_6_xuser_11_reg),
                              .desc_6_xuser_12_reg(desc_6_xuser_12_reg),
                              .desc_6_xuser_13_reg(desc_6_xuser_13_reg),
                              .desc_6_xuser_14_reg(desc_6_xuser_14_reg),
                              .desc_6_xuser_15_reg(desc_6_xuser_15_reg),
                              .desc_6_wuser_0_reg(desc_6_wuser_0_reg),
                              .desc_6_wuser_1_reg(desc_6_wuser_1_reg),
                              .desc_6_wuser_2_reg(desc_6_wuser_2_reg),
                              .desc_6_wuser_3_reg(desc_6_wuser_3_reg),
                              .desc_6_wuser_4_reg(desc_6_wuser_4_reg),
                              .desc_6_wuser_5_reg(desc_6_wuser_5_reg),
                              .desc_6_wuser_6_reg(desc_6_wuser_6_reg),
                              .desc_6_wuser_7_reg(desc_6_wuser_7_reg),
                              .desc_6_wuser_8_reg(desc_6_wuser_8_reg),
                              .desc_6_wuser_9_reg(desc_6_wuser_9_reg),
                              .desc_6_wuser_10_reg(desc_6_wuser_10_reg),
                              .desc_6_wuser_11_reg(desc_6_wuser_11_reg),
                              .desc_6_wuser_12_reg(desc_6_wuser_12_reg),
                              .desc_6_wuser_13_reg(desc_6_wuser_13_reg),
                              .desc_6_wuser_14_reg(desc_6_wuser_14_reg),
                              .desc_6_wuser_15_reg(desc_6_wuser_15_reg),
                              .desc_7_txn_type_reg(desc_7_txn_type_reg),
                              .desc_7_size_reg  (desc_7_size_reg),
                              .desc_7_data_offset_reg(desc_7_data_offset_reg),
                              .desc_7_data_host_addr_0_reg(desc_7_data_host_addr_0_reg),
                              .desc_7_data_host_addr_1_reg(desc_7_data_host_addr_1_reg),
                              .desc_7_data_host_addr_2_reg(desc_7_data_host_addr_2_reg),
                              .desc_7_data_host_addr_3_reg(desc_7_data_host_addr_3_reg),
                              .desc_7_wstrb_host_addr_0_reg(desc_7_wstrb_host_addr_0_reg),
                              .desc_7_wstrb_host_addr_1_reg(desc_7_wstrb_host_addr_1_reg),
                              .desc_7_wstrb_host_addr_2_reg(desc_7_wstrb_host_addr_2_reg),
                              .desc_7_wstrb_host_addr_3_reg(desc_7_wstrb_host_addr_3_reg),
                              .desc_7_axsize_reg(desc_7_axsize_reg),
                              .desc_7_attr_reg  (desc_7_attr_reg),
                              .desc_7_axaddr_0_reg(desc_7_axaddr_0_reg),
                              .desc_7_axaddr_1_reg(desc_7_axaddr_1_reg),
                              .desc_7_axaddr_2_reg(desc_7_axaddr_2_reg),
                              .desc_7_axaddr_3_reg(desc_7_axaddr_3_reg),
                              .desc_7_axid_0_reg(desc_7_axid_0_reg),
                              .desc_7_axid_1_reg(desc_7_axid_1_reg),
                              .desc_7_axid_2_reg(desc_7_axid_2_reg),
                              .desc_7_axid_3_reg(desc_7_axid_3_reg),
                              .desc_7_axuser_0_reg(desc_7_axuser_0_reg),
                              .desc_7_axuser_1_reg(desc_7_axuser_1_reg),
                              .desc_7_axuser_2_reg(desc_7_axuser_2_reg),
                              .desc_7_axuser_3_reg(desc_7_axuser_3_reg),
                              .desc_7_axuser_4_reg(desc_7_axuser_4_reg),
                              .desc_7_axuser_5_reg(desc_7_axuser_5_reg),
                              .desc_7_axuser_6_reg(desc_7_axuser_6_reg),
                              .desc_7_axuser_7_reg(desc_7_axuser_7_reg),
                              .desc_7_axuser_8_reg(desc_7_axuser_8_reg),
                              .desc_7_axuser_9_reg(desc_7_axuser_9_reg),
                              .desc_7_axuser_10_reg(desc_7_axuser_10_reg),
                              .desc_7_axuser_11_reg(desc_7_axuser_11_reg),
                              .desc_7_axuser_12_reg(desc_7_axuser_12_reg),
                              .desc_7_axuser_13_reg(desc_7_axuser_13_reg),
                              .desc_7_axuser_14_reg(desc_7_axuser_14_reg),
                              .desc_7_axuser_15_reg(desc_7_axuser_15_reg),
                              .desc_7_xuser_0_reg(desc_7_xuser_0_reg),
                              .desc_7_xuser_1_reg(desc_7_xuser_1_reg),
                              .desc_7_xuser_2_reg(desc_7_xuser_2_reg),
                              .desc_7_xuser_3_reg(desc_7_xuser_3_reg),
                              .desc_7_xuser_4_reg(desc_7_xuser_4_reg),
                              .desc_7_xuser_5_reg(desc_7_xuser_5_reg),
                              .desc_7_xuser_6_reg(desc_7_xuser_6_reg),
                              .desc_7_xuser_7_reg(desc_7_xuser_7_reg),
                              .desc_7_xuser_8_reg(desc_7_xuser_8_reg),
                              .desc_7_xuser_9_reg(desc_7_xuser_9_reg),
                              .desc_7_xuser_10_reg(desc_7_xuser_10_reg),
                              .desc_7_xuser_11_reg(desc_7_xuser_11_reg),
                              .desc_7_xuser_12_reg(desc_7_xuser_12_reg),
                              .desc_7_xuser_13_reg(desc_7_xuser_13_reg),
                              .desc_7_xuser_14_reg(desc_7_xuser_14_reg),
                              .desc_7_xuser_15_reg(desc_7_xuser_15_reg),
                              .desc_7_wuser_0_reg(desc_7_wuser_0_reg),
                              .desc_7_wuser_1_reg(desc_7_wuser_1_reg),
                              .desc_7_wuser_2_reg(desc_7_wuser_2_reg),
                              .desc_7_wuser_3_reg(desc_7_wuser_3_reg),
                              .desc_7_wuser_4_reg(desc_7_wuser_4_reg),
                              .desc_7_wuser_5_reg(desc_7_wuser_5_reg),
                              .desc_7_wuser_6_reg(desc_7_wuser_6_reg),
                              .desc_7_wuser_7_reg(desc_7_wuser_7_reg),
                              .desc_7_wuser_8_reg(desc_7_wuser_8_reg),
                              .desc_7_wuser_9_reg(desc_7_wuser_9_reg),
                              .desc_7_wuser_10_reg(desc_7_wuser_10_reg),
                              .desc_7_wuser_11_reg(desc_7_wuser_11_reg),
                              .desc_7_wuser_12_reg(desc_7_wuser_12_reg),
                              .desc_7_wuser_13_reg(desc_7_wuser_13_reg),
                              .desc_7_wuser_14_reg(desc_7_wuser_14_reg),
                              .desc_7_wuser_15_reg(desc_7_wuser_15_reg),
                              .desc_8_txn_type_reg(desc_8_txn_type_reg),
                              .desc_8_size_reg  (desc_8_size_reg),
                              .desc_8_data_offset_reg(desc_8_data_offset_reg),
                              .desc_8_data_host_addr_0_reg(desc_8_data_host_addr_0_reg),
                              .desc_8_data_host_addr_1_reg(desc_8_data_host_addr_1_reg),
                              .desc_8_data_host_addr_2_reg(desc_8_data_host_addr_2_reg),
                              .desc_8_data_host_addr_3_reg(desc_8_data_host_addr_3_reg),
                              .desc_8_wstrb_host_addr_0_reg(desc_8_wstrb_host_addr_0_reg),
                              .desc_8_wstrb_host_addr_1_reg(desc_8_wstrb_host_addr_1_reg),
                              .desc_8_wstrb_host_addr_2_reg(desc_8_wstrb_host_addr_2_reg),
                              .desc_8_wstrb_host_addr_3_reg(desc_8_wstrb_host_addr_3_reg),
                              .desc_8_axsize_reg(desc_8_axsize_reg),
                              .desc_8_attr_reg  (desc_8_attr_reg),
                              .desc_8_axaddr_0_reg(desc_8_axaddr_0_reg),
                              .desc_8_axaddr_1_reg(desc_8_axaddr_1_reg),
                              .desc_8_axaddr_2_reg(desc_8_axaddr_2_reg),
                              .desc_8_axaddr_3_reg(desc_8_axaddr_3_reg),
                              .desc_8_axid_0_reg(desc_8_axid_0_reg),
                              .desc_8_axid_1_reg(desc_8_axid_1_reg),
                              .desc_8_axid_2_reg(desc_8_axid_2_reg),
                              .desc_8_axid_3_reg(desc_8_axid_3_reg),
                              .desc_8_axuser_0_reg(desc_8_axuser_0_reg),
                              .desc_8_axuser_1_reg(desc_8_axuser_1_reg),
                              .desc_8_axuser_2_reg(desc_8_axuser_2_reg),
                              .desc_8_axuser_3_reg(desc_8_axuser_3_reg),
                              .desc_8_axuser_4_reg(desc_8_axuser_4_reg),
                              .desc_8_axuser_5_reg(desc_8_axuser_5_reg),
                              .desc_8_axuser_6_reg(desc_8_axuser_6_reg),
                              .desc_8_axuser_7_reg(desc_8_axuser_7_reg),
                              .desc_8_axuser_8_reg(desc_8_axuser_8_reg),
                              .desc_8_axuser_9_reg(desc_8_axuser_9_reg),
                              .desc_8_axuser_10_reg(desc_8_axuser_10_reg),
                              .desc_8_axuser_11_reg(desc_8_axuser_11_reg),
                              .desc_8_axuser_12_reg(desc_8_axuser_12_reg),
                              .desc_8_axuser_13_reg(desc_8_axuser_13_reg),
                              .desc_8_axuser_14_reg(desc_8_axuser_14_reg),
                              .desc_8_axuser_15_reg(desc_8_axuser_15_reg),
                              .desc_8_xuser_0_reg(desc_8_xuser_0_reg),
                              .desc_8_xuser_1_reg(desc_8_xuser_1_reg),
                              .desc_8_xuser_2_reg(desc_8_xuser_2_reg),
                              .desc_8_xuser_3_reg(desc_8_xuser_3_reg),
                              .desc_8_xuser_4_reg(desc_8_xuser_4_reg),
                              .desc_8_xuser_5_reg(desc_8_xuser_5_reg),
                              .desc_8_xuser_6_reg(desc_8_xuser_6_reg),
                              .desc_8_xuser_7_reg(desc_8_xuser_7_reg),
                              .desc_8_xuser_8_reg(desc_8_xuser_8_reg),
                              .desc_8_xuser_9_reg(desc_8_xuser_9_reg),
                              .desc_8_xuser_10_reg(desc_8_xuser_10_reg),
                              .desc_8_xuser_11_reg(desc_8_xuser_11_reg),
                              .desc_8_xuser_12_reg(desc_8_xuser_12_reg),
                              .desc_8_xuser_13_reg(desc_8_xuser_13_reg),
                              .desc_8_xuser_14_reg(desc_8_xuser_14_reg),
                              .desc_8_xuser_15_reg(desc_8_xuser_15_reg),
                              .desc_8_wuser_0_reg(desc_8_wuser_0_reg),
                              .desc_8_wuser_1_reg(desc_8_wuser_1_reg),
                              .desc_8_wuser_2_reg(desc_8_wuser_2_reg),
                              .desc_8_wuser_3_reg(desc_8_wuser_3_reg),
                              .desc_8_wuser_4_reg(desc_8_wuser_4_reg),
                              .desc_8_wuser_5_reg(desc_8_wuser_5_reg),
                              .desc_8_wuser_6_reg(desc_8_wuser_6_reg),
                              .desc_8_wuser_7_reg(desc_8_wuser_7_reg),
                              .desc_8_wuser_8_reg(desc_8_wuser_8_reg),
                              .desc_8_wuser_9_reg(desc_8_wuser_9_reg),
                              .desc_8_wuser_10_reg(desc_8_wuser_10_reg),
                              .desc_8_wuser_11_reg(desc_8_wuser_11_reg),
                              .desc_8_wuser_12_reg(desc_8_wuser_12_reg),
                              .desc_8_wuser_13_reg(desc_8_wuser_13_reg),
                              .desc_8_wuser_14_reg(desc_8_wuser_14_reg),
                              .desc_8_wuser_15_reg(desc_8_wuser_15_reg),
                              .desc_9_txn_type_reg(desc_9_txn_type_reg),
                              .desc_9_size_reg  (desc_9_size_reg),
                              .desc_9_data_offset_reg(desc_9_data_offset_reg),
                              .desc_9_data_host_addr_0_reg(desc_9_data_host_addr_0_reg),
                              .desc_9_data_host_addr_1_reg(desc_9_data_host_addr_1_reg),
                              .desc_9_data_host_addr_2_reg(desc_9_data_host_addr_2_reg),
                              .desc_9_data_host_addr_3_reg(desc_9_data_host_addr_3_reg),
                              .desc_9_wstrb_host_addr_0_reg(desc_9_wstrb_host_addr_0_reg),
                              .desc_9_wstrb_host_addr_1_reg(desc_9_wstrb_host_addr_1_reg),
                              .desc_9_wstrb_host_addr_2_reg(desc_9_wstrb_host_addr_2_reg),
                              .desc_9_wstrb_host_addr_3_reg(desc_9_wstrb_host_addr_3_reg),
                              .desc_9_axsize_reg(desc_9_axsize_reg),
                              .desc_9_attr_reg  (desc_9_attr_reg),
                              .desc_9_axaddr_0_reg(desc_9_axaddr_0_reg),
                              .desc_9_axaddr_1_reg(desc_9_axaddr_1_reg),
                              .desc_9_axaddr_2_reg(desc_9_axaddr_2_reg),
                              .desc_9_axaddr_3_reg(desc_9_axaddr_3_reg),
                              .desc_9_axid_0_reg(desc_9_axid_0_reg),
                              .desc_9_axid_1_reg(desc_9_axid_1_reg),
                              .desc_9_axid_2_reg(desc_9_axid_2_reg),
                              .desc_9_axid_3_reg(desc_9_axid_3_reg),
                              .desc_9_axuser_0_reg(desc_9_axuser_0_reg),
                              .desc_9_axuser_1_reg(desc_9_axuser_1_reg),
                              .desc_9_axuser_2_reg(desc_9_axuser_2_reg),
                              .desc_9_axuser_3_reg(desc_9_axuser_3_reg),
                              .desc_9_axuser_4_reg(desc_9_axuser_4_reg),
                              .desc_9_axuser_5_reg(desc_9_axuser_5_reg),
                              .desc_9_axuser_6_reg(desc_9_axuser_6_reg),
                              .desc_9_axuser_7_reg(desc_9_axuser_7_reg),
                              .desc_9_axuser_8_reg(desc_9_axuser_8_reg),
                              .desc_9_axuser_9_reg(desc_9_axuser_9_reg),
                              .desc_9_axuser_10_reg(desc_9_axuser_10_reg),
                              .desc_9_axuser_11_reg(desc_9_axuser_11_reg),
                              .desc_9_axuser_12_reg(desc_9_axuser_12_reg),
                              .desc_9_axuser_13_reg(desc_9_axuser_13_reg),
                              .desc_9_axuser_14_reg(desc_9_axuser_14_reg),
                              .desc_9_axuser_15_reg(desc_9_axuser_15_reg),
                              .desc_9_xuser_0_reg(desc_9_xuser_0_reg),
                              .desc_9_xuser_1_reg(desc_9_xuser_1_reg),
                              .desc_9_xuser_2_reg(desc_9_xuser_2_reg),
                              .desc_9_xuser_3_reg(desc_9_xuser_3_reg),
                              .desc_9_xuser_4_reg(desc_9_xuser_4_reg),
                              .desc_9_xuser_5_reg(desc_9_xuser_5_reg),
                              .desc_9_xuser_6_reg(desc_9_xuser_6_reg),
                              .desc_9_xuser_7_reg(desc_9_xuser_7_reg),
                              .desc_9_xuser_8_reg(desc_9_xuser_8_reg),
                              .desc_9_xuser_9_reg(desc_9_xuser_9_reg),
                              .desc_9_xuser_10_reg(desc_9_xuser_10_reg),
                              .desc_9_xuser_11_reg(desc_9_xuser_11_reg),
                              .desc_9_xuser_12_reg(desc_9_xuser_12_reg),
                              .desc_9_xuser_13_reg(desc_9_xuser_13_reg),
                              .desc_9_xuser_14_reg(desc_9_xuser_14_reg),
                              .desc_9_xuser_15_reg(desc_9_xuser_15_reg),
                              .desc_9_wuser_0_reg(desc_9_wuser_0_reg),
                              .desc_9_wuser_1_reg(desc_9_wuser_1_reg),
                              .desc_9_wuser_2_reg(desc_9_wuser_2_reg),
                              .desc_9_wuser_3_reg(desc_9_wuser_3_reg),
                              .desc_9_wuser_4_reg(desc_9_wuser_4_reg),
                              .desc_9_wuser_5_reg(desc_9_wuser_5_reg),
                              .desc_9_wuser_6_reg(desc_9_wuser_6_reg),
                              .desc_9_wuser_7_reg(desc_9_wuser_7_reg),
                              .desc_9_wuser_8_reg(desc_9_wuser_8_reg),
                              .desc_9_wuser_9_reg(desc_9_wuser_9_reg),
                              .desc_9_wuser_10_reg(desc_9_wuser_10_reg),
                              .desc_9_wuser_11_reg(desc_9_wuser_11_reg),
                              .desc_9_wuser_12_reg(desc_9_wuser_12_reg),
                              .desc_9_wuser_13_reg(desc_9_wuser_13_reg),
                              .desc_9_wuser_14_reg(desc_9_wuser_14_reg),
                              .desc_9_wuser_15_reg(desc_9_wuser_15_reg),
                              .desc_10_txn_type_reg(desc_10_txn_type_reg),
                              .desc_10_size_reg (desc_10_size_reg),
                              .desc_10_data_offset_reg(desc_10_data_offset_reg),
                              .desc_10_data_host_addr_0_reg(desc_10_data_host_addr_0_reg),
                              .desc_10_data_host_addr_1_reg(desc_10_data_host_addr_1_reg),
                              .desc_10_data_host_addr_2_reg(desc_10_data_host_addr_2_reg),
                              .desc_10_data_host_addr_3_reg(desc_10_data_host_addr_3_reg),
                              .desc_10_wstrb_host_addr_0_reg(desc_10_wstrb_host_addr_0_reg),
                              .desc_10_wstrb_host_addr_1_reg(desc_10_wstrb_host_addr_1_reg),
                              .desc_10_wstrb_host_addr_2_reg(desc_10_wstrb_host_addr_2_reg),
                              .desc_10_wstrb_host_addr_3_reg(desc_10_wstrb_host_addr_3_reg),
                              .desc_10_axsize_reg(desc_10_axsize_reg),
                              .desc_10_attr_reg (desc_10_attr_reg),
                              .desc_10_axaddr_0_reg(desc_10_axaddr_0_reg),
                              .desc_10_axaddr_1_reg(desc_10_axaddr_1_reg),
                              .desc_10_axaddr_2_reg(desc_10_axaddr_2_reg),
                              .desc_10_axaddr_3_reg(desc_10_axaddr_3_reg),
                              .desc_10_axid_0_reg(desc_10_axid_0_reg),
                              .desc_10_axid_1_reg(desc_10_axid_1_reg),
                              .desc_10_axid_2_reg(desc_10_axid_2_reg),
                              .desc_10_axid_3_reg(desc_10_axid_3_reg),
                              .desc_10_axuser_0_reg(desc_10_axuser_0_reg),
                              .desc_10_axuser_1_reg(desc_10_axuser_1_reg),
                              .desc_10_axuser_2_reg(desc_10_axuser_2_reg),
                              .desc_10_axuser_3_reg(desc_10_axuser_3_reg),
                              .desc_10_axuser_4_reg(desc_10_axuser_4_reg),
                              .desc_10_axuser_5_reg(desc_10_axuser_5_reg),
                              .desc_10_axuser_6_reg(desc_10_axuser_6_reg),
                              .desc_10_axuser_7_reg(desc_10_axuser_7_reg),
                              .desc_10_axuser_8_reg(desc_10_axuser_8_reg),
                              .desc_10_axuser_9_reg(desc_10_axuser_9_reg),
                              .desc_10_axuser_10_reg(desc_10_axuser_10_reg),
                              .desc_10_axuser_11_reg(desc_10_axuser_11_reg),
                              .desc_10_axuser_12_reg(desc_10_axuser_12_reg),
                              .desc_10_axuser_13_reg(desc_10_axuser_13_reg),
                              .desc_10_axuser_14_reg(desc_10_axuser_14_reg),
                              .desc_10_axuser_15_reg(desc_10_axuser_15_reg),
                              .desc_10_xuser_0_reg(desc_10_xuser_0_reg),
                              .desc_10_xuser_1_reg(desc_10_xuser_1_reg),
                              .desc_10_xuser_2_reg(desc_10_xuser_2_reg),
                              .desc_10_xuser_3_reg(desc_10_xuser_3_reg),
                              .desc_10_xuser_4_reg(desc_10_xuser_4_reg),
                              .desc_10_xuser_5_reg(desc_10_xuser_5_reg),
                              .desc_10_xuser_6_reg(desc_10_xuser_6_reg),
                              .desc_10_xuser_7_reg(desc_10_xuser_7_reg),
                              .desc_10_xuser_8_reg(desc_10_xuser_8_reg),
                              .desc_10_xuser_9_reg(desc_10_xuser_9_reg),
                              .desc_10_xuser_10_reg(desc_10_xuser_10_reg),
                              .desc_10_xuser_11_reg(desc_10_xuser_11_reg),
                              .desc_10_xuser_12_reg(desc_10_xuser_12_reg),
                              .desc_10_xuser_13_reg(desc_10_xuser_13_reg),
                              .desc_10_xuser_14_reg(desc_10_xuser_14_reg),
                              .desc_10_xuser_15_reg(desc_10_xuser_15_reg),
                              .desc_10_wuser_0_reg(desc_10_wuser_0_reg),
                              .desc_10_wuser_1_reg(desc_10_wuser_1_reg),
                              .desc_10_wuser_2_reg(desc_10_wuser_2_reg),
                              .desc_10_wuser_3_reg(desc_10_wuser_3_reg),
                              .desc_10_wuser_4_reg(desc_10_wuser_4_reg),
                              .desc_10_wuser_5_reg(desc_10_wuser_5_reg),
                              .desc_10_wuser_6_reg(desc_10_wuser_6_reg),
                              .desc_10_wuser_7_reg(desc_10_wuser_7_reg),
                              .desc_10_wuser_8_reg(desc_10_wuser_8_reg),
                              .desc_10_wuser_9_reg(desc_10_wuser_9_reg),
                              .desc_10_wuser_10_reg(desc_10_wuser_10_reg),
                              .desc_10_wuser_11_reg(desc_10_wuser_11_reg),
                              .desc_10_wuser_12_reg(desc_10_wuser_12_reg),
                              .desc_10_wuser_13_reg(desc_10_wuser_13_reg),
                              .desc_10_wuser_14_reg(desc_10_wuser_14_reg),
                              .desc_10_wuser_15_reg(desc_10_wuser_15_reg),
                              .desc_11_txn_type_reg(desc_11_txn_type_reg),
                              .desc_11_size_reg (desc_11_size_reg),
                              .desc_11_data_offset_reg(desc_11_data_offset_reg),
                              .desc_11_data_host_addr_0_reg(desc_11_data_host_addr_0_reg),
                              .desc_11_data_host_addr_1_reg(desc_11_data_host_addr_1_reg),
                              .desc_11_data_host_addr_2_reg(desc_11_data_host_addr_2_reg),
                              .desc_11_data_host_addr_3_reg(desc_11_data_host_addr_3_reg),
                              .desc_11_wstrb_host_addr_0_reg(desc_11_wstrb_host_addr_0_reg),
                              .desc_11_wstrb_host_addr_1_reg(desc_11_wstrb_host_addr_1_reg),
                              .desc_11_wstrb_host_addr_2_reg(desc_11_wstrb_host_addr_2_reg),
                              .desc_11_wstrb_host_addr_3_reg(desc_11_wstrb_host_addr_3_reg),
                              .desc_11_axsize_reg(desc_11_axsize_reg),
                              .desc_11_attr_reg (desc_11_attr_reg),
                              .desc_11_axaddr_0_reg(desc_11_axaddr_0_reg),
                              .desc_11_axaddr_1_reg(desc_11_axaddr_1_reg),
                              .desc_11_axaddr_2_reg(desc_11_axaddr_2_reg),
                              .desc_11_axaddr_3_reg(desc_11_axaddr_3_reg),
                              .desc_11_axid_0_reg(desc_11_axid_0_reg),
                              .desc_11_axid_1_reg(desc_11_axid_1_reg),
                              .desc_11_axid_2_reg(desc_11_axid_2_reg),
                              .desc_11_axid_3_reg(desc_11_axid_3_reg),
                              .desc_11_axuser_0_reg(desc_11_axuser_0_reg),
                              .desc_11_axuser_1_reg(desc_11_axuser_1_reg),
                              .desc_11_axuser_2_reg(desc_11_axuser_2_reg),
                              .desc_11_axuser_3_reg(desc_11_axuser_3_reg),
                              .desc_11_axuser_4_reg(desc_11_axuser_4_reg),
                              .desc_11_axuser_5_reg(desc_11_axuser_5_reg),
                              .desc_11_axuser_6_reg(desc_11_axuser_6_reg),
                              .desc_11_axuser_7_reg(desc_11_axuser_7_reg),
                              .desc_11_axuser_8_reg(desc_11_axuser_8_reg),
                              .desc_11_axuser_9_reg(desc_11_axuser_9_reg),
                              .desc_11_axuser_10_reg(desc_11_axuser_10_reg),
                              .desc_11_axuser_11_reg(desc_11_axuser_11_reg),
                              .desc_11_axuser_12_reg(desc_11_axuser_12_reg),
                              .desc_11_axuser_13_reg(desc_11_axuser_13_reg),
                              .desc_11_axuser_14_reg(desc_11_axuser_14_reg),
                              .desc_11_axuser_15_reg(desc_11_axuser_15_reg),
                              .desc_11_xuser_0_reg(desc_11_xuser_0_reg),
                              .desc_11_xuser_1_reg(desc_11_xuser_1_reg),
                              .desc_11_xuser_2_reg(desc_11_xuser_2_reg),
                              .desc_11_xuser_3_reg(desc_11_xuser_3_reg),
                              .desc_11_xuser_4_reg(desc_11_xuser_4_reg),
                              .desc_11_xuser_5_reg(desc_11_xuser_5_reg),
                              .desc_11_xuser_6_reg(desc_11_xuser_6_reg),
                              .desc_11_xuser_7_reg(desc_11_xuser_7_reg),
                              .desc_11_xuser_8_reg(desc_11_xuser_8_reg),
                              .desc_11_xuser_9_reg(desc_11_xuser_9_reg),
                              .desc_11_xuser_10_reg(desc_11_xuser_10_reg),
                              .desc_11_xuser_11_reg(desc_11_xuser_11_reg),
                              .desc_11_xuser_12_reg(desc_11_xuser_12_reg),
                              .desc_11_xuser_13_reg(desc_11_xuser_13_reg),
                              .desc_11_xuser_14_reg(desc_11_xuser_14_reg),
                              .desc_11_xuser_15_reg(desc_11_xuser_15_reg),
                              .desc_11_wuser_0_reg(desc_11_wuser_0_reg),
                              .desc_11_wuser_1_reg(desc_11_wuser_1_reg),
                              .desc_11_wuser_2_reg(desc_11_wuser_2_reg),
                              .desc_11_wuser_3_reg(desc_11_wuser_3_reg),
                              .desc_11_wuser_4_reg(desc_11_wuser_4_reg),
                              .desc_11_wuser_5_reg(desc_11_wuser_5_reg),
                              .desc_11_wuser_6_reg(desc_11_wuser_6_reg),
                              .desc_11_wuser_7_reg(desc_11_wuser_7_reg),
                              .desc_11_wuser_8_reg(desc_11_wuser_8_reg),
                              .desc_11_wuser_9_reg(desc_11_wuser_9_reg),
                              .desc_11_wuser_10_reg(desc_11_wuser_10_reg),
                              .desc_11_wuser_11_reg(desc_11_wuser_11_reg),
                              .desc_11_wuser_12_reg(desc_11_wuser_12_reg),
                              .desc_11_wuser_13_reg(desc_11_wuser_13_reg),
                              .desc_11_wuser_14_reg(desc_11_wuser_14_reg),
                              .desc_11_wuser_15_reg(desc_11_wuser_15_reg),
                              .desc_12_txn_type_reg(desc_12_txn_type_reg),
                              .desc_12_size_reg (desc_12_size_reg),
                              .desc_12_data_offset_reg(desc_12_data_offset_reg),
                              .desc_12_data_host_addr_0_reg(desc_12_data_host_addr_0_reg),
                              .desc_12_data_host_addr_1_reg(desc_12_data_host_addr_1_reg),
                              .desc_12_data_host_addr_2_reg(desc_12_data_host_addr_2_reg),
                              .desc_12_data_host_addr_3_reg(desc_12_data_host_addr_3_reg),
                              .desc_12_wstrb_host_addr_0_reg(desc_12_wstrb_host_addr_0_reg),
                              .desc_12_wstrb_host_addr_1_reg(desc_12_wstrb_host_addr_1_reg),
                              .desc_12_wstrb_host_addr_2_reg(desc_12_wstrb_host_addr_2_reg),
                              .desc_12_wstrb_host_addr_3_reg(desc_12_wstrb_host_addr_3_reg),
                              .desc_12_axsize_reg(desc_12_axsize_reg),
                              .desc_12_attr_reg (desc_12_attr_reg),
                              .desc_12_axaddr_0_reg(desc_12_axaddr_0_reg),
                              .desc_12_axaddr_1_reg(desc_12_axaddr_1_reg),
                              .desc_12_axaddr_2_reg(desc_12_axaddr_2_reg),
                              .desc_12_axaddr_3_reg(desc_12_axaddr_3_reg),
                              .desc_12_axid_0_reg(desc_12_axid_0_reg),
                              .desc_12_axid_1_reg(desc_12_axid_1_reg),
                              .desc_12_axid_2_reg(desc_12_axid_2_reg),
                              .desc_12_axid_3_reg(desc_12_axid_3_reg),
                              .desc_12_axuser_0_reg(desc_12_axuser_0_reg),
                              .desc_12_axuser_1_reg(desc_12_axuser_1_reg),
                              .desc_12_axuser_2_reg(desc_12_axuser_2_reg),
                              .desc_12_axuser_3_reg(desc_12_axuser_3_reg),
                              .desc_12_axuser_4_reg(desc_12_axuser_4_reg),
                              .desc_12_axuser_5_reg(desc_12_axuser_5_reg),
                              .desc_12_axuser_6_reg(desc_12_axuser_6_reg),
                              .desc_12_axuser_7_reg(desc_12_axuser_7_reg),
                              .desc_12_axuser_8_reg(desc_12_axuser_8_reg),
                              .desc_12_axuser_9_reg(desc_12_axuser_9_reg),
                              .desc_12_axuser_10_reg(desc_12_axuser_10_reg),
                              .desc_12_axuser_11_reg(desc_12_axuser_11_reg),
                              .desc_12_axuser_12_reg(desc_12_axuser_12_reg),
                              .desc_12_axuser_13_reg(desc_12_axuser_13_reg),
                              .desc_12_axuser_14_reg(desc_12_axuser_14_reg),
                              .desc_12_axuser_15_reg(desc_12_axuser_15_reg),
                              .desc_12_xuser_0_reg(desc_12_xuser_0_reg),
                              .desc_12_xuser_1_reg(desc_12_xuser_1_reg),
                              .desc_12_xuser_2_reg(desc_12_xuser_2_reg),
                              .desc_12_xuser_3_reg(desc_12_xuser_3_reg),
                              .desc_12_xuser_4_reg(desc_12_xuser_4_reg),
                              .desc_12_xuser_5_reg(desc_12_xuser_5_reg),
                              .desc_12_xuser_6_reg(desc_12_xuser_6_reg),
                              .desc_12_xuser_7_reg(desc_12_xuser_7_reg),
                              .desc_12_xuser_8_reg(desc_12_xuser_8_reg),
                              .desc_12_xuser_9_reg(desc_12_xuser_9_reg),
                              .desc_12_xuser_10_reg(desc_12_xuser_10_reg),
                              .desc_12_xuser_11_reg(desc_12_xuser_11_reg),
                              .desc_12_xuser_12_reg(desc_12_xuser_12_reg),
                              .desc_12_xuser_13_reg(desc_12_xuser_13_reg),
                              .desc_12_xuser_14_reg(desc_12_xuser_14_reg),
                              .desc_12_xuser_15_reg(desc_12_xuser_15_reg),
                              .desc_12_wuser_0_reg(desc_12_wuser_0_reg),
                              .desc_12_wuser_1_reg(desc_12_wuser_1_reg),
                              .desc_12_wuser_2_reg(desc_12_wuser_2_reg),
                              .desc_12_wuser_3_reg(desc_12_wuser_3_reg),
                              .desc_12_wuser_4_reg(desc_12_wuser_4_reg),
                              .desc_12_wuser_5_reg(desc_12_wuser_5_reg),
                              .desc_12_wuser_6_reg(desc_12_wuser_6_reg),
                              .desc_12_wuser_7_reg(desc_12_wuser_7_reg),
                              .desc_12_wuser_8_reg(desc_12_wuser_8_reg),
                              .desc_12_wuser_9_reg(desc_12_wuser_9_reg),
                              .desc_12_wuser_10_reg(desc_12_wuser_10_reg),
                              .desc_12_wuser_11_reg(desc_12_wuser_11_reg),
                              .desc_12_wuser_12_reg(desc_12_wuser_12_reg),
                              .desc_12_wuser_13_reg(desc_12_wuser_13_reg),
                              .desc_12_wuser_14_reg(desc_12_wuser_14_reg),
                              .desc_12_wuser_15_reg(desc_12_wuser_15_reg),
                              .desc_13_txn_type_reg(desc_13_txn_type_reg),
                              .desc_13_size_reg (desc_13_size_reg),
                              .desc_13_data_offset_reg(desc_13_data_offset_reg),
                              .desc_13_data_host_addr_0_reg(desc_13_data_host_addr_0_reg),
                              .desc_13_data_host_addr_1_reg(desc_13_data_host_addr_1_reg),
                              .desc_13_data_host_addr_2_reg(desc_13_data_host_addr_2_reg),
                              .desc_13_data_host_addr_3_reg(desc_13_data_host_addr_3_reg),
                              .desc_13_wstrb_host_addr_0_reg(desc_13_wstrb_host_addr_0_reg),
                              .desc_13_wstrb_host_addr_1_reg(desc_13_wstrb_host_addr_1_reg),
                              .desc_13_wstrb_host_addr_2_reg(desc_13_wstrb_host_addr_2_reg),
                              .desc_13_wstrb_host_addr_3_reg(desc_13_wstrb_host_addr_3_reg),
                              .desc_13_axsize_reg(desc_13_axsize_reg),
                              .desc_13_attr_reg (desc_13_attr_reg),
                              .desc_13_axaddr_0_reg(desc_13_axaddr_0_reg),
                              .desc_13_axaddr_1_reg(desc_13_axaddr_1_reg),
                              .desc_13_axaddr_2_reg(desc_13_axaddr_2_reg),
                              .desc_13_axaddr_3_reg(desc_13_axaddr_3_reg),
                              .desc_13_axid_0_reg(desc_13_axid_0_reg),
                              .desc_13_axid_1_reg(desc_13_axid_1_reg),
                              .desc_13_axid_2_reg(desc_13_axid_2_reg),
                              .desc_13_axid_3_reg(desc_13_axid_3_reg),
                              .desc_13_axuser_0_reg(desc_13_axuser_0_reg),
                              .desc_13_axuser_1_reg(desc_13_axuser_1_reg),
                              .desc_13_axuser_2_reg(desc_13_axuser_2_reg),
                              .desc_13_axuser_3_reg(desc_13_axuser_3_reg),
                              .desc_13_axuser_4_reg(desc_13_axuser_4_reg),
                              .desc_13_axuser_5_reg(desc_13_axuser_5_reg),
                              .desc_13_axuser_6_reg(desc_13_axuser_6_reg),
                              .desc_13_axuser_7_reg(desc_13_axuser_7_reg),
                              .desc_13_axuser_8_reg(desc_13_axuser_8_reg),
                              .desc_13_axuser_9_reg(desc_13_axuser_9_reg),
                              .desc_13_axuser_10_reg(desc_13_axuser_10_reg),
                              .desc_13_axuser_11_reg(desc_13_axuser_11_reg),
                              .desc_13_axuser_12_reg(desc_13_axuser_12_reg),
                              .desc_13_axuser_13_reg(desc_13_axuser_13_reg),
                              .desc_13_axuser_14_reg(desc_13_axuser_14_reg),
                              .desc_13_axuser_15_reg(desc_13_axuser_15_reg),
                              .desc_13_xuser_0_reg(desc_13_xuser_0_reg),
                              .desc_13_xuser_1_reg(desc_13_xuser_1_reg),
                              .desc_13_xuser_2_reg(desc_13_xuser_2_reg),
                              .desc_13_xuser_3_reg(desc_13_xuser_3_reg),
                              .desc_13_xuser_4_reg(desc_13_xuser_4_reg),
                              .desc_13_xuser_5_reg(desc_13_xuser_5_reg),
                              .desc_13_xuser_6_reg(desc_13_xuser_6_reg),
                              .desc_13_xuser_7_reg(desc_13_xuser_7_reg),
                              .desc_13_xuser_8_reg(desc_13_xuser_8_reg),
                              .desc_13_xuser_9_reg(desc_13_xuser_9_reg),
                              .desc_13_xuser_10_reg(desc_13_xuser_10_reg),
                              .desc_13_xuser_11_reg(desc_13_xuser_11_reg),
                              .desc_13_xuser_12_reg(desc_13_xuser_12_reg),
                              .desc_13_xuser_13_reg(desc_13_xuser_13_reg),
                              .desc_13_xuser_14_reg(desc_13_xuser_14_reg),
                              .desc_13_xuser_15_reg(desc_13_xuser_15_reg),
                              .desc_13_wuser_0_reg(desc_13_wuser_0_reg),
                              .desc_13_wuser_1_reg(desc_13_wuser_1_reg),
                              .desc_13_wuser_2_reg(desc_13_wuser_2_reg),
                              .desc_13_wuser_3_reg(desc_13_wuser_3_reg),
                              .desc_13_wuser_4_reg(desc_13_wuser_4_reg),
                              .desc_13_wuser_5_reg(desc_13_wuser_5_reg),
                              .desc_13_wuser_6_reg(desc_13_wuser_6_reg),
                              .desc_13_wuser_7_reg(desc_13_wuser_7_reg),
                              .desc_13_wuser_8_reg(desc_13_wuser_8_reg),
                              .desc_13_wuser_9_reg(desc_13_wuser_9_reg),
                              .desc_13_wuser_10_reg(desc_13_wuser_10_reg),
                              .desc_13_wuser_11_reg(desc_13_wuser_11_reg),
                              .desc_13_wuser_12_reg(desc_13_wuser_12_reg),
                              .desc_13_wuser_13_reg(desc_13_wuser_13_reg),
                              .desc_13_wuser_14_reg(desc_13_wuser_14_reg),
                              .desc_13_wuser_15_reg(desc_13_wuser_15_reg),
                              .desc_14_txn_type_reg(desc_14_txn_type_reg),
                              .desc_14_size_reg (desc_14_size_reg),
                              .desc_14_data_offset_reg(desc_14_data_offset_reg),
                              .desc_14_data_host_addr_0_reg(desc_14_data_host_addr_0_reg),
                              .desc_14_data_host_addr_1_reg(desc_14_data_host_addr_1_reg),
                              .desc_14_data_host_addr_2_reg(desc_14_data_host_addr_2_reg),
                              .desc_14_data_host_addr_3_reg(desc_14_data_host_addr_3_reg),
                              .desc_14_wstrb_host_addr_0_reg(desc_14_wstrb_host_addr_0_reg),
                              .desc_14_wstrb_host_addr_1_reg(desc_14_wstrb_host_addr_1_reg),
                              .desc_14_wstrb_host_addr_2_reg(desc_14_wstrb_host_addr_2_reg),
                              .desc_14_wstrb_host_addr_3_reg(desc_14_wstrb_host_addr_3_reg),
                              .desc_14_axsize_reg(desc_14_axsize_reg),
                              .desc_14_attr_reg (desc_14_attr_reg),
                              .desc_14_axaddr_0_reg(desc_14_axaddr_0_reg),
                              .desc_14_axaddr_1_reg(desc_14_axaddr_1_reg),
                              .desc_14_axaddr_2_reg(desc_14_axaddr_2_reg),
                              .desc_14_axaddr_3_reg(desc_14_axaddr_3_reg),
                              .desc_14_axid_0_reg(desc_14_axid_0_reg),
                              .desc_14_axid_1_reg(desc_14_axid_1_reg),
                              .desc_14_axid_2_reg(desc_14_axid_2_reg),
                              .desc_14_axid_3_reg(desc_14_axid_3_reg),
                              .desc_14_axuser_0_reg(desc_14_axuser_0_reg),
                              .desc_14_axuser_1_reg(desc_14_axuser_1_reg),
                              .desc_14_axuser_2_reg(desc_14_axuser_2_reg),
                              .desc_14_axuser_3_reg(desc_14_axuser_3_reg),
                              .desc_14_axuser_4_reg(desc_14_axuser_4_reg),
                              .desc_14_axuser_5_reg(desc_14_axuser_5_reg),
                              .desc_14_axuser_6_reg(desc_14_axuser_6_reg),
                              .desc_14_axuser_7_reg(desc_14_axuser_7_reg),
                              .desc_14_axuser_8_reg(desc_14_axuser_8_reg),
                              .desc_14_axuser_9_reg(desc_14_axuser_9_reg),
                              .desc_14_axuser_10_reg(desc_14_axuser_10_reg),
                              .desc_14_axuser_11_reg(desc_14_axuser_11_reg),
                              .desc_14_axuser_12_reg(desc_14_axuser_12_reg),
                              .desc_14_axuser_13_reg(desc_14_axuser_13_reg),
                              .desc_14_axuser_14_reg(desc_14_axuser_14_reg),
                              .desc_14_axuser_15_reg(desc_14_axuser_15_reg),
                              .desc_14_xuser_0_reg(desc_14_xuser_0_reg),
                              .desc_14_xuser_1_reg(desc_14_xuser_1_reg),
                              .desc_14_xuser_2_reg(desc_14_xuser_2_reg),
                              .desc_14_xuser_3_reg(desc_14_xuser_3_reg),
                              .desc_14_xuser_4_reg(desc_14_xuser_4_reg),
                              .desc_14_xuser_5_reg(desc_14_xuser_5_reg),
                              .desc_14_xuser_6_reg(desc_14_xuser_6_reg),
                              .desc_14_xuser_7_reg(desc_14_xuser_7_reg),
                              .desc_14_xuser_8_reg(desc_14_xuser_8_reg),
                              .desc_14_xuser_9_reg(desc_14_xuser_9_reg),
                              .desc_14_xuser_10_reg(desc_14_xuser_10_reg),
                              .desc_14_xuser_11_reg(desc_14_xuser_11_reg),
                              .desc_14_xuser_12_reg(desc_14_xuser_12_reg),
                              .desc_14_xuser_13_reg(desc_14_xuser_13_reg),
                              .desc_14_xuser_14_reg(desc_14_xuser_14_reg),
                              .desc_14_xuser_15_reg(desc_14_xuser_15_reg),
                              .desc_14_wuser_0_reg(desc_14_wuser_0_reg),
                              .desc_14_wuser_1_reg(desc_14_wuser_1_reg),
                              .desc_14_wuser_2_reg(desc_14_wuser_2_reg),
                              .desc_14_wuser_3_reg(desc_14_wuser_3_reg),
                              .desc_14_wuser_4_reg(desc_14_wuser_4_reg),
                              .desc_14_wuser_5_reg(desc_14_wuser_5_reg),
                              .desc_14_wuser_6_reg(desc_14_wuser_6_reg),
                              .desc_14_wuser_7_reg(desc_14_wuser_7_reg),
                              .desc_14_wuser_8_reg(desc_14_wuser_8_reg),
                              .desc_14_wuser_9_reg(desc_14_wuser_9_reg),
                              .desc_14_wuser_10_reg(desc_14_wuser_10_reg),
                              .desc_14_wuser_11_reg(desc_14_wuser_11_reg),
                              .desc_14_wuser_12_reg(desc_14_wuser_12_reg),
                              .desc_14_wuser_13_reg(desc_14_wuser_13_reg),
                              .desc_14_wuser_14_reg(desc_14_wuser_14_reg),
                              .desc_14_wuser_15_reg(desc_14_wuser_15_reg),
                              .desc_15_txn_type_reg(desc_15_txn_type_reg),
                              .desc_15_size_reg (desc_15_size_reg),
                              .desc_15_data_offset_reg(desc_15_data_offset_reg),
                              .desc_15_data_host_addr_0_reg(desc_15_data_host_addr_0_reg),
                              .desc_15_data_host_addr_1_reg(desc_15_data_host_addr_1_reg),
                              .desc_15_data_host_addr_2_reg(desc_15_data_host_addr_2_reg),
                              .desc_15_data_host_addr_3_reg(desc_15_data_host_addr_3_reg),
                              .desc_15_wstrb_host_addr_0_reg(desc_15_wstrb_host_addr_0_reg),
                              .desc_15_wstrb_host_addr_1_reg(desc_15_wstrb_host_addr_1_reg),
                              .desc_15_wstrb_host_addr_2_reg(desc_15_wstrb_host_addr_2_reg),
                              .desc_15_wstrb_host_addr_3_reg(desc_15_wstrb_host_addr_3_reg),
                              .desc_15_axsize_reg(desc_15_axsize_reg),
                              .desc_15_attr_reg (desc_15_attr_reg),
                              .desc_15_axaddr_0_reg(desc_15_axaddr_0_reg),
                              .desc_15_axaddr_1_reg(desc_15_axaddr_1_reg),
                              .desc_15_axaddr_2_reg(desc_15_axaddr_2_reg),
                              .desc_15_axaddr_3_reg(desc_15_axaddr_3_reg),
                              .desc_15_axid_0_reg(desc_15_axid_0_reg),
                              .desc_15_axid_1_reg(desc_15_axid_1_reg),
                              .desc_15_axid_2_reg(desc_15_axid_2_reg),
                              .desc_15_axid_3_reg(desc_15_axid_3_reg),
                              .desc_15_axuser_0_reg(desc_15_axuser_0_reg),
                              .desc_15_axuser_1_reg(desc_15_axuser_1_reg),
                              .desc_15_axuser_2_reg(desc_15_axuser_2_reg),
                              .desc_15_axuser_3_reg(desc_15_axuser_3_reg),
                              .desc_15_axuser_4_reg(desc_15_axuser_4_reg),
                              .desc_15_axuser_5_reg(desc_15_axuser_5_reg),
                              .desc_15_axuser_6_reg(desc_15_axuser_6_reg),
                              .desc_15_axuser_7_reg(desc_15_axuser_7_reg),
                              .desc_15_axuser_8_reg(desc_15_axuser_8_reg),
                              .desc_15_axuser_9_reg(desc_15_axuser_9_reg),
                              .desc_15_axuser_10_reg(desc_15_axuser_10_reg),
                              .desc_15_axuser_11_reg(desc_15_axuser_11_reg),
                              .desc_15_axuser_12_reg(desc_15_axuser_12_reg),
                              .desc_15_axuser_13_reg(desc_15_axuser_13_reg),
                              .desc_15_axuser_14_reg(desc_15_axuser_14_reg),
                              .desc_15_axuser_15_reg(desc_15_axuser_15_reg),
                              .desc_15_xuser_0_reg(desc_15_xuser_0_reg),
                              .desc_15_xuser_1_reg(desc_15_xuser_1_reg),
                              .desc_15_xuser_2_reg(desc_15_xuser_2_reg),
                              .desc_15_xuser_3_reg(desc_15_xuser_3_reg),
                              .desc_15_xuser_4_reg(desc_15_xuser_4_reg),
                              .desc_15_xuser_5_reg(desc_15_xuser_5_reg),
                              .desc_15_xuser_6_reg(desc_15_xuser_6_reg),
                              .desc_15_xuser_7_reg(desc_15_xuser_7_reg),
                              .desc_15_xuser_8_reg(desc_15_xuser_8_reg),
                              .desc_15_xuser_9_reg(desc_15_xuser_9_reg),
                              .desc_15_xuser_10_reg(desc_15_xuser_10_reg),
                              .desc_15_xuser_11_reg(desc_15_xuser_11_reg),
                              .desc_15_xuser_12_reg(desc_15_xuser_12_reg),
                              .desc_15_xuser_13_reg(desc_15_xuser_13_reg),
                              .desc_15_xuser_14_reg(desc_15_xuser_14_reg),
                              .desc_15_xuser_15_reg(desc_15_xuser_15_reg),
                              .desc_15_wuser_0_reg(desc_15_wuser_0_reg),
                              .desc_15_wuser_1_reg(desc_15_wuser_1_reg),
                              .desc_15_wuser_2_reg(desc_15_wuser_2_reg),
                              .desc_15_wuser_3_reg(desc_15_wuser_3_reg),
                              .desc_15_wuser_4_reg(desc_15_wuser_4_reg),
                              .desc_15_wuser_5_reg(desc_15_wuser_5_reg),
                              .desc_15_wuser_6_reg(desc_15_wuser_6_reg),
                              .desc_15_wuser_7_reg(desc_15_wuser_7_reg),
                              .desc_15_wuser_8_reg(desc_15_wuser_8_reg),
                              .desc_15_wuser_9_reg(desc_15_wuser_9_reg),
                              .desc_15_wuser_10_reg(desc_15_wuser_10_reg),
                              .desc_15_wuser_11_reg(desc_15_wuser_11_reg),
                              .desc_15_wuser_12_reg(desc_15_wuser_12_reg),
                              .desc_15_wuser_13_reg(desc_15_wuser_13_reg),
                              .desc_15_wuser_14_reg(desc_15_wuser_14_reg),
                              .desc_15_wuser_15_reg(desc_15_wuser_15_reg),
                              // Inputs
                              .hm2rb_intr_error_status_reg_we({31'h0,hm2rb_intr_error_status_reg_we[0]}),
                              .hm2rb_intr_error_status_reg({31'h0,hm2rb_intr_error_status_reg[0]}),
                              .axi_aclk         (axi_aclk),
                              .axi_aresetn      (axi_aresetn),
                              .rst_n            (rst_n),
                              .s_axi_awaddr     (s_axi_awaddr),
                              .s_axi_awprot     (s_axi_awprot),
                              .s_axi_awvalid    (s_axi_awvalid),
                              .s_axi_wdata      (s_axi_wdata),
                              .s_axi_wstrb      (s_axi_wstrb),
                              .s_axi_wvalid     (s_axi_wvalid),
                              .s_axi_bready     (s_axi_bready),
                              .s_axi_araddr     (s_axi_araddr),
                              .s_axi_arprot     (s_axi_arprot),
                              .s_axi_arvalid    (s_axi_arvalid),
                              .s_axi_rready     (s_axi_rready),
                              .rb2uc_rd_data    (rb2uc_rd_data),
                              .hm2rb_rd_addr    (hm2rb_rd_addr),
                              .hm2rb_wr_we      (hm2rb_wr_we),
                              .hm2rb_wr_bwe     (hm2rb_wr_bwe),
                              .hm2rb_wr_addr    (hm2rb_wr_addr),
                              .hm2rb_wr_data    (hm2rb_wr_data),
                              .hm2uc_done       (hm2uc_done),
                              .uc2rb_intr_error_status_reg(uc2rb_intr_error_status_reg),
                              .uc2rb_ownership_reg(uc2rb_ownership_reg),
                              .uc2rb_intr_txn_avail_status_reg(uc2rb_intr_txn_avail_status_reg),
                              .uc2rb_intr_comp_status_reg(uc2rb_intr_comp_status_reg),
                              .uc2rb_status_busy_reg(uc2rb_status_busy_reg),
                              .uc2rb_resp_fifo_free_level_reg(uc2rb_resp_fifo_free_level_reg),
                              .uc2rb_desc_0_txn_type_reg(uc2rb_desc_0_txn_type_reg),
                              .uc2rb_desc_0_size_reg(uc2rb_desc_0_size_reg),
                              .uc2rb_desc_0_data_offset_reg(uc2rb_desc_0_data_offset_reg),
                              .uc2rb_desc_0_axsize_reg(uc2rb_desc_0_axsize_reg),
                              .uc2rb_desc_0_attr_reg(uc2rb_desc_0_attr_reg),
                              .uc2rb_desc_0_axaddr_0_reg(uc2rb_desc_0_axaddr_0_reg),
                              .uc2rb_desc_0_axaddr_1_reg(uc2rb_desc_0_axaddr_1_reg),
                              .uc2rb_desc_0_axaddr_2_reg(uc2rb_desc_0_axaddr_2_reg),
                              .uc2rb_desc_0_axaddr_3_reg(uc2rb_desc_0_axaddr_3_reg),
                              .uc2rb_desc_0_axid_0_reg(uc2rb_desc_0_axid_0_reg),
                              .uc2rb_desc_0_axid_1_reg(uc2rb_desc_0_axid_1_reg),
                              .uc2rb_desc_0_axid_2_reg(uc2rb_desc_0_axid_2_reg),
                              .uc2rb_desc_0_axid_3_reg(uc2rb_desc_0_axid_3_reg),
                              .uc2rb_desc_0_axuser_0_reg(uc2rb_desc_0_axuser_0_reg),
                              .uc2rb_desc_0_axuser_1_reg(uc2rb_desc_0_axuser_1_reg),
                              .uc2rb_desc_0_axuser_2_reg(uc2rb_desc_0_axuser_2_reg),
                              .uc2rb_desc_0_axuser_3_reg(uc2rb_desc_0_axuser_3_reg),
                              .uc2rb_desc_0_axuser_4_reg(uc2rb_desc_0_axuser_4_reg),
                              .uc2rb_desc_0_axuser_5_reg(uc2rb_desc_0_axuser_5_reg),
                              .uc2rb_desc_0_axuser_6_reg(uc2rb_desc_0_axuser_6_reg),
                              .uc2rb_desc_0_axuser_7_reg(uc2rb_desc_0_axuser_7_reg),
                              .uc2rb_desc_0_axuser_8_reg(uc2rb_desc_0_axuser_8_reg),
                              .uc2rb_desc_0_axuser_9_reg(uc2rb_desc_0_axuser_9_reg),
                              .uc2rb_desc_0_axuser_10_reg(uc2rb_desc_0_axuser_10_reg),
                              .uc2rb_desc_0_axuser_11_reg(uc2rb_desc_0_axuser_11_reg),
                              .uc2rb_desc_0_axuser_12_reg(uc2rb_desc_0_axuser_12_reg),
                              .uc2rb_desc_0_axuser_13_reg(uc2rb_desc_0_axuser_13_reg),
                              .uc2rb_desc_0_axuser_14_reg(uc2rb_desc_0_axuser_14_reg),
                              .uc2rb_desc_0_axuser_15_reg(uc2rb_desc_0_axuser_15_reg),
                              .uc2rb_desc_0_wuser_0_reg(uc2rb_desc_0_wuser_0_reg),
                              .uc2rb_desc_0_wuser_1_reg(uc2rb_desc_0_wuser_1_reg),
                              .uc2rb_desc_0_wuser_2_reg(uc2rb_desc_0_wuser_2_reg),
                              .uc2rb_desc_0_wuser_3_reg(uc2rb_desc_0_wuser_3_reg),
                              .uc2rb_desc_0_wuser_4_reg(uc2rb_desc_0_wuser_4_reg),
                              .uc2rb_desc_0_wuser_5_reg(uc2rb_desc_0_wuser_5_reg),
                              .uc2rb_desc_0_wuser_6_reg(uc2rb_desc_0_wuser_6_reg),
                              .uc2rb_desc_0_wuser_7_reg(uc2rb_desc_0_wuser_7_reg),
                              .uc2rb_desc_0_wuser_8_reg(uc2rb_desc_0_wuser_8_reg),
                              .uc2rb_desc_0_wuser_9_reg(uc2rb_desc_0_wuser_9_reg),
                              .uc2rb_desc_0_wuser_10_reg(uc2rb_desc_0_wuser_10_reg),
                              .uc2rb_desc_0_wuser_11_reg(uc2rb_desc_0_wuser_11_reg),
                              .uc2rb_desc_0_wuser_12_reg(uc2rb_desc_0_wuser_12_reg),
                              .uc2rb_desc_0_wuser_13_reg(uc2rb_desc_0_wuser_13_reg),
                              .uc2rb_desc_0_wuser_14_reg(uc2rb_desc_0_wuser_14_reg),
                              .uc2rb_desc_0_wuser_15_reg(uc2rb_desc_0_wuser_15_reg),
                              .uc2rb_desc_1_txn_type_reg(uc2rb_desc_1_txn_type_reg),
                              .uc2rb_desc_1_size_reg(uc2rb_desc_1_size_reg),
                              .uc2rb_desc_1_data_offset_reg(uc2rb_desc_1_data_offset_reg),
                              .uc2rb_desc_1_axsize_reg(uc2rb_desc_1_axsize_reg),
                              .uc2rb_desc_1_attr_reg(uc2rb_desc_1_attr_reg),
                              .uc2rb_desc_1_axaddr_0_reg(uc2rb_desc_1_axaddr_0_reg),
                              .uc2rb_desc_1_axaddr_1_reg(uc2rb_desc_1_axaddr_1_reg),
                              .uc2rb_desc_1_axaddr_2_reg(uc2rb_desc_1_axaddr_2_reg),
                              .uc2rb_desc_1_axaddr_3_reg(uc2rb_desc_1_axaddr_3_reg),
                              .uc2rb_desc_1_axid_0_reg(uc2rb_desc_1_axid_0_reg),
                              .uc2rb_desc_1_axid_1_reg(uc2rb_desc_1_axid_1_reg),
                              .uc2rb_desc_1_axid_2_reg(uc2rb_desc_1_axid_2_reg),
                              .uc2rb_desc_1_axid_3_reg(uc2rb_desc_1_axid_3_reg),
                              .uc2rb_desc_1_axuser_0_reg(uc2rb_desc_1_axuser_0_reg),
                              .uc2rb_desc_1_axuser_1_reg(uc2rb_desc_1_axuser_1_reg),
                              .uc2rb_desc_1_axuser_2_reg(uc2rb_desc_1_axuser_2_reg),
                              .uc2rb_desc_1_axuser_3_reg(uc2rb_desc_1_axuser_3_reg),
                              .uc2rb_desc_1_axuser_4_reg(uc2rb_desc_1_axuser_4_reg),
                              .uc2rb_desc_1_axuser_5_reg(uc2rb_desc_1_axuser_5_reg),
                              .uc2rb_desc_1_axuser_6_reg(uc2rb_desc_1_axuser_6_reg),
                              .uc2rb_desc_1_axuser_7_reg(uc2rb_desc_1_axuser_7_reg),
                              .uc2rb_desc_1_axuser_8_reg(uc2rb_desc_1_axuser_8_reg),
                              .uc2rb_desc_1_axuser_9_reg(uc2rb_desc_1_axuser_9_reg),
                              .uc2rb_desc_1_axuser_10_reg(uc2rb_desc_1_axuser_10_reg),
                              .uc2rb_desc_1_axuser_11_reg(uc2rb_desc_1_axuser_11_reg),
                              .uc2rb_desc_1_axuser_12_reg(uc2rb_desc_1_axuser_12_reg),
                              .uc2rb_desc_1_axuser_13_reg(uc2rb_desc_1_axuser_13_reg),
                              .uc2rb_desc_1_axuser_14_reg(uc2rb_desc_1_axuser_14_reg),
                              .uc2rb_desc_1_axuser_15_reg(uc2rb_desc_1_axuser_15_reg),
                              .uc2rb_desc_1_wuser_0_reg(uc2rb_desc_1_wuser_0_reg),
                              .uc2rb_desc_1_wuser_1_reg(uc2rb_desc_1_wuser_1_reg),
                              .uc2rb_desc_1_wuser_2_reg(uc2rb_desc_1_wuser_2_reg),
                              .uc2rb_desc_1_wuser_3_reg(uc2rb_desc_1_wuser_3_reg),
                              .uc2rb_desc_1_wuser_4_reg(uc2rb_desc_1_wuser_4_reg),
                              .uc2rb_desc_1_wuser_5_reg(uc2rb_desc_1_wuser_5_reg),
                              .uc2rb_desc_1_wuser_6_reg(uc2rb_desc_1_wuser_6_reg),
                              .uc2rb_desc_1_wuser_7_reg(uc2rb_desc_1_wuser_7_reg),
                              .uc2rb_desc_1_wuser_8_reg(uc2rb_desc_1_wuser_8_reg),
                              .uc2rb_desc_1_wuser_9_reg(uc2rb_desc_1_wuser_9_reg),
                              .uc2rb_desc_1_wuser_10_reg(uc2rb_desc_1_wuser_10_reg),
                              .uc2rb_desc_1_wuser_11_reg(uc2rb_desc_1_wuser_11_reg),
                              .uc2rb_desc_1_wuser_12_reg(uc2rb_desc_1_wuser_12_reg),
                              .uc2rb_desc_1_wuser_13_reg(uc2rb_desc_1_wuser_13_reg),
                              .uc2rb_desc_1_wuser_14_reg(uc2rb_desc_1_wuser_14_reg),
                              .uc2rb_desc_1_wuser_15_reg(uc2rb_desc_1_wuser_15_reg),
                              .uc2rb_desc_2_txn_type_reg(uc2rb_desc_2_txn_type_reg),
                              .uc2rb_desc_2_size_reg(uc2rb_desc_2_size_reg),
                              .uc2rb_desc_2_data_offset_reg(uc2rb_desc_2_data_offset_reg),
                              .uc2rb_desc_2_axsize_reg(uc2rb_desc_2_axsize_reg),
                              .uc2rb_desc_2_attr_reg(uc2rb_desc_2_attr_reg),
                              .uc2rb_desc_2_axaddr_0_reg(uc2rb_desc_2_axaddr_0_reg),
                              .uc2rb_desc_2_axaddr_1_reg(uc2rb_desc_2_axaddr_1_reg),
                              .uc2rb_desc_2_axaddr_2_reg(uc2rb_desc_2_axaddr_2_reg),
                              .uc2rb_desc_2_axaddr_3_reg(uc2rb_desc_2_axaddr_3_reg),
                              .uc2rb_desc_2_axid_0_reg(uc2rb_desc_2_axid_0_reg),
                              .uc2rb_desc_2_axid_1_reg(uc2rb_desc_2_axid_1_reg),
                              .uc2rb_desc_2_axid_2_reg(uc2rb_desc_2_axid_2_reg),
                              .uc2rb_desc_2_axid_3_reg(uc2rb_desc_2_axid_3_reg),
                              .uc2rb_desc_2_axuser_0_reg(uc2rb_desc_2_axuser_0_reg),
                              .uc2rb_desc_2_axuser_1_reg(uc2rb_desc_2_axuser_1_reg),
                              .uc2rb_desc_2_axuser_2_reg(uc2rb_desc_2_axuser_2_reg),
                              .uc2rb_desc_2_axuser_3_reg(uc2rb_desc_2_axuser_3_reg),
                              .uc2rb_desc_2_axuser_4_reg(uc2rb_desc_2_axuser_4_reg),
                              .uc2rb_desc_2_axuser_5_reg(uc2rb_desc_2_axuser_5_reg),
                              .uc2rb_desc_2_axuser_6_reg(uc2rb_desc_2_axuser_6_reg),
                              .uc2rb_desc_2_axuser_7_reg(uc2rb_desc_2_axuser_7_reg),
                              .uc2rb_desc_2_axuser_8_reg(uc2rb_desc_2_axuser_8_reg),
                              .uc2rb_desc_2_axuser_9_reg(uc2rb_desc_2_axuser_9_reg),
                              .uc2rb_desc_2_axuser_10_reg(uc2rb_desc_2_axuser_10_reg),
                              .uc2rb_desc_2_axuser_11_reg(uc2rb_desc_2_axuser_11_reg),
                              .uc2rb_desc_2_axuser_12_reg(uc2rb_desc_2_axuser_12_reg),
                              .uc2rb_desc_2_axuser_13_reg(uc2rb_desc_2_axuser_13_reg),
                              .uc2rb_desc_2_axuser_14_reg(uc2rb_desc_2_axuser_14_reg),
                              .uc2rb_desc_2_axuser_15_reg(uc2rb_desc_2_axuser_15_reg),
                              .uc2rb_desc_2_wuser_0_reg(uc2rb_desc_2_wuser_0_reg),
                              .uc2rb_desc_2_wuser_1_reg(uc2rb_desc_2_wuser_1_reg),
                              .uc2rb_desc_2_wuser_2_reg(uc2rb_desc_2_wuser_2_reg),
                              .uc2rb_desc_2_wuser_3_reg(uc2rb_desc_2_wuser_3_reg),
                              .uc2rb_desc_2_wuser_4_reg(uc2rb_desc_2_wuser_4_reg),
                              .uc2rb_desc_2_wuser_5_reg(uc2rb_desc_2_wuser_5_reg),
                              .uc2rb_desc_2_wuser_6_reg(uc2rb_desc_2_wuser_6_reg),
                              .uc2rb_desc_2_wuser_7_reg(uc2rb_desc_2_wuser_7_reg),
                              .uc2rb_desc_2_wuser_8_reg(uc2rb_desc_2_wuser_8_reg),
                              .uc2rb_desc_2_wuser_9_reg(uc2rb_desc_2_wuser_9_reg),
                              .uc2rb_desc_2_wuser_10_reg(uc2rb_desc_2_wuser_10_reg),
                              .uc2rb_desc_2_wuser_11_reg(uc2rb_desc_2_wuser_11_reg),
                              .uc2rb_desc_2_wuser_12_reg(uc2rb_desc_2_wuser_12_reg),
                              .uc2rb_desc_2_wuser_13_reg(uc2rb_desc_2_wuser_13_reg),
                              .uc2rb_desc_2_wuser_14_reg(uc2rb_desc_2_wuser_14_reg),
                              .uc2rb_desc_2_wuser_15_reg(uc2rb_desc_2_wuser_15_reg),
                              .uc2rb_desc_3_txn_type_reg(uc2rb_desc_3_txn_type_reg),
                              .uc2rb_desc_3_size_reg(uc2rb_desc_3_size_reg),
                              .uc2rb_desc_3_data_offset_reg(uc2rb_desc_3_data_offset_reg),
                              .uc2rb_desc_3_axsize_reg(uc2rb_desc_3_axsize_reg),
                              .uc2rb_desc_3_attr_reg(uc2rb_desc_3_attr_reg),
                              .uc2rb_desc_3_axaddr_0_reg(uc2rb_desc_3_axaddr_0_reg),
                              .uc2rb_desc_3_axaddr_1_reg(uc2rb_desc_3_axaddr_1_reg),
                              .uc2rb_desc_3_axaddr_2_reg(uc2rb_desc_3_axaddr_2_reg),
                              .uc2rb_desc_3_axaddr_3_reg(uc2rb_desc_3_axaddr_3_reg),
                              .uc2rb_desc_3_axid_0_reg(uc2rb_desc_3_axid_0_reg),
                              .uc2rb_desc_3_axid_1_reg(uc2rb_desc_3_axid_1_reg),
                              .uc2rb_desc_3_axid_2_reg(uc2rb_desc_3_axid_2_reg),
                              .uc2rb_desc_3_axid_3_reg(uc2rb_desc_3_axid_3_reg),
                              .uc2rb_desc_3_axuser_0_reg(uc2rb_desc_3_axuser_0_reg),
                              .uc2rb_desc_3_axuser_1_reg(uc2rb_desc_3_axuser_1_reg),
                              .uc2rb_desc_3_axuser_2_reg(uc2rb_desc_3_axuser_2_reg),
                              .uc2rb_desc_3_axuser_3_reg(uc2rb_desc_3_axuser_3_reg),
                              .uc2rb_desc_3_axuser_4_reg(uc2rb_desc_3_axuser_4_reg),
                              .uc2rb_desc_3_axuser_5_reg(uc2rb_desc_3_axuser_5_reg),
                              .uc2rb_desc_3_axuser_6_reg(uc2rb_desc_3_axuser_6_reg),
                              .uc2rb_desc_3_axuser_7_reg(uc2rb_desc_3_axuser_7_reg),
                              .uc2rb_desc_3_axuser_8_reg(uc2rb_desc_3_axuser_8_reg),
                              .uc2rb_desc_3_axuser_9_reg(uc2rb_desc_3_axuser_9_reg),
                              .uc2rb_desc_3_axuser_10_reg(uc2rb_desc_3_axuser_10_reg),
                              .uc2rb_desc_3_axuser_11_reg(uc2rb_desc_3_axuser_11_reg),
                              .uc2rb_desc_3_axuser_12_reg(uc2rb_desc_3_axuser_12_reg),
                              .uc2rb_desc_3_axuser_13_reg(uc2rb_desc_3_axuser_13_reg),
                              .uc2rb_desc_3_axuser_14_reg(uc2rb_desc_3_axuser_14_reg),
                              .uc2rb_desc_3_axuser_15_reg(uc2rb_desc_3_axuser_15_reg),
                              .uc2rb_desc_3_wuser_0_reg(uc2rb_desc_3_wuser_0_reg),
                              .uc2rb_desc_3_wuser_1_reg(uc2rb_desc_3_wuser_1_reg),
                              .uc2rb_desc_3_wuser_2_reg(uc2rb_desc_3_wuser_2_reg),
                              .uc2rb_desc_3_wuser_3_reg(uc2rb_desc_3_wuser_3_reg),
                              .uc2rb_desc_3_wuser_4_reg(uc2rb_desc_3_wuser_4_reg),
                              .uc2rb_desc_3_wuser_5_reg(uc2rb_desc_3_wuser_5_reg),
                              .uc2rb_desc_3_wuser_6_reg(uc2rb_desc_3_wuser_6_reg),
                              .uc2rb_desc_3_wuser_7_reg(uc2rb_desc_3_wuser_7_reg),
                              .uc2rb_desc_3_wuser_8_reg(uc2rb_desc_3_wuser_8_reg),
                              .uc2rb_desc_3_wuser_9_reg(uc2rb_desc_3_wuser_9_reg),
                              .uc2rb_desc_3_wuser_10_reg(uc2rb_desc_3_wuser_10_reg),
                              .uc2rb_desc_3_wuser_11_reg(uc2rb_desc_3_wuser_11_reg),
                              .uc2rb_desc_3_wuser_12_reg(uc2rb_desc_3_wuser_12_reg),
                              .uc2rb_desc_3_wuser_13_reg(uc2rb_desc_3_wuser_13_reg),
                              .uc2rb_desc_3_wuser_14_reg(uc2rb_desc_3_wuser_14_reg),
                              .uc2rb_desc_3_wuser_15_reg(uc2rb_desc_3_wuser_15_reg),
                              .uc2rb_desc_4_txn_type_reg(uc2rb_desc_4_txn_type_reg),
                              .uc2rb_desc_4_size_reg(uc2rb_desc_4_size_reg),
                              .uc2rb_desc_4_data_offset_reg(uc2rb_desc_4_data_offset_reg),
                              .uc2rb_desc_4_axsize_reg(uc2rb_desc_4_axsize_reg),
                              .uc2rb_desc_4_attr_reg(uc2rb_desc_4_attr_reg),
                              .uc2rb_desc_4_axaddr_0_reg(uc2rb_desc_4_axaddr_0_reg),
                              .uc2rb_desc_4_axaddr_1_reg(uc2rb_desc_4_axaddr_1_reg),
                              .uc2rb_desc_4_axaddr_2_reg(uc2rb_desc_4_axaddr_2_reg),
                              .uc2rb_desc_4_axaddr_3_reg(uc2rb_desc_4_axaddr_3_reg),
                              .uc2rb_desc_4_axid_0_reg(uc2rb_desc_4_axid_0_reg),
                              .uc2rb_desc_4_axid_1_reg(uc2rb_desc_4_axid_1_reg),
                              .uc2rb_desc_4_axid_2_reg(uc2rb_desc_4_axid_2_reg),
                              .uc2rb_desc_4_axid_3_reg(uc2rb_desc_4_axid_3_reg),
                              .uc2rb_desc_4_axuser_0_reg(uc2rb_desc_4_axuser_0_reg),
                              .uc2rb_desc_4_axuser_1_reg(uc2rb_desc_4_axuser_1_reg),
                              .uc2rb_desc_4_axuser_2_reg(uc2rb_desc_4_axuser_2_reg),
                              .uc2rb_desc_4_axuser_3_reg(uc2rb_desc_4_axuser_3_reg),
                              .uc2rb_desc_4_axuser_4_reg(uc2rb_desc_4_axuser_4_reg),
                              .uc2rb_desc_4_axuser_5_reg(uc2rb_desc_4_axuser_5_reg),
                              .uc2rb_desc_4_axuser_6_reg(uc2rb_desc_4_axuser_6_reg),
                              .uc2rb_desc_4_axuser_7_reg(uc2rb_desc_4_axuser_7_reg),
                              .uc2rb_desc_4_axuser_8_reg(uc2rb_desc_4_axuser_8_reg),
                              .uc2rb_desc_4_axuser_9_reg(uc2rb_desc_4_axuser_9_reg),
                              .uc2rb_desc_4_axuser_10_reg(uc2rb_desc_4_axuser_10_reg),
                              .uc2rb_desc_4_axuser_11_reg(uc2rb_desc_4_axuser_11_reg),
                              .uc2rb_desc_4_axuser_12_reg(uc2rb_desc_4_axuser_12_reg),
                              .uc2rb_desc_4_axuser_13_reg(uc2rb_desc_4_axuser_13_reg),
                              .uc2rb_desc_4_axuser_14_reg(uc2rb_desc_4_axuser_14_reg),
                              .uc2rb_desc_4_axuser_15_reg(uc2rb_desc_4_axuser_15_reg),
                              .uc2rb_desc_4_wuser_0_reg(uc2rb_desc_4_wuser_0_reg),
                              .uc2rb_desc_4_wuser_1_reg(uc2rb_desc_4_wuser_1_reg),
                              .uc2rb_desc_4_wuser_2_reg(uc2rb_desc_4_wuser_2_reg),
                              .uc2rb_desc_4_wuser_3_reg(uc2rb_desc_4_wuser_3_reg),
                              .uc2rb_desc_4_wuser_4_reg(uc2rb_desc_4_wuser_4_reg),
                              .uc2rb_desc_4_wuser_5_reg(uc2rb_desc_4_wuser_5_reg),
                              .uc2rb_desc_4_wuser_6_reg(uc2rb_desc_4_wuser_6_reg),
                              .uc2rb_desc_4_wuser_7_reg(uc2rb_desc_4_wuser_7_reg),
                              .uc2rb_desc_4_wuser_8_reg(uc2rb_desc_4_wuser_8_reg),
                              .uc2rb_desc_4_wuser_9_reg(uc2rb_desc_4_wuser_9_reg),
                              .uc2rb_desc_4_wuser_10_reg(uc2rb_desc_4_wuser_10_reg),
                              .uc2rb_desc_4_wuser_11_reg(uc2rb_desc_4_wuser_11_reg),
                              .uc2rb_desc_4_wuser_12_reg(uc2rb_desc_4_wuser_12_reg),
                              .uc2rb_desc_4_wuser_13_reg(uc2rb_desc_4_wuser_13_reg),
                              .uc2rb_desc_4_wuser_14_reg(uc2rb_desc_4_wuser_14_reg),
                              .uc2rb_desc_4_wuser_15_reg(uc2rb_desc_4_wuser_15_reg),
                              .uc2rb_desc_5_txn_type_reg(uc2rb_desc_5_txn_type_reg),
                              .uc2rb_desc_5_size_reg(uc2rb_desc_5_size_reg),
                              .uc2rb_desc_5_data_offset_reg(uc2rb_desc_5_data_offset_reg),
                              .uc2rb_desc_5_axsize_reg(uc2rb_desc_5_axsize_reg),
                              .uc2rb_desc_5_attr_reg(uc2rb_desc_5_attr_reg),
                              .uc2rb_desc_5_axaddr_0_reg(uc2rb_desc_5_axaddr_0_reg),
                              .uc2rb_desc_5_axaddr_1_reg(uc2rb_desc_5_axaddr_1_reg),
                              .uc2rb_desc_5_axaddr_2_reg(uc2rb_desc_5_axaddr_2_reg),
                              .uc2rb_desc_5_axaddr_3_reg(uc2rb_desc_5_axaddr_3_reg),
                              .uc2rb_desc_5_axid_0_reg(uc2rb_desc_5_axid_0_reg),
                              .uc2rb_desc_5_axid_1_reg(uc2rb_desc_5_axid_1_reg),
                              .uc2rb_desc_5_axid_2_reg(uc2rb_desc_5_axid_2_reg),
                              .uc2rb_desc_5_axid_3_reg(uc2rb_desc_5_axid_3_reg),
                              .uc2rb_desc_5_axuser_0_reg(uc2rb_desc_5_axuser_0_reg),
                              .uc2rb_desc_5_axuser_1_reg(uc2rb_desc_5_axuser_1_reg),
                              .uc2rb_desc_5_axuser_2_reg(uc2rb_desc_5_axuser_2_reg),
                              .uc2rb_desc_5_axuser_3_reg(uc2rb_desc_5_axuser_3_reg),
                              .uc2rb_desc_5_axuser_4_reg(uc2rb_desc_5_axuser_4_reg),
                              .uc2rb_desc_5_axuser_5_reg(uc2rb_desc_5_axuser_5_reg),
                              .uc2rb_desc_5_axuser_6_reg(uc2rb_desc_5_axuser_6_reg),
                              .uc2rb_desc_5_axuser_7_reg(uc2rb_desc_5_axuser_7_reg),
                              .uc2rb_desc_5_axuser_8_reg(uc2rb_desc_5_axuser_8_reg),
                              .uc2rb_desc_5_axuser_9_reg(uc2rb_desc_5_axuser_9_reg),
                              .uc2rb_desc_5_axuser_10_reg(uc2rb_desc_5_axuser_10_reg),
                              .uc2rb_desc_5_axuser_11_reg(uc2rb_desc_5_axuser_11_reg),
                              .uc2rb_desc_5_axuser_12_reg(uc2rb_desc_5_axuser_12_reg),
                              .uc2rb_desc_5_axuser_13_reg(uc2rb_desc_5_axuser_13_reg),
                              .uc2rb_desc_5_axuser_14_reg(uc2rb_desc_5_axuser_14_reg),
                              .uc2rb_desc_5_axuser_15_reg(uc2rb_desc_5_axuser_15_reg),
                              .uc2rb_desc_5_wuser_0_reg(uc2rb_desc_5_wuser_0_reg),
                              .uc2rb_desc_5_wuser_1_reg(uc2rb_desc_5_wuser_1_reg),
                              .uc2rb_desc_5_wuser_2_reg(uc2rb_desc_5_wuser_2_reg),
                              .uc2rb_desc_5_wuser_3_reg(uc2rb_desc_5_wuser_3_reg),
                              .uc2rb_desc_5_wuser_4_reg(uc2rb_desc_5_wuser_4_reg),
                              .uc2rb_desc_5_wuser_5_reg(uc2rb_desc_5_wuser_5_reg),
                              .uc2rb_desc_5_wuser_6_reg(uc2rb_desc_5_wuser_6_reg),
                              .uc2rb_desc_5_wuser_7_reg(uc2rb_desc_5_wuser_7_reg),
                              .uc2rb_desc_5_wuser_8_reg(uc2rb_desc_5_wuser_8_reg),
                              .uc2rb_desc_5_wuser_9_reg(uc2rb_desc_5_wuser_9_reg),
                              .uc2rb_desc_5_wuser_10_reg(uc2rb_desc_5_wuser_10_reg),
                              .uc2rb_desc_5_wuser_11_reg(uc2rb_desc_5_wuser_11_reg),
                              .uc2rb_desc_5_wuser_12_reg(uc2rb_desc_5_wuser_12_reg),
                              .uc2rb_desc_5_wuser_13_reg(uc2rb_desc_5_wuser_13_reg),
                              .uc2rb_desc_5_wuser_14_reg(uc2rb_desc_5_wuser_14_reg),
                              .uc2rb_desc_5_wuser_15_reg(uc2rb_desc_5_wuser_15_reg),
                              .uc2rb_desc_6_txn_type_reg(uc2rb_desc_6_txn_type_reg),
                              .uc2rb_desc_6_size_reg(uc2rb_desc_6_size_reg),
                              .uc2rb_desc_6_data_offset_reg(uc2rb_desc_6_data_offset_reg),
                              .uc2rb_desc_6_axsize_reg(uc2rb_desc_6_axsize_reg),
                              .uc2rb_desc_6_attr_reg(uc2rb_desc_6_attr_reg),
                              .uc2rb_desc_6_axaddr_0_reg(uc2rb_desc_6_axaddr_0_reg),
                              .uc2rb_desc_6_axaddr_1_reg(uc2rb_desc_6_axaddr_1_reg),
                              .uc2rb_desc_6_axaddr_2_reg(uc2rb_desc_6_axaddr_2_reg),
                              .uc2rb_desc_6_axaddr_3_reg(uc2rb_desc_6_axaddr_3_reg),
                              .uc2rb_desc_6_axid_0_reg(uc2rb_desc_6_axid_0_reg),
                              .uc2rb_desc_6_axid_1_reg(uc2rb_desc_6_axid_1_reg),
                              .uc2rb_desc_6_axid_2_reg(uc2rb_desc_6_axid_2_reg),
                              .uc2rb_desc_6_axid_3_reg(uc2rb_desc_6_axid_3_reg),
                              .uc2rb_desc_6_axuser_0_reg(uc2rb_desc_6_axuser_0_reg),
                              .uc2rb_desc_6_axuser_1_reg(uc2rb_desc_6_axuser_1_reg),
                              .uc2rb_desc_6_axuser_2_reg(uc2rb_desc_6_axuser_2_reg),
                              .uc2rb_desc_6_axuser_3_reg(uc2rb_desc_6_axuser_3_reg),
                              .uc2rb_desc_6_axuser_4_reg(uc2rb_desc_6_axuser_4_reg),
                              .uc2rb_desc_6_axuser_5_reg(uc2rb_desc_6_axuser_5_reg),
                              .uc2rb_desc_6_axuser_6_reg(uc2rb_desc_6_axuser_6_reg),
                              .uc2rb_desc_6_axuser_7_reg(uc2rb_desc_6_axuser_7_reg),
                              .uc2rb_desc_6_axuser_8_reg(uc2rb_desc_6_axuser_8_reg),
                              .uc2rb_desc_6_axuser_9_reg(uc2rb_desc_6_axuser_9_reg),
                              .uc2rb_desc_6_axuser_10_reg(uc2rb_desc_6_axuser_10_reg),
                              .uc2rb_desc_6_axuser_11_reg(uc2rb_desc_6_axuser_11_reg),
                              .uc2rb_desc_6_axuser_12_reg(uc2rb_desc_6_axuser_12_reg),
                              .uc2rb_desc_6_axuser_13_reg(uc2rb_desc_6_axuser_13_reg),
                              .uc2rb_desc_6_axuser_14_reg(uc2rb_desc_6_axuser_14_reg),
                              .uc2rb_desc_6_axuser_15_reg(uc2rb_desc_6_axuser_15_reg),
                              .uc2rb_desc_6_wuser_0_reg(uc2rb_desc_6_wuser_0_reg),
                              .uc2rb_desc_6_wuser_1_reg(uc2rb_desc_6_wuser_1_reg),
                              .uc2rb_desc_6_wuser_2_reg(uc2rb_desc_6_wuser_2_reg),
                              .uc2rb_desc_6_wuser_3_reg(uc2rb_desc_6_wuser_3_reg),
                              .uc2rb_desc_6_wuser_4_reg(uc2rb_desc_6_wuser_4_reg),
                              .uc2rb_desc_6_wuser_5_reg(uc2rb_desc_6_wuser_5_reg),
                              .uc2rb_desc_6_wuser_6_reg(uc2rb_desc_6_wuser_6_reg),
                              .uc2rb_desc_6_wuser_7_reg(uc2rb_desc_6_wuser_7_reg),
                              .uc2rb_desc_6_wuser_8_reg(uc2rb_desc_6_wuser_8_reg),
                              .uc2rb_desc_6_wuser_9_reg(uc2rb_desc_6_wuser_9_reg),
                              .uc2rb_desc_6_wuser_10_reg(uc2rb_desc_6_wuser_10_reg),
                              .uc2rb_desc_6_wuser_11_reg(uc2rb_desc_6_wuser_11_reg),
                              .uc2rb_desc_6_wuser_12_reg(uc2rb_desc_6_wuser_12_reg),
                              .uc2rb_desc_6_wuser_13_reg(uc2rb_desc_6_wuser_13_reg),
                              .uc2rb_desc_6_wuser_14_reg(uc2rb_desc_6_wuser_14_reg),
                              .uc2rb_desc_6_wuser_15_reg(uc2rb_desc_6_wuser_15_reg),
                              .uc2rb_desc_7_txn_type_reg(uc2rb_desc_7_txn_type_reg),
                              .uc2rb_desc_7_size_reg(uc2rb_desc_7_size_reg),
                              .uc2rb_desc_7_data_offset_reg(uc2rb_desc_7_data_offset_reg),
                              .uc2rb_desc_7_axsize_reg(uc2rb_desc_7_axsize_reg),
                              .uc2rb_desc_7_attr_reg(uc2rb_desc_7_attr_reg),
                              .uc2rb_desc_7_axaddr_0_reg(uc2rb_desc_7_axaddr_0_reg),
                              .uc2rb_desc_7_axaddr_1_reg(uc2rb_desc_7_axaddr_1_reg),
                              .uc2rb_desc_7_axaddr_2_reg(uc2rb_desc_7_axaddr_2_reg),
                              .uc2rb_desc_7_axaddr_3_reg(uc2rb_desc_7_axaddr_3_reg),
                              .uc2rb_desc_7_axid_0_reg(uc2rb_desc_7_axid_0_reg),
                              .uc2rb_desc_7_axid_1_reg(uc2rb_desc_7_axid_1_reg),
                              .uc2rb_desc_7_axid_2_reg(uc2rb_desc_7_axid_2_reg),
                              .uc2rb_desc_7_axid_3_reg(uc2rb_desc_7_axid_3_reg),
                              .uc2rb_desc_7_axuser_0_reg(uc2rb_desc_7_axuser_0_reg),
                              .uc2rb_desc_7_axuser_1_reg(uc2rb_desc_7_axuser_1_reg),
                              .uc2rb_desc_7_axuser_2_reg(uc2rb_desc_7_axuser_2_reg),
                              .uc2rb_desc_7_axuser_3_reg(uc2rb_desc_7_axuser_3_reg),
                              .uc2rb_desc_7_axuser_4_reg(uc2rb_desc_7_axuser_4_reg),
                              .uc2rb_desc_7_axuser_5_reg(uc2rb_desc_7_axuser_5_reg),
                              .uc2rb_desc_7_axuser_6_reg(uc2rb_desc_7_axuser_6_reg),
                              .uc2rb_desc_7_axuser_7_reg(uc2rb_desc_7_axuser_7_reg),
                              .uc2rb_desc_7_axuser_8_reg(uc2rb_desc_7_axuser_8_reg),
                              .uc2rb_desc_7_axuser_9_reg(uc2rb_desc_7_axuser_9_reg),
                              .uc2rb_desc_7_axuser_10_reg(uc2rb_desc_7_axuser_10_reg),
                              .uc2rb_desc_7_axuser_11_reg(uc2rb_desc_7_axuser_11_reg),
                              .uc2rb_desc_7_axuser_12_reg(uc2rb_desc_7_axuser_12_reg),
                              .uc2rb_desc_7_axuser_13_reg(uc2rb_desc_7_axuser_13_reg),
                              .uc2rb_desc_7_axuser_14_reg(uc2rb_desc_7_axuser_14_reg),
                              .uc2rb_desc_7_axuser_15_reg(uc2rb_desc_7_axuser_15_reg),
                              .uc2rb_desc_7_wuser_0_reg(uc2rb_desc_7_wuser_0_reg),
                              .uc2rb_desc_7_wuser_1_reg(uc2rb_desc_7_wuser_1_reg),
                              .uc2rb_desc_7_wuser_2_reg(uc2rb_desc_7_wuser_2_reg),
                              .uc2rb_desc_7_wuser_3_reg(uc2rb_desc_7_wuser_3_reg),
                              .uc2rb_desc_7_wuser_4_reg(uc2rb_desc_7_wuser_4_reg),
                              .uc2rb_desc_7_wuser_5_reg(uc2rb_desc_7_wuser_5_reg),
                              .uc2rb_desc_7_wuser_6_reg(uc2rb_desc_7_wuser_6_reg),
                              .uc2rb_desc_7_wuser_7_reg(uc2rb_desc_7_wuser_7_reg),
                              .uc2rb_desc_7_wuser_8_reg(uc2rb_desc_7_wuser_8_reg),
                              .uc2rb_desc_7_wuser_9_reg(uc2rb_desc_7_wuser_9_reg),
                              .uc2rb_desc_7_wuser_10_reg(uc2rb_desc_7_wuser_10_reg),
                              .uc2rb_desc_7_wuser_11_reg(uc2rb_desc_7_wuser_11_reg),
                              .uc2rb_desc_7_wuser_12_reg(uc2rb_desc_7_wuser_12_reg),
                              .uc2rb_desc_7_wuser_13_reg(uc2rb_desc_7_wuser_13_reg),
                              .uc2rb_desc_7_wuser_14_reg(uc2rb_desc_7_wuser_14_reg),
                              .uc2rb_desc_7_wuser_15_reg(uc2rb_desc_7_wuser_15_reg),
                              .uc2rb_desc_8_txn_type_reg(uc2rb_desc_8_txn_type_reg),
                              .uc2rb_desc_8_size_reg(uc2rb_desc_8_size_reg),
                              .uc2rb_desc_8_data_offset_reg(uc2rb_desc_8_data_offset_reg),
                              .uc2rb_desc_8_axsize_reg(uc2rb_desc_8_axsize_reg),
                              .uc2rb_desc_8_attr_reg(uc2rb_desc_8_attr_reg),
                              .uc2rb_desc_8_axaddr_0_reg(uc2rb_desc_8_axaddr_0_reg),
                              .uc2rb_desc_8_axaddr_1_reg(uc2rb_desc_8_axaddr_1_reg),
                              .uc2rb_desc_8_axaddr_2_reg(uc2rb_desc_8_axaddr_2_reg),
                              .uc2rb_desc_8_axaddr_3_reg(uc2rb_desc_8_axaddr_3_reg),
                              .uc2rb_desc_8_axid_0_reg(uc2rb_desc_8_axid_0_reg),
                              .uc2rb_desc_8_axid_1_reg(uc2rb_desc_8_axid_1_reg),
                              .uc2rb_desc_8_axid_2_reg(uc2rb_desc_8_axid_2_reg),
                              .uc2rb_desc_8_axid_3_reg(uc2rb_desc_8_axid_3_reg),
                              .uc2rb_desc_8_axuser_0_reg(uc2rb_desc_8_axuser_0_reg),
                              .uc2rb_desc_8_axuser_1_reg(uc2rb_desc_8_axuser_1_reg),
                              .uc2rb_desc_8_axuser_2_reg(uc2rb_desc_8_axuser_2_reg),
                              .uc2rb_desc_8_axuser_3_reg(uc2rb_desc_8_axuser_3_reg),
                              .uc2rb_desc_8_axuser_4_reg(uc2rb_desc_8_axuser_4_reg),
                              .uc2rb_desc_8_axuser_5_reg(uc2rb_desc_8_axuser_5_reg),
                              .uc2rb_desc_8_axuser_6_reg(uc2rb_desc_8_axuser_6_reg),
                              .uc2rb_desc_8_axuser_7_reg(uc2rb_desc_8_axuser_7_reg),
                              .uc2rb_desc_8_axuser_8_reg(uc2rb_desc_8_axuser_8_reg),
                              .uc2rb_desc_8_axuser_9_reg(uc2rb_desc_8_axuser_9_reg),
                              .uc2rb_desc_8_axuser_10_reg(uc2rb_desc_8_axuser_10_reg),
                              .uc2rb_desc_8_axuser_11_reg(uc2rb_desc_8_axuser_11_reg),
                              .uc2rb_desc_8_axuser_12_reg(uc2rb_desc_8_axuser_12_reg),
                              .uc2rb_desc_8_axuser_13_reg(uc2rb_desc_8_axuser_13_reg),
                              .uc2rb_desc_8_axuser_14_reg(uc2rb_desc_8_axuser_14_reg),
                              .uc2rb_desc_8_axuser_15_reg(uc2rb_desc_8_axuser_15_reg),
                              .uc2rb_desc_8_wuser_0_reg(uc2rb_desc_8_wuser_0_reg),
                              .uc2rb_desc_8_wuser_1_reg(uc2rb_desc_8_wuser_1_reg),
                              .uc2rb_desc_8_wuser_2_reg(uc2rb_desc_8_wuser_2_reg),
                              .uc2rb_desc_8_wuser_3_reg(uc2rb_desc_8_wuser_3_reg),
                              .uc2rb_desc_8_wuser_4_reg(uc2rb_desc_8_wuser_4_reg),
                              .uc2rb_desc_8_wuser_5_reg(uc2rb_desc_8_wuser_5_reg),
                              .uc2rb_desc_8_wuser_6_reg(uc2rb_desc_8_wuser_6_reg),
                              .uc2rb_desc_8_wuser_7_reg(uc2rb_desc_8_wuser_7_reg),
                              .uc2rb_desc_8_wuser_8_reg(uc2rb_desc_8_wuser_8_reg),
                              .uc2rb_desc_8_wuser_9_reg(uc2rb_desc_8_wuser_9_reg),
                              .uc2rb_desc_8_wuser_10_reg(uc2rb_desc_8_wuser_10_reg),
                              .uc2rb_desc_8_wuser_11_reg(uc2rb_desc_8_wuser_11_reg),
                              .uc2rb_desc_8_wuser_12_reg(uc2rb_desc_8_wuser_12_reg),
                              .uc2rb_desc_8_wuser_13_reg(uc2rb_desc_8_wuser_13_reg),
                              .uc2rb_desc_8_wuser_14_reg(uc2rb_desc_8_wuser_14_reg),
                              .uc2rb_desc_8_wuser_15_reg(uc2rb_desc_8_wuser_15_reg),
                              .uc2rb_desc_9_txn_type_reg(uc2rb_desc_9_txn_type_reg),
                              .uc2rb_desc_9_size_reg(uc2rb_desc_9_size_reg),
                              .uc2rb_desc_9_data_offset_reg(uc2rb_desc_9_data_offset_reg),
                              .uc2rb_desc_9_axsize_reg(uc2rb_desc_9_axsize_reg),
                              .uc2rb_desc_9_attr_reg(uc2rb_desc_9_attr_reg),
                              .uc2rb_desc_9_axaddr_0_reg(uc2rb_desc_9_axaddr_0_reg),
                              .uc2rb_desc_9_axaddr_1_reg(uc2rb_desc_9_axaddr_1_reg),
                              .uc2rb_desc_9_axaddr_2_reg(uc2rb_desc_9_axaddr_2_reg),
                              .uc2rb_desc_9_axaddr_3_reg(uc2rb_desc_9_axaddr_3_reg),
                              .uc2rb_desc_9_axid_0_reg(uc2rb_desc_9_axid_0_reg),
                              .uc2rb_desc_9_axid_1_reg(uc2rb_desc_9_axid_1_reg),
                              .uc2rb_desc_9_axid_2_reg(uc2rb_desc_9_axid_2_reg),
                              .uc2rb_desc_9_axid_3_reg(uc2rb_desc_9_axid_3_reg),
                              .uc2rb_desc_9_axuser_0_reg(uc2rb_desc_9_axuser_0_reg),
                              .uc2rb_desc_9_axuser_1_reg(uc2rb_desc_9_axuser_1_reg),
                              .uc2rb_desc_9_axuser_2_reg(uc2rb_desc_9_axuser_2_reg),
                              .uc2rb_desc_9_axuser_3_reg(uc2rb_desc_9_axuser_3_reg),
                              .uc2rb_desc_9_axuser_4_reg(uc2rb_desc_9_axuser_4_reg),
                              .uc2rb_desc_9_axuser_5_reg(uc2rb_desc_9_axuser_5_reg),
                              .uc2rb_desc_9_axuser_6_reg(uc2rb_desc_9_axuser_6_reg),
                              .uc2rb_desc_9_axuser_7_reg(uc2rb_desc_9_axuser_7_reg),
                              .uc2rb_desc_9_axuser_8_reg(uc2rb_desc_9_axuser_8_reg),
                              .uc2rb_desc_9_axuser_9_reg(uc2rb_desc_9_axuser_9_reg),
                              .uc2rb_desc_9_axuser_10_reg(uc2rb_desc_9_axuser_10_reg),
                              .uc2rb_desc_9_axuser_11_reg(uc2rb_desc_9_axuser_11_reg),
                              .uc2rb_desc_9_axuser_12_reg(uc2rb_desc_9_axuser_12_reg),
                              .uc2rb_desc_9_axuser_13_reg(uc2rb_desc_9_axuser_13_reg),
                              .uc2rb_desc_9_axuser_14_reg(uc2rb_desc_9_axuser_14_reg),
                              .uc2rb_desc_9_axuser_15_reg(uc2rb_desc_9_axuser_15_reg),
                              .uc2rb_desc_9_wuser_0_reg(uc2rb_desc_9_wuser_0_reg),
                              .uc2rb_desc_9_wuser_1_reg(uc2rb_desc_9_wuser_1_reg),
                              .uc2rb_desc_9_wuser_2_reg(uc2rb_desc_9_wuser_2_reg),
                              .uc2rb_desc_9_wuser_3_reg(uc2rb_desc_9_wuser_3_reg),
                              .uc2rb_desc_9_wuser_4_reg(uc2rb_desc_9_wuser_4_reg),
                              .uc2rb_desc_9_wuser_5_reg(uc2rb_desc_9_wuser_5_reg),
                              .uc2rb_desc_9_wuser_6_reg(uc2rb_desc_9_wuser_6_reg),
                              .uc2rb_desc_9_wuser_7_reg(uc2rb_desc_9_wuser_7_reg),
                              .uc2rb_desc_9_wuser_8_reg(uc2rb_desc_9_wuser_8_reg),
                              .uc2rb_desc_9_wuser_9_reg(uc2rb_desc_9_wuser_9_reg),
                              .uc2rb_desc_9_wuser_10_reg(uc2rb_desc_9_wuser_10_reg),
                              .uc2rb_desc_9_wuser_11_reg(uc2rb_desc_9_wuser_11_reg),
                              .uc2rb_desc_9_wuser_12_reg(uc2rb_desc_9_wuser_12_reg),
                              .uc2rb_desc_9_wuser_13_reg(uc2rb_desc_9_wuser_13_reg),
                              .uc2rb_desc_9_wuser_14_reg(uc2rb_desc_9_wuser_14_reg),
                              .uc2rb_desc_9_wuser_15_reg(uc2rb_desc_9_wuser_15_reg),
                              .uc2rb_desc_10_txn_type_reg(uc2rb_desc_10_txn_type_reg),
                              .uc2rb_desc_10_size_reg(uc2rb_desc_10_size_reg),
                              .uc2rb_desc_10_data_offset_reg(uc2rb_desc_10_data_offset_reg),
                              .uc2rb_desc_10_axsize_reg(uc2rb_desc_10_axsize_reg),
                              .uc2rb_desc_10_attr_reg(uc2rb_desc_10_attr_reg),
                              .uc2rb_desc_10_axaddr_0_reg(uc2rb_desc_10_axaddr_0_reg),
                              .uc2rb_desc_10_axaddr_1_reg(uc2rb_desc_10_axaddr_1_reg),
                              .uc2rb_desc_10_axaddr_2_reg(uc2rb_desc_10_axaddr_2_reg),
                              .uc2rb_desc_10_axaddr_3_reg(uc2rb_desc_10_axaddr_3_reg),
                              .uc2rb_desc_10_axid_0_reg(uc2rb_desc_10_axid_0_reg),
                              .uc2rb_desc_10_axid_1_reg(uc2rb_desc_10_axid_1_reg),
                              .uc2rb_desc_10_axid_2_reg(uc2rb_desc_10_axid_2_reg),
                              .uc2rb_desc_10_axid_3_reg(uc2rb_desc_10_axid_3_reg),
                              .uc2rb_desc_10_axuser_0_reg(uc2rb_desc_10_axuser_0_reg),
                              .uc2rb_desc_10_axuser_1_reg(uc2rb_desc_10_axuser_1_reg),
                              .uc2rb_desc_10_axuser_2_reg(uc2rb_desc_10_axuser_2_reg),
                              .uc2rb_desc_10_axuser_3_reg(uc2rb_desc_10_axuser_3_reg),
                              .uc2rb_desc_10_axuser_4_reg(uc2rb_desc_10_axuser_4_reg),
                              .uc2rb_desc_10_axuser_5_reg(uc2rb_desc_10_axuser_5_reg),
                              .uc2rb_desc_10_axuser_6_reg(uc2rb_desc_10_axuser_6_reg),
                              .uc2rb_desc_10_axuser_7_reg(uc2rb_desc_10_axuser_7_reg),
                              .uc2rb_desc_10_axuser_8_reg(uc2rb_desc_10_axuser_8_reg),
                              .uc2rb_desc_10_axuser_9_reg(uc2rb_desc_10_axuser_9_reg),
                              .uc2rb_desc_10_axuser_10_reg(uc2rb_desc_10_axuser_10_reg),
                              .uc2rb_desc_10_axuser_11_reg(uc2rb_desc_10_axuser_11_reg),
                              .uc2rb_desc_10_axuser_12_reg(uc2rb_desc_10_axuser_12_reg),
                              .uc2rb_desc_10_axuser_13_reg(uc2rb_desc_10_axuser_13_reg),
                              .uc2rb_desc_10_axuser_14_reg(uc2rb_desc_10_axuser_14_reg),
                              .uc2rb_desc_10_axuser_15_reg(uc2rb_desc_10_axuser_15_reg),
                              .uc2rb_desc_10_wuser_0_reg(uc2rb_desc_10_wuser_0_reg),
                              .uc2rb_desc_10_wuser_1_reg(uc2rb_desc_10_wuser_1_reg),
                              .uc2rb_desc_10_wuser_2_reg(uc2rb_desc_10_wuser_2_reg),
                              .uc2rb_desc_10_wuser_3_reg(uc2rb_desc_10_wuser_3_reg),
                              .uc2rb_desc_10_wuser_4_reg(uc2rb_desc_10_wuser_4_reg),
                              .uc2rb_desc_10_wuser_5_reg(uc2rb_desc_10_wuser_5_reg),
                              .uc2rb_desc_10_wuser_6_reg(uc2rb_desc_10_wuser_6_reg),
                              .uc2rb_desc_10_wuser_7_reg(uc2rb_desc_10_wuser_7_reg),
                              .uc2rb_desc_10_wuser_8_reg(uc2rb_desc_10_wuser_8_reg),
                              .uc2rb_desc_10_wuser_9_reg(uc2rb_desc_10_wuser_9_reg),
                              .uc2rb_desc_10_wuser_10_reg(uc2rb_desc_10_wuser_10_reg),
                              .uc2rb_desc_10_wuser_11_reg(uc2rb_desc_10_wuser_11_reg),
                              .uc2rb_desc_10_wuser_12_reg(uc2rb_desc_10_wuser_12_reg),
                              .uc2rb_desc_10_wuser_13_reg(uc2rb_desc_10_wuser_13_reg),
                              .uc2rb_desc_10_wuser_14_reg(uc2rb_desc_10_wuser_14_reg),
                              .uc2rb_desc_10_wuser_15_reg(uc2rb_desc_10_wuser_15_reg),
                              .uc2rb_desc_11_txn_type_reg(uc2rb_desc_11_txn_type_reg),
                              .uc2rb_desc_11_size_reg(uc2rb_desc_11_size_reg),
                              .uc2rb_desc_11_data_offset_reg(uc2rb_desc_11_data_offset_reg),
                              .uc2rb_desc_11_axsize_reg(uc2rb_desc_11_axsize_reg),
                              .uc2rb_desc_11_attr_reg(uc2rb_desc_11_attr_reg),
                              .uc2rb_desc_11_axaddr_0_reg(uc2rb_desc_11_axaddr_0_reg),
                              .uc2rb_desc_11_axaddr_1_reg(uc2rb_desc_11_axaddr_1_reg),
                              .uc2rb_desc_11_axaddr_2_reg(uc2rb_desc_11_axaddr_2_reg),
                              .uc2rb_desc_11_axaddr_3_reg(uc2rb_desc_11_axaddr_3_reg),
                              .uc2rb_desc_11_axid_0_reg(uc2rb_desc_11_axid_0_reg),
                              .uc2rb_desc_11_axid_1_reg(uc2rb_desc_11_axid_1_reg),
                              .uc2rb_desc_11_axid_2_reg(uc2rb_desc_11_axid_2_reg),
                              .uc2rb_desc_11_axid_3_reg(uc2rb_desc_11_axid_3_reg),
                              .uc2rb_desc_11_axuser_0_reg(uc2rb_desc_11_axuser_0_reg),
                              .uc2rb_desc_11_axuser_1_reg(uc2rb_desc_11_axuser_1_reg),
                              .uc2rb_desc_11_axuser_2_reg(uc2rb_desc_11_axuser_2_reg),
                              .uc2rb_desc_11_axuser_3_reg(uc2rb_desc_11_axuser_3_reg),
                              .uc2rb_desc_11_axuser_4_reg(uc2rb_desc_11_axuser_4_reg),
                              .uc2rb_desc_11_axuser_5_reg(uc2rb_desc_11_axuser_5_reg),
                              .uc2rb_desc_11_axuser_6_reg(uc2rb_desc_11_axuser_6_reg),
                              .uc2rb_desc_11_axuser_7_reg(uc2rb_desc_11_axuser_7_reg),
                              .uc2rb_desc_11_axuser_8_reg(uc2rb_desc_11_axuser_8_reg),
                              .uc2rb_desc_11_axuser_9_reg(uc2rb_desc_11_axuser_9_reg),
                              .uc2rb_desc_11_axuser_10_reg(uc2rb_desc_11_axuser_10_reg),
                              .uc2rb_desc_11_axuser_11_reg(uc2rb_desc_11_axuser_11_reg),
                              .uc2rb_desc_11_axuser_12_reg(uc2rb_desc_11_axuser_12_reg),
                              .uc2rb_desc_11_axuser_13_reg(uc2rb_desc_11_axuser_13_reg),
                              .uc2rb_desc_11_axuser_14_reg(uc2rb_desc_11_axuser_14_reg),
                              .uc2rb_desc_11_axuser_15_reg(uc2rb_desc_11_axuser_15_reg),
                              .uc2rb_desc_11_wuser_0_reg(uc2rb_desc_11_wuser_0_reg),
                              .uc2rb_desc_11_wuser_1_reg(uc2rb_desc_11_wuser_1_reg),
                              .uc2rb_desc_11_wuser_2_reg(uc2rb_desc_11_wuser_2_reg),
                              .uc2rb_desc_11_wuser_3_reg(uc2rb_desc_11_wuser_3_reg),
                              .uc2rb_desc_11_wuser_4_reg(uc2rb_desc_11_wuser_4_reg),
                              .uc2rb_desc_11_wuser_5_reg(uc2rb_desc_11_wuser_5_reg),
                              .uc2rb_desc_11_wuser_6_reg(uc2rb_desc_11_wuser_6_reg),
                              .uc2rb_desc_11_wuser_7_reg(uc2rb_desc_11_wuser_7_reg),
                              .uc2rb_desc_11_wuser_8_reg(uc2rb_desc_11_wuser_8_reg),
                              .uc2rb_desc_11_wuser_9_reg(uc2rb_desc_11_wuser_9_reg),
                              .uc2rb_desc_11_wuser_10_reg(uc2rb_desc_11_wuser_10_reg),
                              .uc2rb_desc_11_wuser_11_reg(uc2rb_desc_11_wuser_11_reg),
                              .uc2rb_desc_11_wuser_12_reg(uc2rb_desc_11_wuser_12_reg),
                              .uc2rb_desc_11_wuser_13_reg(uc2rb_desc_11_wuser_13_reg),
                              .uc2rb_desc_11_wuser_14_reg(uc2rb_desc_11_wuser_14_reg),
                              .uc2rb_desc_11_wuser_15_reg(uc2rb_desc_11_wuser_15_reg),
                              .uc2rb_desc_12_txn_type_reg(uc2rb_desc_12_txn_type_reg),
                              .uc2rb_desc_12_size_reg(uc2rb_desc_12_size_reg),
                              .uc2rb_desc_12_data_offset_reg(uc2rb_desc_12_data_offset_reg),
                              .uc2rb_desc_12_axsize_reg(uc2rb_desc_12_axsize_reg),
                              .uc2rb_desc_12_attr_reg(uc2rb_desc_12_attr_reg),
                              .uc2rb_desc_12_axaddr_0_reg(uc2rb_desc_12_axaddr_0_reg),
                              .uc2rb_desc_12_axaddr_1_reg(uc2rb_desc_12_axaddr_1_reg),
                              .uc2rb_desc_12_axaddr_2_reg(uc2rb_desc_12_axaddr_2_reg),
                              .uc2rb_desc_12_axaddr_3_reg(uc2rb_desc_12_axaddr_3_reg),
                              .uc2rb_desc_12_axid_0_reg(uc2rb_desc_12_axid_0_reg),
                              .uc2rb_desc_12_axid_1_reg(uc2rb_desc_12_axid_1_reg),
                              .uc2rb_desc_12_axid_2_reg(uc2rb_desc_12_axid_2_reg),
                              .uc2rb_desc_12_axid_3_reg(uc2rb_desc_12_axid_3_reg),
                              .uc2rb_desc_12_axuser_0_reg(uc2rb_desc_12_axuser_0_reg),
                              .uc2rb_desc_12_axuser_1_reg(uc2rb_desc_12_axuser_1_reg),
                              .uc2rb_desc_12_axuser_2_reg(uc2rb_desc_12_axuser_2_reg),
                              .uc2rb_desc_12_axuser_3_reg(uc2rb_desc_12_axuser_3_reg),
                              .uc2rb_desc_12_axuser_4_reg(uc2rb_desc_12_axuser_4_reg),
                              .uc2rb_desc_12_axuser_5_reg(uc2rb_desc_12_axuser_5_reg),
                              .uc2rb_desc_12_axuser_6_reg(uc2rb_desc_12_axuser_6_reg),
                              .uc2rb_desc_12_axuser_7_reg(uc2rb_desc_12_axuser_7_reg),
                              .uc2rb_desc_12_axuser_8_reg(uc2rb_desc_12_axuser_8_reg),
                              .uc2rb_desc_12_axuser_9_reg(uc2rb_desc_12_axuser_9_reg),
                              .uc2rb_desc_12_axuser_10_reg(uc2rb_desc_12_axuser_10_reg),
                              .uc2rb_desc_12_axuser_11_reg(uc2rb_desc_12_axuser_11_reg),
                              .uc2rb_desc_12_axuser_12_reg(uc2rb_desc_12_axuser_12_reg),
                              .uc2rb_desc_12_axuser_13_reg(uc2rb_desc_12_axuser_13_reg),
                              .uc2rb_desc_12_axuser_14_reg(uc2rb_desc_12_axuser_14_reg),
                              .uc2rb_desc_12_axuser_15_reg(uc2rb_desc_12_axuser_15_reg),
                              .uc2rb_desc_12_wuser_0_reg(uc2rb_desc_12_wuser_0_reg),
                              .uc2rb_desc_12_wuser_1_reg(uc2rb_desc_12_wuser_1_reg),
                              .uc2rb_desc_12_wuser_2_reg(uc2rb_desc_12_wuser_2_reg),
                              .uc2rb_desc_12_wuser_3_reg(uc2rb_desc_12_wuser_3_reg),
                              .uc2rb_desc_12_wuser_4_reg(uc2rb_desc_12_wuser_4_reg),
                              .uc2rb_desc_12_wuser_5_reg(uc2rb_desc_12_wuser_5_reg),
                              .uc2rb_desc_12_wuser_6_reg(uc2rb_desc_12_wuser_6_reg),
                              .uc2rb_desc_12_wuser_7_reg(uc2rb_desc_12_wuser_7_reg),
                              .uc2rb_desc_12_wuser_8_reg(uc2rb_desc_12_wuser_8_reg),
                              .uc2rb_desc_12_wuser_9_reg(uc2rb_desc_12_wuser_9_reg),
                              .uc2rb_desc_12_wuser_10_reg(uc2rb_desc_12_wuser_10_reg),
                              .uc2rb_desc_12_wuser_11_reg(uc2rb_desc_12_wuser_11_reg),
                              .uc2rb_desc_12_wuser_12_reg(uc2rb_desc_12_wuser_12_reg),
                              .uc2rb_desc_12_wuser_13_reg(uc2rb_desc_12_wuser_13_reg),
                              .uc2rb_desc_12_wuser_14_reg(uc2rb_desc_12_wuser_14_reg),
                              .uc2rb_desc_12_wuser_15_reg(uc2rb_desc_12_wuser_15_reg),
                              .uc2rb_desc_13_txn_type_reg(uc2rb_desc_13_txn_type_reg),
                              .uc2rb_desc_13_size_reg(uc2rb_desc_13_size_reg),
                              .uc2rb_desc_13_data_offset_reg(uc2rb_desc_13_data_offset_reg),
                              .uc2rb_desc_13_axsize_reg(uc2rb_desc_13_axsize_reg),
                              .uc2rb_desc_13_attr_reg(uc2rb_desc_13_attr_reg),
                              .uc2rb_desc_13_axaddr_0_reg(uc2rb_desc_13_axaddr_0_reg),
                              .uc2rb_desc_13_axaddr_1_reg(uc2rb_desc_13_axaddr_1_reg),
                              .uc2rb_desc_13_axaddr_2_reg(uc2rb_desc_13_axaddr_2_reg),
                              .uc2rb_desc_13_axaddr_3_reg(uc2rb_desc_13_axaddr_3_reg),
                              .uc2rb_desc_13_axid_0_reg(uc2rb_desc_13_axid_0_reg),
                              .uc2rb_desc_13_axid_1_reg(uc2rb_desc_13_axid_1_reg),
                              .uc2rb_desc_13_axid_2_reg(uc2rb_desc_13_axid_2_reg),
                              .uc2rb_desc_13_axid_3_reg(uc2rb_desc_13_axid_3_reg),
                              .uc2rb_desc_13_axuser_0_reg(uc2rb_desc_13_axuser_0_reg),
                              .uc2rb_desc_13_axuser_1_reg(uc2rb_desc_13_axuser_1_reg),
                              .uc2rb_desc_13_axuser_2_reg(uc2rb_desc_13_axuser_2_reg),
                              .uc2rb_desc_13_axuser_3_reg(uc2rb_desc_13_axuser_3_reg),
                              .uc2rb_desc_13_axuser_4_reg(uc2rb_desc_13_axuser_4_reg),
                              .uc2rb_desc_13_axuser_5_reg(uc2rb_desc_13_axuser_5_reg),
                              .uc2rb_desc_13_axuser_6_reg(uc2rb_desc_13_axuser_6_reg),
                              .uc2rb_desc_13_axuser_7_reg(uc2rb_desc_13_axuser_7_reg),
                              .uc2rb_desc_13_axuser_8_reg(uc2rb_desc_13_axuser_8_reg),
                              .uc2rb_desc_13_axuser_9_reg(uc2rb_desc_13_axuser_9_reg),
                              .uc2rb_desc_13_axuser_10_reg(uc2rb_desc_13_axuser_10_reg),
                              .uc2rb_desc_13_axuser_11_reg(uc2rb_desc_13_axuser_11_reg),
                              .uc2rb_desc_13_axuser_12_reg(uc2rb_desc_13_axuser_12_reg),
                              .uc2rb_desc_13_axuser_13_reg(uc2rb_desc_13_axuser_13_reg),
                              .uc2rb_desc_13_axuser_14_reg(uc2rb_desc_13_axuser_14_reg),
                              .uc2rb_desc_13_axuser_15_reg(uc2rb_desc_13_axuser_15_reg),
                              .uc2rb_desc_13_wuser_0_reg(uc2rb_desc_13_wuser_0_reg),
                              .uc2rb_desc_13_wuser_1_reg(uc2rb_desc_13_wuser_1_reg),
                              .uc2rb_desc_13_wuser_2_reg(uc2rb_desc_13_wuser_2_reg),
                              .uc2rb_desc_13_wuser_3_reg(uc2rb_desc_13_wuser_3_reg),
                              .uc2rb_desc_13_wuser_4_reg(uc2rb_desc_13_wuser_4_reg),
                              .uc2rb_desc_13_wuser_5_reg(uc2rb_desc_13_wuser_5_reg),
                              .uc2rb_desc_13_wuser_6_reg(uc2rb_desc_13_wuser_6_reg),
                              .uc2rb_desc_13_wuser_7_reg(uc2rb_desc_13_wuser_7_reg),
                              .uc2rb_desc_13_wuser_8_reg(uc2rb_desc_13_wuser_8_reg),
                              .uc2rb_desc_13_wuser_9_reg(uc2rb_desc_13_wuser_9_reg),
                              .uc2rb_desc_13_wuser_10_reg(uc2rb_desc_13_wuser_10_reg),
                              .uc2rb_desc_13_wuser_11_reg(uc2rb_desc_13_wuser_11_reg),
                              .uc2rb_desc_13_wuser_12_reg(uc2rb_desc_13_wuser_12_reg),
                              .uc2rb_desc_13_wuser_13_reg(uc2rb_desc_13_wuser_13_reg),
                              .uc2rb_desc_13_wuser_14_reg(uc2rb_desc_13_wuser_14_reg),
                              .uc2rb_desc_13_wuser_15_reg(uc2rb_desc_13_wuser_15_reg),
                              .uc2rb_desc_14_txn_type_reg(uc2rb_desc_14_txn_type_reg),
                              .uc2rb_desc_14_size_reg(uc2rb_desc_14_size_reg),
                              .uc2rb_desc_14_data_offset_reg(uc2rb_desc_14_data_offset_reg),
                              .uc2rb_desc_14_axsize_reg(uc2rb_desc_14_axsize_reg),
                              .uc2rb_desc_14_attr_reg(uc2rb_desc_14_attr_reg),
                              .uc2rb_desc_14_axaddr_0_reg(uc2rb_desc_14_axaddr_0_reg),
                              .uc2rb_desc_14_axaddr_1_reg(uc2rb_desc_14_axaddr_1_reg),
                              .uc2rb_desc_14_axaddr_2_reg(uc2rb_desc_14_axaddr_2_reg),
                              .uc2rb_desc_14_axaddr_3_reg(uc2rb_desc_14_axaddr_3_reg),
                              .uc2rb_desc_14_axid_0_reg(uc2rb_desc_14_axid_0_reg),
                              .uc2rb_desc_14_axid_1_reg(uc2rb_desc_14_axid_1_reg),
                              .uc2rb_desc_14_axid_2_reg(uc2rb_desc_14_axid_2_reg),
                              .uc2rb_desc_14_axid_3_reg(uc2rb_desc_14_axid_3_reg),
                              .uc2rb_desc_14_axuser_0_reg(uc2rb_desc_14_axuser_0_reg),
                              .uc2rb_desc_14_axuser_1_reg(uc2rb_desc_14_axuser_1_reg),
                              .uc2rb_desc_14_axuser_2_reg(uc2rb_desc_14_axuser_2_reg),
                              .uc2rb_desc_14_axuser_3_reg(uc2rb_desc_14_axuser_3_reg),
                              .uc2rb_desc_14_axuser_4_reg(uc2rb_desc_14_axuser_4_reg),
                              .uc2rb_desc_14_axuser_5_reg(uc2rb_desc_14_axuser_5_reg),
                              .uc2rb_desc_14_axuser_6_reg(uc2rb_desc_14_axuser_6_reg),
                              .uc2rb_desc_14_axuser_7_reg(uc2rb_desc_14_axuser_7_reg),
                              .uc2rb_desc_14_axuser_8_reg(uc2rb_desc_14_axuser_8_reg),
                              .uc2rb_desc_14_axuser_9_reg(uc2rb_desc_14_axuser_9_reg),
                              .uc2rb_desc_14_axuser_10_reg(uc2rb_desc_14_axuser_10_reg),
                              .uc2rb_desc_14_axuser_11_reg(uc2rb_desc_14_axuser_11_reg),
                              .uc2rb_desc_14_axuser_12_reg(uc2rb_desc_14_axuser_12_reg),
                              .uc2rb_desc_14_axuser_13_reg(uc2rb_desc_14_axuser_13_reg),
                              .uc2rb_desc_14_axuser_14_reg(uc2rb_desc_14_axuser_14_reg),
                              .uc2rb_desc_14_axuser_15_reg(uc2rb_desc_14_axuser_15_reg),
                              .uc2rb_desc_14_wuser_0_reg(uc2rb_desc_14_wuser_0_reg),
                              .uc2rb_desc_14_wuser_1_reg(uc2rb_desc_14_wuser_1_reg),
                              .uc2rb_desc_14_wuser_2_reg(uc2rb_desc_14_wuser_2_reg),
                              .uc2rb_desc_14_wuser_3_reg(uc2rb_desc_14_wuser_3_reg),
                              .uc2rb_desc_14_wuser_4_reg(uc2rb_desc_14_wuser_4_reg),
                              .uc2rb_desc_14_wuser_5_reg(uc2rb_desc_14_wuser_5_reg),
                              .uc2rb_desc_14_wuser_6_reg(uc2rb_desc_14_wuser_6_reg),
                              .uc2rb_desc_14_wuser_7_reg(uc2rb_desc_14_wuser_7_reg),
                              .uc2rb_desc_14_wuser_8_reg(uc2rb_desc_14_wuser_8_reg),
                              .uc2rb_desc_14_wuser_9_reg(uc2rb_desc_14_wuser_9_reg),
                              .uc2rb_desc_14_wuser_10_reg(uc2rb_desc_14_wuser_10_reg),
                              .uc2rb_desc_14_wuser_11_reg(uc2rb_desc_14_wuser_11_reg),
                              .uc2rb_desc_14_wuser_12_reg(uc2rb_desc_14_wuser_12_reg),
                              .uc2rb_desc_14_wuser_13_reg(uc2rb_desc_14_wuser_13_reg),
                              .uc2rb_desc_14_wuser_14_reg(uc2rb_desc_14_wuser_14_reg),
                              .uc2rb_desc_14_wuser_15_reg(uc2rb_desc_14_wuser_15_reg),
                              .uc2rb_desc_15_txn_type_reg(uc2rb_desc_15_txn_type_reg),
                              .uc2rb_desc_15_size_reg(uc2rb_desc_15_size_reg),
                              .uc2rb_desc_15_data_offset_reg(uc2rb_desc_15_data_offset_reg),
                              .uc2rb_desc_15_axsize_reg(uc2rb_desc_15_axsize_reg),
                              .uc2rb_desc_15_attr_reg(uc2rb_desc_15_attr_reg),
                              .uc2rb_desc_15_axaddr_0_reg(uc2rb_desc_15_axaddr_0_reg),
                              .uc2rb_desc_15_axaddr_1_reg(uc2rb_desc_15_axaddr_1_reg),
                              .uc2rb_desc_15_axaddr_2_reg(uc2rb_desc_15_axaddr_2_reg),
                              .uc2rb_desc_15_axaddr_3_reg(uc2rb_desc_15_axaddr_3_reg),
                              .uc2rb_desc_15_axid_0_reg(uc2rb_desc_15_axid_0_reg),
                              .uc2rb_desc_15_axid_1_reg(uc2rb_desc_15_axid_1_reg),
                              .uc2rb_desc_15_axid_2_reg(uc2rb_desc_15_axid_2_reg),
                              .uc2rb_desc_15_axid_3_reg(uc2rb_desc_15_axid_3_reg),
                              .uc2rb_desc_15_axuser_0_reg(uc2rb_desc_15_axuser_0_reg),
                              .uc2rb_desc_15_axuser_1_reg(uc2rb_desc_15_axuser_1_reg),
                              .uc2rb_desc_15_axuser_2_reg(uc2rb_desc_15_axuser_2_reg),
                              .uc2rb_desc_15_axuser_3_reg(uc2rb_desc_15_axuser_3_reg),
                              .uc2rb_desc_15_axuser_4_reg(uc2rb_desc_15_axuser_4_reg),
                              .uc2rb_desc_15_axuser_5_reg(uc2rb_desc_15_axuser_5_reg),
                              .uc2rb_desc_15_axuser_6_reg(uc2rb_desc_15_axuser_6_reg),
                              .uc2rb_desc_15_axuser_7_reg(uc2rb_desc_15_axuser_7_reg),
                              .uc2rb_desc_15_axuser_8_reg(uc2rb_desc_15_axuser_8_reg),
                              .uc2rb_desc_15_axuser_9_reg(uc2rb_desc_15_axuser_9_reg),
                              .uc2rb_desc_15_axuser_10_reg(uc2rb_desc_15_axuser_10_reg),
                              .uc2rb_desc_15_axuser_11_reg(uc2rb_desc_15_axuser_11_reg),
                              .uc2rb_desc_15_axuser_12_reg(uc2rb_desc_15_axuser_12_reg),
                              .uc2rb_desc_15_axuser_13_reg(uc2rb_desc_15_axuser_13_reg),
                              .uc2rb_desc_15_axuser_14_reg(uc2rb_desc_15_axuser_14_reg),
                              .uc2rb_desc_15_axuser_15_reg(uc2rb_desc_15_axuser_15_reg),
                              .uc2rb_desc_15_wuser_0_reg(uc2rb_desc_15_wuser_0_reg),
                              .uc2rb_desc_15_wuser_1_reg(uc2rb_desc_15_wuser_1_reg),
                              .uc2rb_desc_15_wuser_2_reg(uc2rb_desc_15_wuser_2_reg),
                              .uc2rb_desc_15_wuser_3_reg(uc2rb_desc_15_wuser_3_reg),
                              .uc2rb_desc_15_wuser_4_reg(uc2rb_desc_15_wuser_4_reg),
                              .uc2rb_desc_15_wuser_5_reg(uc2rb_desc_15_wuser_5_reg),
                              .uc2rb_desc_15_wuser_6_reg(uc2rb_desc_15_wuser_6_reg),
                              .uc2rb_desc_15_wuser_7_reg(uc2rb_desc_15_wuser_7_reg),
                              .uc2rb_desc_15_wuser_8_reg(uc2rb_desc_15_wuser_8_reg),
                              .uc2rb_desc_15_wuser_9_reg(uc2rb_desc_15_wuser_9_reg),
                              .uc2rb_desc_15_wuser_10_reg(uc2rb_desc_15_wuser_10_reg),
                              .uc2rb_desc_15_wuser_11_reg(uc2rb_desc_15_wuser_11_reg),
                              .uc2rb_desc_15_wuser_12_reg(uc2rb_desc_15_wuser_12_reg),
                              .uc2rb_desc_15_wuser_13_reg(uc2rb_desc_15_wuser_13_reg),
                              .uc2rb_desc_15_wuser_14_reg(uc2rb_desc_15_wuser_14_reg),
                              .uc2rb_desc_15_wuser_15_reg(uc2rb_desc_15_wuser_15_reg),
                              .uc2rb_intr_error_status_reg_we(uc2rb_intr_error_status_reg_we),
                              .uc2rb_ownership_reg_we(uc2rb_ownership_reg_we),
                              .uc2rb_intr_txn_avail_status_reg_we(uc2rb_intr_txn_avail_status_reg_we),
                              .uc2rb_intr_comp_status_reg_we(uc2rb_intr_comp_status_reg_we),
                              .uc2rb_status_busy_reg_we(uc2rb_status_busy_reg_we),
                              .uc2rb_resp_fifo_free_level_reg_we(uc2rb_resp_fifo_free_level_reg_we),
                              .uc2rb_desc_0_txn_type_reg_we(uc2rb_desc_0_txn_type_reg_we),
                              .uc2rb_desc_0_size_reg_we(uc2rb_desc_0_size_reg_we),
                              .uc2rb_desc_0_data_offset_reg_we(uc2rb_desc_0_data_offset_reg_we),
                              .uc2rb_desc_0_axsize_reg_we(uc2rb_desc_0_axsize_reg_we),
                              .uc2rb_desc_0_attr_reg_we(uc2rb_desc_0_attr_reg_we),
                              .uc2rb_desc_0_axaddr_0_reg_we(uc2rb_desc_0_axaddr_0_reg_we),
                              .uc2rb_desc_0_axaddr_1_reg_we(uc2rb_desc_0_axaddr_1_reg_we),
                              .uc2rb_desc_0_axaddr_2_reg_we(uc2rb_desc_0_axaddr_2_reg_we),
                              .uc2rb_desc_0_axaddr_3_reg_we(uc2rb_desc_0_axaddr_3_reg_we),
                              .uc2rb_desc_0_axid_0_reg_we(uc2rb_desc_0_axid_0_reg_we),
                              .uc2rb_desc_0_axid_1_reg_we(uc2rb_desc_0_axid_1_reg_we),
                              .uc2rb_desc_0_axid_2_reg_we(uc2rb_desc_0_axid_2_reg_we),
                              .uc2rb_desc_0_axid_3_reg_we(uc2rb_desc_0_axid_3_reg_we),
                              .uc2rb_desc_0_axuser_0_reg_we(uc2rb_desc_0_axuser_0_reg_we),
                              .uc2rb_desc_0_axuser_1_reg_we(uc2rb_desc_0_axuser_1_reg_we),
                              .uc2rb_desc_0_axuser_2_reg_we(uc2rb_desc_0_axuser_2_reg_we),
                              .uc2rb_desc_0_axuser_3_reg_we(uc2rb_desc_0_axuser_3_reg_we),
                              .uc2rb_desc_0_axuser_4_reg_we(uc2rb_desc_0_axuser_4_reg_we),
                              .uc2rb_desc_0_axuser_5_reg_we(uc2rb_desc_0_axuser_5_reg_we),
                              .uc2rb_desc_0_axuser_6_reg_we(uc2rb_desc_0_axuser_6_reg_we),
                              .uc2rb_desc_0_axuser_7_reg_we(uc2rb_desc_0_axuser_7_reg_we),
                              .uc2rb_desc_0_axuser_8_reg_we(uc2rb_desc_0_axuser_8_reg_we),
                              .uc2rb_desc_0_axuser_9_reg_we(uc2rb_desc_0_axuser_9_reg_we),
                              .uc2rb_desc_0_axuser_10_reg_we(uc2rb_desc_0_axuser_10_reg_we),
                              .uc2rb_desc_0_axuser_11_reg_we(uc2rb_desc_0_axuser_11_reg_we),
                              .uc2rb_desc_0_axuser_12_reg_we(uc2rb_desc_0_axuser_12_reg_we),
                              .uc2rb_desc_0_axuser_13_reg_we(uc2rb_desc_0_axuser_13_reg_we),
                              .uc2rb_desc_0_axuser_14_reg_we(uc2rb_desc_0_axuser_14_reg_we),
                              .uc2rb_desc_0_axuser_15_reg_we(uc2rb_desc_0_axuser_15_reg_we),
                              .uc2rb_desc_0_wuser_0_reg_we(uc2rb_desc_0_wuser_0_reg_we),
                              .uc2rb_desc_0_wuser_1_reg_we(uc2rb_desc_0_wuser_1_reg_we),
                              .uc2rb_desc_0_wuser_2_reg_we(uc2rb_desc_0_wuser_2_reg_we),
                              .uc2rb_desc_0_wuser_3_reg_we(uc2rb_desc_0_wuser_3_reg_we),
                              .uc2rb_desc_0_wuser_4_reg_we(uc2rb_desc_0_wuser_4_reg_we),
                              .uc2rb_desc_0_wuser_5_reg_we(uc2rb_desc_0_wuser_5_reg_we),
                              .uc2rb_desc_0_wuser_6_reg_we(uc2rb_desc_0_wuser_6_reg_we),
                              .uc2rb_desc_0_wuser_7_reg_we(uc2rb_desc_0_wuser_7_reg_we),
                              .uc2rb_desc_0_wuser_8_reg_we(uc2rb_desc_0_wuser_8_reg_we),
                              .uc2rb_desc_0_wuser_9_reg_we(uc2rb_desc_0_wuser_9_reg_we),
                              .uc2rb_desc_0_wuser_10_reg_we(uc2rb_desc_0_wuser_10_reg_we),
                              .uc2rb_desc_0_wuser_11_reg_we(uc2rb_desc_0_wuser_11_reg_we),
                              .uc2rb_desc_0_wuser_12_reg_we(uc2rb_desc_0_wuser_12_reg_we),
                              .uc2rb_desc_0_wuser_13_reg_we(uc2rb_desc_0_wuser_13_reg_we),
                              .uc2rb_desc_0_wuser_14_reg_we(uc2rb_desc_0_wuser_14_reg_we),
                              .uc2rb_desc_0_wuser_15_reg_we(uc2rb_desc_0_wuser_15_reg_we),
                              .uc2rb_desc_1_txn_type_reg_we(uc2rb_desc_1_txn_type_reg_we),
                              .uc2rb_desc_1_size_reg_we(uc2rb_desc_1_size_reg_we),
                              .uc2rb_desc_1_data_offset_reg_we(uc2rb_desc_1_data_offset_reg_we),
                              .uc2rb_desc_1_axsize_reg_we(uc2rb_desc_1_axsize_reg_we),
                              .uc2rb_desc_1_attr_reg_we(uc2rb_desc_1_attr_reg_we),
                              .uc2rb_desc_1_axaddr_0_reg_we(uc2rb_desc_1_axaddr_0_reg_we),
                              .uc2rb_desc_1_axaddr_1_reg_we(uc2rb_desc_1_axaddr_1_reg_we),
                              .uc2rb_desc_1_axaddr_2_reg_we(uc2rb_desc_1_axaddr_2_reg_we),
                              .uc2rb_desc_1_axaddr_3_reg_we(uc2rb_desc_1_axaddr_3_reg_we),
                              .uc2rb_desc_1_axid_0_reg_we(uc2rb_desc_1_axid_0_reg_we),
                              .uc2rb_desc_1_axid_1_reg_we(uc2rb_desc_1_axid_1_reg_we),
                              .uc2rb_desc_1_axid_2_reg_we(uc2rb_desc_1_axid_2_reg_we),
                              .uc2rb_desc_1_axid_3_reg_we(uc2rb_desc_1_axid_3_reg_we),
                              .uc2rb_desc_1_axuser_0_reg_we(uc2rb_desc_1_axuser_0_reg_we),
                              .uc2rb_desc_1_axuser_1_reg_we(uc2rb_desc_1_axuser_1_reg_we),
                              .uc2rb_desc_1_axuser_2_reg_we(uc2rb_desc_1_axuser_2_reg_we),
                              .uc2rb_desc_1_axuser_3_reg_we(uc2rb_desc_1_axuser_3_reg_we),
                              .uc2rb_desc_1_axuser_4_reg_we(uc2rb_desc_1_axuser_4_reg_we),
                              .uc2rb_desc_1_axuser_5_reg_we(uc2rb_desc_1_axuser_5_reg_we),
                              .uc2rb_desc_1_axuser_6_reg_we(uc2rb_desc_1_axuser_6_reg_we),
                              .uc2rb_desc_1_axuser_7_reg_we(uc2rb_desc_1_axuser_7_reg_we),
                              .uc2rb_desc_1_axuser_8_reg_we(uc2rb_desc_1_axuser_8_reg_we),
                              .uc2rb_desc_1_axuser_9_reg_we(uc2rb_desc_1_axuser_9_reg_we),
                              .uc2rb_desc_1_axuser_10_reg_we(uc2rb_desc_1_axuser_10_reg_we),
                              .uc2rb_desc_1_axuser_11_reg_we(uc2rb_desc_1_axuser_11_reg_we),
                              .uc2rb_desc_1_axuser_12_reg_we(uc2rb_desc_1_axuser_12_reg_we),
                              .uc2rb_desc_1_axuser_13_reg_we(uc2rb_desc_1_axuser_13_reg_we),
                              .uc2rb_desc_1_axuser_14_reg_we(uc2rb_desc_1_axuser_14_reg_we),
                              .uc2rb_desc_1_axuser_15_reg_we(uc2rb_desc_1_axuser_15_reg_we),
                              .uc2rb_desc_1_wuser_0_reg_we(uc2rb_desc_1_wuser_0_reg_we),
                              .uc2rb_desc_1_wuser_1_reg_we(uc2rb_desc_1_wuser_1_reg_we),
                              .uc2rb_desc_1_wuser_2_reg_we(uc2rb_desc_1_wuser_2_reg_we),
                              .uc2rb_desc_1_wuser_3_reg_we(uc2rb_desc_1_wuser_3_reg_we),
                              .uc2rb_desc_1_wuser_4_reg_we(uc2rb_desc_1_wuser_4_reg_we),
                              .uc2rb_desc_1_wuser_5_reg_we(uc2rb_desc_1_wuser_5_reg_we),
                              .uc2rb_desc_1_wuser_6_reg_we(uc2rb_desc_1_wuser_6_reg_we),
                              .uc2rb_desc_1_wuser_7_reg_we(uc2rb_desc_1_wuser_7_reg_we),
                              .uc2rb_desc_1_wuser_8_reg_we(uc2rb_desc_1_wuser_8_reg_we),
                              .uc2rb_desc_1_wuser_9_reg_we(uc2rb_desc_1_wuser_9_reg_we),
                              .uc2rb_desc_1_wuser_10_reg_we(uc2rb_desc_1_wuser_10_reg_we),
                              .uc2rb_desc_1_wuser_11_reg_we(uc2rb_desc_1_wuser_11_reg_we),
                              .uc2rb_desc_1_wuser_12_reg_we(uc2rb_desc_1_wuser_12_reg_we),
                              .uc2rb_desc_1_wuser_13_reg_we(uc2rb_desc_1_wuser_13_reg_we),
                              .uc2rb_desc_1_wuser_14_reg_we(uc2rb_desc_1_wuser_14_reg_we),
                              .uc2rb_desc_1_wuser_15_reg_we(uc2rb_desc_1_wuser_15_reg_we),
                              .uc2rb_desc_2_txn_type_reg_we(uc2rb_desc_2_txn_type_reg_we),
                              .uc2rb_desc_2_size_reg_we(uc2rb_desc_2_size_reg_we),
                              .uc2rb_desc_2_data_offset_reg_we(uc2rb_desc_2_data_offset_reg_we),
                              .uc2rb_desc_2_axsize_reg_we(uc2rb_desc_2_axsize_reg_we),
                              .uc2rb_desc_2_attr_reg_we(uc2rb_desc_2_attr_reg_we),
                              .uc2rb_desc_2_axaddr_0_reg_we(uc2rb_desc_2_axaddr_0_reg_we),
                              .uc2rb_desc_2_axaddr_1_reg_we(uc2rb_desc_2_axaddr_1_reg_we),
                              .uc2rb_desc_2_axaddr_2_reg_we(uc2rb_desc_2_axaddr_2_reg_we),
                              .uc2rb_desc_2_axaddr_3_reg_we(uc2rb_desc_2_axaddr_3_reg_we),
                              .uc2rb_desc_2_axid_0_reg_we(uc2rb_desc_2_axid_0_reg_we),
                              .uc2rb_desc_2_axid_1_reg_we(uc2rb_desc_2_axid_1_reg_we),
                              .uc2rb_desc_2_axid_2_reg_we(uc2rb_desc_2_axid_2_reg_we),
                              .uc2rb_desc_2_axid_3_reg_we(uc2rb_desc_2_axid_3_reg_we),
                              .uc2rb_desc_2_axuser_0_reg_we(uc2rb_desc_2_axuser_0_reg_we),
                              .uc2rb_desc_2_axuser_1_reg_we(uc2rb_desc_2_axuser_1_reg_we),
                              .uc2rb_desc_2_axuser_2_reg_we(uc2rb_desc_2_axuser_2_reg_we),
                              .uc2rb_desc_2_axuser_3_reg_we(uc2rb_desc_2_axuser_3_reg_we),
                              .uc2rb_desc_2_axuser_4_reg_we(uc2rb_desc_2_axuser_4_reg_we),
                              .uc2rb_desc_2_axuser_5_reg_we(uc2rb_desc_2_axuser_5_reg_we),
                              .uc2rb_desc_2_axuser_6_reg_we(uc2rb_desc_2_axuser_6_reg_we),
                              .uc2rb_desc_2_axuser_7_reg_we(uc2rb_desc_2_axuser_7_reg_we),
                              .uc2rb_desc_2_axuser_8_reg_we(uc2rb_desc_2_axuser_8_reg_we),
                              .uc2rb_desc_2_axuser_9_reg_we(uc2rb_desc_2_axuser_9_reg_we),
                              .uc2rb_desc_2_axuser_10_reg_we(uc2rb_desc_2_axuser_10_reg_we),
                              .uc2rb_desc_2_axuser_11_reg_we(uc2rb_desc_2_axuser_11_reg_we),
                              .uc2rb_desc_2_axuser_12_reg_we(uc2rb_desc_2_axuser_12_reg_we),
                              .uc2rb_desc_2_axuser_13_reg_we(uc2rb_desc_2_axuser_13_reg_we),
                              .uc2rb_desc_2_axuser_14_reg_we(uc2rb_desc_2_axuser_14_reg_we),
                              .uc2rb_desc_2_axuser_15_reg_we(uc2rb_desc_2_axuser_15_reg_we),
                              .uc2rb_desc_2_wuser_0_reg_we(uc2rb_desc_2_wuser_0_reg_we),
                              .uc2rb_desc_2_wuser_1_reg_we(uc2rb_desc_2_wuser_1_reg_we),
                              .uc2rb_desc_2_wuser_2_reg_we(uc2rb_desc_2_wuser_2_reg_we),
                              .uc2rb_desc_2_wuser_3_reg_we(uc2rb_desc_2_wuser_3_reg_we),
                              .uc2rb_desc_2_wuser_4_reg_we(uc2rb_desc_2_wuser_4_reg_we),
                              .uc2rb_desc_2_wuser_5_reg_we(uc2rb_desc_2_wuser_5_reg_we),
                              .uc2rb_desc_2_wuser_6_reg_we(uc2rb_desc_2_wuser_6_reg_we),
                              .uc2rb_desc_2_wuser_7_reg_we(uc2rb_desc_2_wuser_7_reg_we),
                              .uc2rb_desc_2_wuser_8_reg_we(uc2rb_desc_2_wuser_8_reg_we),
                              .uc2rb_desc_2_wuser_9_reg_we(uc2rb_desc_2_wuser_9_reg_we),
                              .uc2rb_desc_2_wuser_10_reg_we(uc2rb_desc_2_wuser_10_reg_we),
                              .uc2rb_desc_2_wuser_11_reg_we(uc2rb_desc_2_wuser_11_reg_we),
                              .uc2rb_desc_2_wuser_12_reg_we(uc2rb_desc_2_wuser_12_reg_we),
                              .uc2rb_desc_2_wuser_13_reg_we(uc2rb_desc_2_wuser_13_reg_we),
                              .uc2rb_desc_2_wuser_14_reg_we(uc2rb_desc_2_wuser_14_reg_we),
                              .uc2rb_desc_2_wuser_15_reg_we(uc2rb_desc_2_wuser_15_reg_we),
                              .uc2rb_desc_3_txn_type_reg_we(uc2rb_desc_3_txn_type_reg_we),
                              .uc2rb_desc_3_size_reg_we(uc2rb_desc_3_size_reg_we),
                              .uc2rb_desc_3_data_offset_reg_we(uc2rb_desc_3_data_offset_reg_we),
                              .uc2rb_desc_3_axsize_reg_we(uc2rb_desc_3_axsize_reg_we),
                              .uc2rb_desc_3_attr_reg_we(uc2rb_desc_3_attr_reg_we),
                              .uc2rb_desc_3_axaddr_0_reg_we(uc2rb_desc_3_axaddr_0_reg_we),
                              .uc2rb_desc_3_axaddr_1_reg_we(uc2rb_desc_3_axaddr_1_reg_we),
                              .uc2rb_desc_3_axaddr_2_reg_we(uc2rb_desc_3_axaddr_2_reg_we),
                              .uc2rb_desc_3_axaddr_3_reg_we(uc2rb_desc_3_axaddr_3_reg_we),
                              .uc2rb_desc_3_axid_0_reg_we(uc2rb_desc_3_axid_0_reg_we),
                              .uc2rb_desc_3_axid_1_reg_we(uc2rb_desc_3_axid_1_reg_we),
                              .uc2rb_desc_3_axid_2_reg_we(uc2rb_desc_3_axid_2_reg_we),
                              .uc2rb_desc_3_axid_3_reg_we(uc2rb_desc_3_axid_3_reg_we),
                              .uc2rb_desc_3_axuser_0_reg_we(uc2rb_desc_3_axuser_0_reg_we),
                              .uc2rb_desc_3_axuser_1_reg_we(uc2rb_desc_3_axuser_1_reg_we),
                              .uc2rb_desc_3_axuser_2_reg_we(uc2rb_desc_3_axuser_2_reg_we),
                              .uc2rb_desc_3_axuser_3_reg_we(uc2rb_desc_3_axuser_3_reg_we),
                              .uc2rb_desc_3_axuser_4_reg_we(uc2rb_desc_3_axuser_4_reg_we),
                              .uc2rb_desc_3_axuser_5_reg_we(uc2rb_desc_3_axuser_5_reg_we),
                              .uc2rb_desc_3_axuser_6_reg_we(uc2rb_desc_3_axuser_6_reg_we),
                              .uc2rb_desc_3_axuser_7_reg_we(uc2rb_desc_3_axuser_7_reg_we),
                              .uc2rb_desc_3_axuser_8_reg_we(uc2rb_desc_3_axuser_8_reg_we),
                              .uc2rb_desc_3_axuser_9_reg_we(uc2rb_desc_3_axuser_9_reg_we),
                              .uc2rb_desc_3_axuser_10_reg_we(uc2rb_desc_3_axuser_10_reg_we),
                              .uc2rb_desc_3_axuser_11_reg_we(uc2rb_desc_3_axuser_11_reg_we),
                              .uc2rb_desc_3_axuser_12_reg_we(uc2rb_desc_3_axuser_12_reg_we),
                              .uc2rb_desc_3_axuser_13_reg_we(uc2rb_desc_3_axuser_13_reg_we),
                              .uc2rb_desc_3_axuser_14_reg_we(uc2rb_desc_3_axuser_14_reg_we),
                              .uc2rb_desc_3_axuser_15_reg_we(uc2rb_desc_3_axuser_15_reg_we),
                              .uc2rb_desc_3_wuser_0_reg_we(uc2rb_desc_3_wuser_0_reg_we),
                              .uc2rb_desc_3_wuser_1_reg_we(uc2rb_desc_3_wuser_1_reg_we),
                              .uc2rb_desc_3_wuser_2_reg_we(uc2rb_desc_3_wuser_2_reg_we),
                              .uc2rb_desc_3_wuser_3_reg_we(uc2rb_desc_3_wuser_3_reg_we),
                              .uc2rb_desc_3_wuser_4_reg_we(uc2rb_desc_3_wuser_4_reg_we),
                              .uc2rb_desc_3_wuser_5_reg_we(uc2rb_desc_3_wuser_5_reg_we),
                              .uc2rb_desc_3_wuser_6_reg_we(uc2rb_desc_3_wuser_6_reg_we),
                              .uc2rb_desc_3_wuser_7_reg_we(uc2rb_desc_3_wuser_7_reg_we),
                              .uc2rb_desc_3_wuser_8_reg_we(uc2rb_desc_3_wuser_8_reg_we),
                              .uc2rb_desc_3_wuser_9_reg_we(uc2rb_desc_3_wuser_9_reg_we),
                              .uc2rb_desc_3_wuser_10_reg_we(uc2rb_desc_3_wuser_10_reg_we),
                              .uc2rb_desc_3_wuser_11_reg_we(uc2rb_desc_3_wuser_11_reg_we),
                              .uc2rb_desc_3_wuser_12_reg_we(uc2rb_desc_3_wuser_12_reg_we),
                              .uc2rb_desc_3_wuser_13_reg_we(uc2rb_desc_3_wuser_13_reg_we),
                              .uc2rb_desc_3_wuser_14_reg_we(uc2rb_desc_3_wuser_14_reg_we),
                              .uc2rb_desc_3_wuser_15_reg_we(uc2rb_desc_3_wuser_15_reg_we),
                              .uc2rb_desc_4_txn_type_reg_we(uc2rb_desc_4_txn_type_reg_we),
                              .uc2rb_desc_4_size_reg_we(uc2rb_desc_4_size_reg_we),
                              .uc2rb_desc_4_data_offset_reg_we(uc2rb_desc_4_data_offset_reg_we),
                              .uc2rb_desc_4_axsize_reg_we(uc2rb_desc_4_axsize_reg_we),
                              .uc2rb_desc_4_attr_reg_we(uc2rb_desc_4_attr_reg_we),
                              .uc2rb_desc_4_axaddr_0_reg_we(uc2rb_desc_4_axaddr_0_reg_we),
                              .uc2rb_desc_4_axaddr_1_reg_we(uc2rb_desc_4_axaddr_1_reg_we),
                              .uc2rb_desc_4_axaddr_2_reg_we(uc2rb_desc_4_axaddr_2_reg_we),
                              .uc2rb_desc_4_axaddr_3_reg_we(uc2rb_desc_4_axaddr_3_reg_we),
                              .uc2rb_desc_4_axid_0_reg_we(uc2rb_desc_4_axid_0_reg_we),
                              .uc2rb_desc_4_axid_1_reg_we(uc2rb_desc_4_axid_1_reg_we),
                              .uc2rb_desc_4_axid_2_reg_we(uc2rb_desc_4_axid_2_reg_we),
                              .uc2rb_desc_4_axid_3_reg_we(uc2rb_desc_4_axid_3_reg_we),
                              .uc2rb_desc_4_axuser_0_reg_we(uc2rb_desc_4_axuser_0_reg_we),
                              .uc2rb_desc_4_axuser_1_reg_we(uc2rb_desc_4_axuser_1_reg_we),
                              .uc2rb_desc_4_axuser_2_reg_we(uc2rb_desc_4_axuser_2_reg_we),
                              .uc2rb_desc_4_axuser_3_reg_we(uc2rb_desc_4_axuser_3_reg_we),
                              .uc2rb_desc_4_axuser_4_reg_we(uc2rb_desc_4_axuser_4_reg_we),
                              .uc2rb_desc_4_axuser_5_reg_we(uc2rb_desc_4_axuser_5_reg_we),
                              .uc2rb_desc_4_axuser_6_reg_we(uc2rb_desc_4_axuser_6_reg_we),
                              .uc2rb_desc_4_axuser_7_reg_we(uc2rb_desc_4_axuser_7_reg_we),
                              .uc2rb_desc_4_axuser_8_reg_we(uc2rb_desc_4_axuser_8_reg_we),
                              .uc2rb_desc_4_axuser_9_reg_we(uc2rb_desc_4_axuser_9_reg_we),
                              .uc2rb_desc_4_axuser_10_reg_we(uc2rb_desc_4_axuser_10_reg_we),
                              .uc2rb_desc_4_axuser_11_reg_we(uc2rb_desc_4_axuser_11_reg_we),
                              .uc2rb_desc_4_axuser_12_reg_we(uc2rb_desc_4_axuser_12_reg_we),
                              .uc2rb_desc_4_axuser_13_reg_we(uc2rb_desc_4_axuser_13_reg_we),
                              .uc2rb_desc_4_axuser_14_reg_we(uc2rb_desc_4_axuser_14_reg_we),
                              .uc2rb_desc_4_axuser_15_reg_we(uc2rb_desc_4_axuser_15_reg_we),
                              .uc2rb_desc_4_wuser_0_reg_we(uc2rb_desc_4_wuser_0_reg_we),
                              .uc2rb_desc_4_wuser_1_reg_we(uc2rb_desc_4_wuser_1_reg_we),
                              .uc2rb_desc_4_wuser_2_reg_we(uc2rb_desc_4_wuser_2_reg_we),
                              .uc2rb_desc_4_wuser_3_reg_we(uc2rb_desc_4_wuser_3_reg_we),
                              .uc2rb_desc_4_wuser_4_reg_we(uc2rb_desc_4_wuser_4_reg_we),
                              .uc2rb_desc_4_wuser_5_reg_we(uc2rb_desc_4_wuser_5_reg_we),
                              .uc2rb_desc_4_wuser_6_reg_we(uc2rb_desc_4_wuser_6_reg_we),
                              .uc2rb_desc_4_wuser_7_reg_we(uc2rb_desc_4_wuser_7_reg_we),
                              .uc2rb_desc_4_wuser_8_reg_we(uc2rb_desc_4_wuser_8_reg_we),
                              .uc2rb_desc_4_wuser_9_reg_we(uc2rb_desc_4_wuser_9_reg_we),
                              .uc2rb_desc_4_wuser_10_reg_we(uc2rb_desc_4_wuser_10_reg_we),
                              .uc2rb_desc_4_wuser_11_reg_we(uc2rb_desc_4_wuser_11_reg_we),
                              .uc2rb_desc_4_wuser_12_reg_we(uc2rb_desc_4_wuser_12_reg_we),
                              .uc2rb_desc_4_wuser_13_reg_we(uc2rb_desc_4_wuser_13_reg_we),
                              .uc2rb_desc_4_wuser_14_reg_we(uc2rb_desc_4_wuser_14_reg_we),
                              .uc2rb_desc_4_wuser_15_reg_we(uc2rb_desc_4_wuser_15_reg_we),
                              .uc2rb_desc_5_txn_type_reg_we(uc2rb_desc_5_txn_type_reg_we),
                              .uc2rb_desc_5_size_reg_we(uc2rb_desc_5_size_reg_we),
                              .uc2rb_desc_5_data_offset_reg_we(uc2rb_desc_5_data_offset_reg_we),
                              .uc2rb_desc_5_axsize_reg_we(uc2rb_desc_5_axsize_reg_we),
                              .uc2rb_desc_5_attr_reg_we(uc2rb_desc_5_attr_reg_we),
                              .uc2rb_desc_5_axaddr_0_reg_we(uc2rb_desc_5_axaddr_0_reg_we),
                              .uc2rb_desc_5_axaddr_1_reg_we(uc2rb_desc_5_axaddr_1_reg_we),
                              .uc2rb_desc_5_axaddr_2_reg_we(uc2rb_desc_5_axaddr_2_reg_we),
                              .uc2rb_desc_5_axaddr_3_reg_we(uc2rb_desc_5_axaddr_3_reg_we),
                              .uc2rb_desc_5_axid_0_reg_we(uc2rb_desc_5_axid_0_reg_we),
                              .uc2rb_desc_5_axid_1_reg_we(uc2rb_desc_5_axid_1_reg_we),
                              .uc2rb_desc_5_axid_2_reg_we(uc2rb_desc_5_axid_2_reg_we),
                              .uc2rb_desc_5_axid_3_reg_we(uc2rb_desc_5_axid_3_reg_we),
                              .uc2rb_desc_5_axuser_0_reg_we(uc2rb_desc_5_axuser_0_reg_we),
                              .uc2rb_desc_5_axuser_1_reg_we(uc2rb_desc_5_axuser_1_reg_we),
                              .uc2rb_desc_5_axuser_2_reg_we(uc2rb_desc_5_axuser_2_reg_we),
                              .uc2rb_desc_5_axuser_3_reg_we(uc2rb_desc_5_axuser_3_reg_we),
                              .uc2rb_desc_5_axuser_4_reg_we(uc2rb_desc_5_axuser_4_reg_we),
                              .uc2rb_desc_5_axuser_5_reg_we(uc2rb_desc_5_axuser_5_reg_we),
                              .uc2rb_desc_5_axuser_6_reg_we(uc2rb_desc_5_axuser_6_reg_we),
                              .uc2rb_desc_5_axuser_7_reg_we(uc2rb_desc_5_axuser_7_reg_we),
                              .uc2rb_desc_5_axuser_8_reg_we(uc2rb_desc_5_axuser_8_reg_we),
                              .uc2rb_desc_5_axuser_9_reg_we(uc2rb_desc_5_axuser_9_reg_we),
                              .uc2rb_desc_5_axuser_10_reg_we(uc2rb_desc_5_axuser_10_reg_we),
                              .uc2rb_desc_5_axuser_11_reg_we(uc2rb_desc_5_axuser_11_reg_we),
                              .uc2rb_desc_5_axuser_12_reg_we(uc2rb_desc_5_axuser_12_reg_we),
                              .uc2rb_desc_5_axuser_13_reg_we(uc2rb_desc_5_axuser_13_reg_we),
                              .uc2rb_desc_5_axuser_14_reg_we(uc2rb_desc_5_axuser_14_reg_we),
                              .uc2rb_desc_5_axuser_15_reg_we(uc2rb_desc_5_axuser_15_reg_we),
                              .uc2rb_desc_5_wuser_0_reg_we(uc2rb_desc_5_wuser_0_reg_we),
                              .uc2rb_desc_5_wuser_1_reg_we(uc2rb_desc_5_wuser_1_reg_we),
                              .uc2rb_desc_5_wuser_2_reg_we(uc2rb_desc_5_wuser_2_reg_we),
                              .uc2rb_desc_5_wuser_3_reg_we(uc2rb_desc_5_wuser_3_reg_we),
                              .uc2rb_desc_5_wuser_4_reg_we(uc2rb_desc_5_wuser_4_reg_we),
                              .uc2rb_desc_5_wuser_5_reg_we(uc2rb_desc_5_wuser_5_reg_we),
                              .uc2rb_desc_5_wuser_6_reg_we(uc2rb_desc_5_wuser_6_reg_we),
                              .uc2rb_desc_5_wuser_7_reg_we(uc2rb_desc_5_wuser_7_reg_we),
                              .uc2rb_desc_5_wuser_8_reg_we(uc2rb_desc_5_wuser_8_reg_we),
                              .uc2rb_desc_5_wuser_9_reg_we(uc2rb_desc_5_wuser_9_reg_we),
                              .uc2rb_desc_5_wuser_10_reg_we(uc2rb_desc_5_wuser_10_reg_we),
                              .uc2rb_desc_5_wuser_11_reg_we(uc2rb_desc_5_wuser_11_reg_we),
                              .uc2rb_desc_5_wuser_12_reg_we(uc2rb_desc_5_wuser_12_reg_we),
                              .uc2rb_desc_5_wuser_13_reg_we(uc2rb_desc_5_wuser_13_reg_we),
                              .uc2rb_desc_5_wuser_14_reg_we(uc2rb_desc_5_wuser_14_reg_we),
                              .uc2rb_desc_5_wuser_15_reg_we(uc2rb_desc_5_wuser_15_reg_we),
                              .uc2rb_desc_6_txn_type_reg_we(uc2rb_desc_6_txn_type_reg_we),
                              .uc2rb_desc_6_size_reg_we(uc2rb_desc_6_size_reg_we),
                              .uc2rb_desc_6_data_offset_reg_we(uc2rb_desc_6_data_offset_reg_we),
                              .uc2rb_desc_6_axsize_reg_we(uc2rb_desc_6_axsize_reg_we),
                              .uc2rb_desc_6_attr_reg_we(uc2rb_desc_6_attr_reg_we),
                              .uc2rb_desc_6_axaddr_0_reg_we(uc2rb_desc_6_axaddr_0_reg_we),
                              .uc2rb_desc_6_axaddr_1_reg_we(uc2rb_desc_6_axaddr_1_reg_we),
                              .uc2rb_desc_6_axaddr_2_reg_we(uc2rb_desc_6_axaddr_2_reg_we),
                              .uc2rb_desc_6_axaddr_3_reg_we(uc2rb_desc_6_axaddr_3_reg_we),
                              .uc2rb_desc_6_axid_0_reg_we(uc2rb_desc_6_axid_0_reg_we),
                              .uc2rb_desc_6_axid_1_reg_we(uc2rb_desc_6_axid_1_reg_we),
                              .uc2rb_desc_6_axid_2_reg_we(uc2rb_desc_6_axid_2_reg_we),
                              .uc2rb_desc_6_axid_3_reg_we(uc2rb_desc_6_axid_3_reg_we),
                              .uc2rb_desc_6_axuser_0_reg_we(uc2rb_desc_6_axuser_0_reg_we),
                              .uc2rb_desc_6_axuser_1_reg_we(uc2rb_desc_6_axuser_1_reg_we),
                              .uc2rb_desc_6_axuser_2_reg_we(uc2rb_desc_6_axuser_2_reg_we),
                              .uc2rb_desc_6_axuser_3_reg_we(uc2rb_desc_6_axuser_3_reg_we),
                              .uc2rb_desc_6_axuser_4_reg_we(uc2rb_desc_6_axuser_4_reg_we),
                              .uc2rb_desc_6_axuser_5_reg_we(uc2rb_desc_6_axuser_5_reg_we),
                              .uc2rb_desc_6_axuser_6_reg_we(uc2rb_desc_6_axuser_6_reg_we),
                              .uc2rb_desc_6_axuser_7_reg_we(uc2rb_desc_6_axuser_7_reg_we),
                              .uc2rb_desc_6_axuser_8_reg_we(uc2rb_desc_6_axuser_8_reg_we),
                              .uc2rb_desc_6_axuser_9_reg_we(uc2rb_desc_6_axuser_9_reg_we),
                              .uc2rb_desc_6_axuser_10_reg_we(uc2rb_desc_6_axuser_10_reg_we),
                              .uc2rb_desc_6_axuser_11_reg_we(uc2rb_desc_6_axuser_11_reg_we),
                              .uc2rb_desc_6_axuser_12_reg_we(uc2rb_desc_6_axuser_12_reg_we),
                              .uc2rb_desc_6_axuser_13_reg_we(uc2rb_desc_6_axuser_13_reg_we),
                              .uc2rb_desc_6_axuser_14_reg_we(uc2rb_desc_6_axuser_14_reg_we),
                              .uc2rb_desc_6_axuser_15_reg_we(uc2rb_desc_6_axuser_15_reg_we),
                              .uc2rb_desc_6_wuser_0_reg_we(uc2rb_desc_6_wuser_0_reg_we),
                              .uc2rb_desc_6_wuser_1_reg_we(uc2rb_desc_6_wuser_1_reg_we),
                              .uc2rb_desc_6_wuser_2_reg_we(uc2rb_desc_6_wuser_2_reg_we),
                              .uc2rb_desc_6_wuser_3_reg_we(uc2rb_desc_6_wuser_3_reg_we),
                              .uc2rb_desc_6_wuser_4_reg_we(uc2rb_desc_6_wuser_4_reg_we),
                              .uc2rb_desc_6_wuser_5_reg_we(uc2rb_desc_6_wuser_5_reg_we),
                              .uc2rb_desc_6_wuser_6_reg_we(uc2rb_desc_6_wuser_6_reg_we),
                              .uc2rb_desc_6_wuser_7_reg_we(uc2rb_desc_6_wuser_7_reg_we),
                              .uc2rb_desc_6_wuser_8_reg_we(uc2rb_desc_6_wuser_8_reg_we),
                              .uc2rb_desc_6_wuser_9_reg_we(uc2rb_desc_6_wuser_9_reg_we),
                              .uc2rb_desc_6_wuser_10_reg_we(uc2rb_desc_6_wuser_10_reg_we),
                              .uc2rb_desc_6_wuser_11_reg_we(uc2rb_desc_6_wuser_11_reg_we),
                              .uc2rb_desc_6_wuser_12_reg_we(uc2rb_desc_6_wuser_12_reg_we),
                              .uc2rb_desc_6_wuser_13_reg_we(uc2rb_desc_6_wuser_13_reg_we),
                              .uc2rb_desc_6_wuser_14_reg_we(uc2rb_desc_6_wuser_14_reg_we),
                              .uc2rb_desc_6_wuser_15_reg_we(uc2rb_desc_6_wuser_15_reg_we),
                              .uc2rb_desc_7_txn_type_reg_we(uc2rb_desc_7_txn_type_reg_we),
                              .uc2rb_desc_7_size_reg_we(uc2rb_desc_7_size_reg_we),
                              .uc2rb_desc_7_data_offset_reg_we(uc2rb_desc_7_data_offset_reg_we),
                              .uc2rb_desc_7_axsize_reg_we(uc2rb_desc_7_axsize_reg_we),
                              .uc2rb_desc_7_attr_reg_we(uc2rb_desc_7_attr_reg_we),
                              .uc2rb_desc_7_axaddr_0_reg_we(uc2rb_desc_7_axaddr_0_reg_we),
                              .uc2rb_desc_7_axaddr_1_reg_we(uc2rb_desc_7_axaddr_1_reg_we),
                              .uc2rb_desc_7_axaddr_2_reg_we(uc2rb_desc_7_axaddr_2_reg_we),
                              .uc2rb_desc_7_axaddr_3_reg_we(uc2rb_desc_7_axaddr_3_reg_we),
                              .uc2rb_desc_7_axid_0_reg_we(uc2rb_desc_7_axid_0_reg_we),
                              .uc2rb_desc_7_axid_1_reg_we(uc2rb_desc_7_axid_1_reg_we),
                              .uc2rb_desc_7_axid_2_reg_we(uc2rb_desc_7_axid_2_reg_we),
                              .uc2rb_desc_7_axid_3_reg_we(uc2rb_desc_7_axid_3_reg_we),
                              .uc2rb_desc_7_axuser_0_reg_we(uc2rb_desc_7_axuser_0_reg_we),
                              .uc2rb_desc_7_axuser_1_reg_we(uc2rb_desc_7_axuser_1_reg_we),
                              .uc2rb_desc_7_axuser_2_reg_we(uc2rb_desc_7_axuser_2_reg_we),
                              .uc2rb_desc_7_axuser_3_reg_we(uc2rb_desc_7_axuser_3_reg_we),
                              .uc2rb_desc_7_axuser_4_reg_we(uc2rb_desc_7_axuser_4_reg_we),
                              .uc2rb_desc_7_axuser_5_reg_we(uc2rb_desc_7_axuser_5_reg_we),
                              .uc2rb_desc_7_axuser_6_reg_we(uc2rb_desc_7_axuser_6_reg_we),
                              .uc2rb_desc_7_axuser_7_reg_we(uc2rb_desc_7_axuser_7_reg_we),
                              .uc2rb_desc_7_axuser_8_reg_we(uc2rb_desc_7_axuser_8_reg_we),
                              .uc2rb_desc_7_axuser_9_reg_we(uc2rb_desc_7_axuser_9_reg_we),
                              .uc2rb_desc_7_axuser_10_reg_we(uc2rb_desc_7_axuser_10_reg_we),
                              .uc2rb_desc_7_axuser_11_reg_we(uc2rb_desc_7_axuser_11_reg_we),
                              .uc2rb_desc_7_axuser_12_reg_we(uc2rb_desc_7_axuser_12_reg_we),
                              .uc2rb_desc_7_axuser_13_reg_we(uc2rb_desc_7_axuser_13_reg_we),
                              .uc2rb_desc_7_axuser_14_reg_we(uc2rb_desc_7_axuser_14_reg_we),
                              .uc2rb_desc_7_axuser_15_reg_we(uc2rb_desc_7_axuser_15_reg_we),
                              .uc2rb_desc_7_wuser_0_reg_we(uc2rb_desc_7_wuser_0_reg_we),
                              .uc2rb_desc_7_wuser_1_reg_we(uc2rb_desc_7_wuser_1_reg_we),
                              .uc2rb_desc_7_wuser_2_reg_we(uc2rb_desc_7_wuser_2_reg_we),
                              .uc2rb_desc_7_wuser_3_reg_we(uc2rb_desc_7_wuser_3_reg_we),
                              .uc2rb_desc_7_wuser_4_reg_we(uc2rb_desc_7_wuser_4_reg_we),
                              .uc2rb_desc_7_wuser_5_reg_we(uc2rb_desc_7_wuser_5_reg_we),
                              .uc2rb_desc_7_wuser_6_reg_we(uc2rb_desc_7_wuser_6_reg_we),
                              .uc2rb_desc_7_wuser_7_reg_we(uc2rb_desc_7_wuser_7_reg_we),
                              .uc2rb_desc_7_wuser_8_reg_we(uc2rb_desc_7_wuser_8_reg_we),
                              .uc2rb_desc_7_wuser_9_reg_we(uc2rb_desc_7_wuser_9_reg_we),
                              .uc2rb_desc_7_wuser_10_reg_we(uc2rb_desc_7_wuser_10_reg_we),
                              .uc2rb_desc_7_wuser_11_reg_we(uc2rb_desc_7_wuser_11_reg_we),
                              .uc2rb_desc_7_wuser_12_reg_we(uc2rb_desc_7_wuser_12_reg_we),
                              .uc2rb_desc_7_wuser_13_reg_we(uc2rb_desc_7_wuser_13_reg_we),
                              .uc2rb_desc_7_wuser_14_reg_we(uc2rb_desc_7_wuser_14_reg_we),
                              .uc2rb_desc_7_wuser_15_reg_we(uc2rb_desc_7_wuser_15_reg_we),
                              .uc2rb_desc_8_txn_type_reg_we(uc2rb_desc_8_txn_type_reg_we),
                              .uc2rb_desc_8_size_reg_we(uc2rb_desc_8_size_reg_we),
                              .uc2rb_desc_8_data_offset_reg_we(uc2rb_desc_8_data_offset_reg_we),
                              .uc2rb_desc_8_axsize_reg_we(uc2rb_desc_8_axsize_reg_we),
                              .uc2rb_desc_8_attr_reg_we(uc2rb_desc_8_attr_reg_we),
                              .uc2rb_desc_8_axaddr_0_reg_we(uc2rb_desc_8_axaddr_0_reg_we),
                              .uc2rb_desc_8_axaddr_1_reg_we(uc2rb_desc_8_axaddr_1_reg_we),
                              .uc2rb_desc_8_axaddr_2_reg_we(uc2rb_desc_8_axaddr_2_reg_we),
                              .uc2rb_desc_8_axaddr_3_reg_we(uc2rb_desc_8_axaddr_3_reg_we),
                              .uc2rb_desc_8_axid_0_reg_we(uc2rb_desc_8_axid_0_reg_we),
                              .uc2rb_desc_8_axid_1_reg_we(uc2rb_desc_8_axid_1_reg_we),
                              .uc2rb_desc_8_axid_2_reg_we(uc2rb_desc_8_axid_2_reg_we),
                              .uc2rb_desc_8_axid_3_reg_we(uc2rb_desc_8_axid_3_reg_we),
                              .uc2rb_desc_8_axuser_0_reg_we(uc2rb_desc_8_axuser_0_reg_we),
                              .uc2rb_desc_8_axuser_1_reg_we(uc2rb_desc_8_axuser_1_reg_we),
                              .uc2rb_desc_8_axuser_2_reg_we(uc2rb_desc_8_axuser_2_reg_we),
                              .uc2rb_desc_8_axuser_3_reg_we(uc2rb_desc_8_axuser_3_reg_we),
                              .uc2rb_desc_8_axuser_4_reg_we(uc2rb_desc_8_axuser_4_reg_we),
                              .uc2rb_desc_8_axuser_5_reg_we(uc2rb_desc_8_axuser_5_reg_we),
                              .uc2rb_desc_8_axuser_6_reg_we(uc2rb_desc_8_axuser_6_reg_we),
                              .uc2rb_desc_8_axuser_7_reg_we(uc2rb_desc_8_axuser_7_reg_we),
                              .uc2rb_desc_8_axuser_8_reg_we(uc2rb_desc_8_axuser_8_reg_we),
                              .uc2rb_desc_8_axuser_9_reg_we(uc2rb_desc_8_axuser_9_reg_we),
                              .uc2rb_desc_8_axuser_10_reg_we(uc2rb_desc_8_axuser_10_reg_we),
                              .uc2rb_desc_8_axuser_11_reg_we(uc2rb_desc_8_axuser_11_reg_we),
                              .uc2rb_desc_8_axuser_12_reg_we(uc2rb_desc_8_axuser_12_reg_we),
                              .uc2rb_desc_8_axuser_13_reg_we(uc2rb_desc_8_axuser_13_reg_we),
                              .uc2rb_desc_8_axuser_14_reg_we(uc2rb_desc_8_axuser_14_reg_we),
                              .uc2rb_desc_8_axuser_15_reg_we(uc2rb_desc_8_axuser_15_reg_we),
                              .uc2rb_desc_8_wuser_0_reg_we(uc2rb_desc_8_wuser_0_reg_we),
                              .uc2rb_desc_8_wuser_1_reg_we(uc2rb_desc_8_wuser_1_reg_we),
                              .uc2rb_desc_8_wuser_2_reg_we(uc2rb_desc_8_wuser_2_reg_we),
                              .uc2rb_desc_8_wuser_3_reg_we(uc2rb_desc_8_wuser_3_reg_we),
                              .uc2rb_desc_8_wuser_4_reg_we(uc2rb_desc_8_wuser_4_reg_we),
                              .uc2rb_desc_8_wuser_5_reg_we(uc2rb_desc_8_wuser_5_reg_we),
                              .uc2rb_desc_8_wuser_6_reg_we(uc2rb_desc_8_wuser_6_reg_we),
                              .uc2rb_desc_8_wuser_7_reg_we(uc2rb_desc_8_wuser_7_reg_we),
                              .uc2rb_desc_8_wuser_8_reg_we(uc2rb_desc_8_wuser_8_reg_we),
                              .uc2rb_desc_8_wuser_9_reg_we(uc2rb_desc_8_wuser_9_reg_we),
                              .uc2rb_desc_8_wuser_10_reg_we(uc2rb_desc_8_wuser_10_reg_we),
                              .uc2rb_desc_8_wuser_11_reg_we(uc2rb_desc_8_wuser_11_reg_we),
                              .uc2rb_desc_8_wuser_12_reg_we(uc2rb_desc_8_wuser_12_reg_we),
                              .uc2rb_desc_8_wuser_13_reg_we(uc2rb_desc_8_wuser_13_reg_we),
                              .uc2rb_desc_8_wuser_14_reg_we(uc2rb_desc_8_wuser_14_reg_we),
                              .uc2rb_desc_8_wuser_15_reg_we(uc2rb_desc_8_wuser_15_reg_we),
                              .uc2rb_desc_9_txn_type_reg_we(uc2rb_desc_9_txn_type_reg_we),
                              .uc2rb_desc_9_size_reg_we(uc2rb_desc_9_size_reg_we),
                              .uc2rb_desc_9_data_offset_reg_we(uc2rb_desc_9_data_offset_reg_we),
                              .uc2rb_desc_9_axsize_reg_we(uc2rb_desc_9_axsize_reg_we),
                              .uc2rb_desc_9_attr_reg_we(uc2rb_desc_9_attr_reg_we),
                              .uc2rb_desc_9_axaddr_0_reg_we(uc2rb_desc_9_axaddr_0_reg_we),
                              .uc2rb_desc_9_axaddr_1_reg_we(uc2rb_desc_9_axaddr_1_reg_we),
                              .uc2rb_desc_9_axaddr_2_reg_we(uc2rb_desc_9_axaddr_2_reg_we),
                              .uc2rb_desc_9_axaddr_3_reg_we(uc2rb_desc_9_axaddr_3_reg_we),
                              .uc2rb_desc_9_axid_0_reg_we(uc2rb_desc_9_axid_0_reg_we),
                              .uc2rb_desc_9_axid_1_reg_we(uc2rb_desc_9_axid_1_reg_we),
                              .uc2rb_desc_9_axid_2_reg_we(uc2rb_desc_9_axid_2_reg_we),
                              .uc2rb_desc_9_axid_3_reg_we(uc2rb_desc_9_axid_3_reg_we),
                              .uc2rb_desc_9_axuser_0_reg_we(uc2rb_desc_9_axuser_0_reg_we),
                              .uc2rb_desc_9_axuser_1_reg_we(uc2rb_desc_9_axuser_1_reg_we),
                              .uc2rb_desc_9_axuser_2_reg_we(uc2rb_desc_9_axuser_2_reg_we),
                              .uc2rb_desc_9_axuser_3_reg_we(uc2rb_desc_9_axuser_3_reg_we),
                              .uc2rb_desc_9_axuser_4_reg_we(uc2rb_desc_9_axuser_4_reg_we),
                              .uc2rb_desc_9_axuser_5_reg_we(uc2rb_desc_9_axuser_5_reg_we),
                              .uc2rb_desc_9_axuser_6_reg_we(uc2rb_desc_9_axuser_6_reg_we),
                              .uc2rb_desc_9_axuser_7_reg_we(uc2rb_desc_9_axuser_7_reg_we),
                              .uc2rb_desc_9_axuser_8_reg_we(uc2rb_desc_9_axuser_8_reg_we),
                              .uc2rb_desc_9_axuser_9_reg_we(uc2rb_desc_9_axuser_9_reg_we),
                              .uc2rb_desc_9_axuser_10_reg_we(uc2rb_desc_9_axuser_10_reg_we),
                              .uc2rb_desc_9_axuser_11_reg_we(uc2rb_desc_9_axuser_11_reg_we),
                              .uc2rb_desc_9_axuser_12_reg_we(uc2rb_desc_9_axuser_12_reg_we),
                              .uc2rb_desc_9_axuser_13_reg_we(uc2rb_desc_9_axuser_13_reg_we),
                              .uc2rb_desc_9_axuser_14_reg_we(uc2rb_desc_9_axuser_14_reg_we),
                              .uc2rb_desc_9_axuser_15_reg_we(uc2rb_desc_9_axuser_15_reg_we),
                              .uc2rb_desc_9_wuser_0_reg_we(uc2rb_desc_9_wuser_0_reg_we),
                              .uc2rb_desc_9_wuser_1_reg_we(uc2rb_desc_9_wuser_1_reg_we),
                              .uc2rb_desc_9_wuser_2_reg_we(uc2rb_desc_9_wuser_2_reg_we),
                              .uc2rb_desc_9_wuser_3_reg_we(uc2rb_desc_9_wuser_3_reg_we),
                              .uc2rb_desc_9_wuser_4_reg_we(uc2rb_desc_9_wuser_4_reg_we),
                              .uc2rb_desc_9_wuser_5_reg_we(uc2rb_desc_9_wuser_5_reg_we),
                              .uc2rb_desc_9_wuser_6_reg_we(uc2rb_desc_9_wuser_6_reg_we),
                              .uc2rb_desc_9_wuser_7_reg_we(uc2rb_desc_9_wuser_7_reg_we),
                              .uc2rb_desc_9_wuser_8_reg_we(uc2rb_desc_9_wuser_8_reg_we),
                              .uc2rb_desc_9_wuser_9_reg_we(uc2rb_desc_9_wuser_9_reg_we),
                              .uc2rb_desc_9_wuser_10_reg_we(uc2rb_desc_9_wuser_10_reg_we),
                              .uc2rb_desc_9_wuser_11_reg_we(uc2rb_desc_9_wuser_11_reg_we),
                              .uc2rb_desc_9_wuser_12_reg_we(uc2rb_desc_9_wuser_12_reg_we),
                              .uc2rb_desc_9_wuser_13_reg_we(uc2rb_desc_9_wuser_13_reg_we),
                              .uc2rb_desc_9_wuser_14_reg_we(uc2rb_desc_9_wuser_14_reg_we),
                              .uc2rb_desc_9_wuser_15_reg_we(uc2rb_desc_9_wuser_15_reg_we),
                              .uc2rb_desc_10_txn_type_reg_we(uc2rb_desc_10_txn_type_reg_we),
                              .uc2rb_desc_10_size_reg_we(uc2rb_desc_10_size_reg_we),
                              .uc2rb_desc_10_data_offset_reg_we(uc2rb_desc_10_data_offset_reg_we),
                              .uc2rb_desc_10_axsize_reg_we(uc2rb_desc_10_axsize_reg_we),
                              .uc2rb_desc_10_attr_reg_we(uc2rb_desc_10_attr_reg_we),
                              .uc2rb_desc_10_axaddr_0_reg_we(uc2rb_desc_10_axaddr_0_reg_we),
                              .uc2rb_desc_10_axaddr_1_reg_we(uc2rb_desc_10_axaddr_1_reg_we),
                              .uc2rb_desc_10_axaddr_2_reg_we(uc2rb_desc_10_axaddr_2_reg_we),
                              .uc2rb_desc_10_axaddr_3_reg_we(uc2rb_desc_10_axaddr_3_reg_we),
                              .uc2rb_desc_10_axid_0_reg_we(uc2rb_desc_10_axid_0_reg_we),
                              .uc2rb_desc_10_axid_1_reg_we(uc2rb_desc_10_axid_1_reg_we),
                              .uc2rb_desc_10_axid_2_reg_we(uc2rb_desc_10_axid_2_reg_we),
                              .uc2rb_desc_10_axid_3_reg_we(uc2rb_desc_10_axid_3_reg_we),
                              .uc2rb_desc_10_axuser_0_reg_we(uc2rb_desc_10_axuser_0_reg_we),
                              .uc2rb_desc_10_axuser_1_reg_we(uc2rb_desc_10_axuser_1_reg_we),
                              .uc2rb_desc_10_axuser_2_reg_we(uc2rb_desc_10_axuser_2_reg_we),
                              .uc2rb_desc_10_axuser_3_reg_we(uc2rb_desc_10_axuser_3_reg_we),
                              .uc2rb_desc_10_axuser_4_reg_we(uc2rb_desc_10_axuser_4_reg_we),
                              .uc2rb_desc_10_axuser_5_reg_we(uc2rb_desc_10_axuser_5_reg_we),
                              .uc2rb_desc_10_axuser_6_reg_we(uc2rb_desc_10_axuser_6_reg_we),
                              .uc2rb_desc_10_axuser_7_reg_we(uc2rb_desc_10_axuser_7_reg_we),
                              .uc2rb_desc_10_axuser_8_reg_we(uc2rb_desc_10_axuser_8_reg_we),
                              .uc2rb_desc_10_axuser_9_reg_we(uc2rb_desc_10_axuser_9_reg_we),
                              .uc2rb_desc_10_axuser_10_reg_we(uc2rb_desc_10_axuser_10_reg_we),
                              .uc2rb_desc_10_axuser_11_reg_we(uc2rb_desc_10_axuser_11_reg_we),
                              .uc2rb_desc_10_axuser_12_reg_we(uc2rb_desc_10_axuser_12_reg_we),
                              .uc2rb_desc_10_axuser_13_reg_we(uc2rb_desc_10_axuser_13_reg_we),
                              .uc2rb_desc_10_axuser_14_reg_we(uc2rb_desc_10_axuser_14_reg_we),
                              .uc2rb_desc_10_axuser_15_reg_we(uc2rb_desc_10_axuser_15_reg_we),
                              .uc2rb_desc_10_wuser_0_reg_we(uc2rb_desc_10_wuser_0_reg_we),
                              .uc2rb_desc_10_wuser_1_reg_we(uc2rb_desc_10_wuser_1_reg_we),
                              .uc2rb_desc_10_wuser_2_reg_we(uc2rb_desc_10_wuser_2_reg_we),
                              .uc2rb_desc_10_wuser_3_reg_we(uc2rb_desc_10_wuser_3_reg_we),
                              .uc2rb_desc_10_wuser_4_reg_we(uc2rb_desc_10_wuser_4_reg_we),
                              .uc2rb_desc_10_wuser_5_reg_we(uc2rb_desc_10_wuser_5_reg_we),
                              .uc2rb_desc_10_wuser_6_reg_we(uc2rb_desc_10_wuser_6_reg_we),
                              .uc2rb_desc_10_wuser_7_reg_we(uc2rb_desc_10_wuser_7_reg_we),
                              .uc2rb_desc_10_wuser_8_reg_we(uc2rb_desc_10_wuser_8_reg_we),
                              .uc2rb_desc_10_wuser_9_reg_we(uc2rb_desc_10_wuser_9_reg_we),
                              .uc2rb_desc_10_wuser_10_reg_we(uc2rb_desc_10_wuser_10_reg_we),
                              .uc2rb_desc_10_wuser_11_reg_we(uc2rb_desc_10_wuser_11_reg_we),
                              .uc2rb_desc_10_wuser_12_reg_we(uc2rb_desc_10_wuser_12_reg_we),
                              .uc2rb_desc_10_wuser_13_reg_we(uc2rb_desc_10_wuser_13_reg_we),
                              .uc2rb_desc_10_wuser_14_reg_we(uc2rb_desc_10_wuser_14_reg_we),
                              .uc2rb_desc_10_wuser_15_reg_we(uc2rb_desc_10_wuser_15_reg_we),
                              .uc2rb_desc_11_txn_type_reg_we(uc2rb_desc_11_txn_type_reg_we),
                              .uc2rb_desc_11_size_reg_we(uc2rb_desc_11_size_reg_we),
                              .uc2rb_desc_11_data_offset_reg_we(uc2rb_desc_11_data_offset_reg_we),
                              .uc2rb_desc_11_axsize_reg_we(uc2rb_desc_11_axsize_reg_we),
                              .uc2rb_desc_11_attr_reg_we(uc2rb_desc_11_attr_reg_we),
                              .uc2rb_desc_11_axaddr_0_reg_we(uc2rb_desc_11_axaddr_0_reg_we),
                              .uc2rb_desc_11_axaddr_1_reg_we(uc2rb_desc_11_axaddr_1_reg_we),
                              .uc2rb_desc_11_axaddr_2_reg_we(uc2rb_desc_11_axaddr_2_reg_we),
                              .uc2rb_desc_11_axaddr_3_reg_we(uc2rb_desc_11_axaddr_3_reg_we),
                              .uc2rb_desc_11_axid_0_reg_we(uc2rb_desc_11_axid_0_reg_we),
                              .uc2rb_desc_11_axid_1_reg_we(uc2rb_desc_11_axid_1_reg_we),
                              .uc2rb_desc_11_axid_2_reg_we(uc2rb_desc_11_axid_2_reg_we),
                              .uc2rb_desc_11_axid_3_reg_we(uc2rb_desc_11_axid_3_reg_we),
                              .uc2rb_desc_11_axuser_0_reg_we(uc2rb_desc_11_axuser_0_reg_we),
                              .uc2rb_desc_11_axuser_1_reg_we(uc2rb_desc_11_axuser_1_reg_we),
                              .uc2rb_desc_11_axuser_2_reg_we(uc2rb_desc_11_axuser_2_reg_we),
                              .uc2rb_desc_11_axuser_3_reg_we(uc2rb_desc_11_axuser_3_reg_we),
                              .uc2rb_desc_11_axuser_4_reg_we(uc2rb_desc_11_axuser_4_reg_we),
                              .uc2rb_desc_11_axuser_5_reg_we(uc2rb_desc_11_axuser_5_reg_we),
                              .uc2rb_desc_11_axuser_6_reg_we(uc2rb_desc_11_axuser_6_reg_we),
                              .uc2rb_desc_11_axuser_7_reg_we(uc2rb_desc_11_axuser_7_reg_we),
                              .uc2rb_desc_11_axuser_8_reg_we(uc2rb_desc_11_axuser_8_reg_we),
                              .uc2rb_desc_11_axuser_9_reg_we(uc2rb_desc_11_axuser_9_reg_we),
                              .uc2rb_desc_11_axuser_10_reg_we(uc2rb_desc_11_axuser_10_reg_we),
                              .uc2rb_desc_11_axuser_11_reg_we(uc2rb_desc_11_axuser_11_reg_we),
                              .uc2rb_desc_11_axuser_12_reg_we(uc2rb_desc_11_axuser_12_reg_we),
                              .uc2rb_desc_11_axuser_13_reg_we(uc2rb_desc_11_axuser_13_reg_we),
                              .uc2rb_desc_11_axuser_14_reg_we(uc2rb_desc_11_axuser_14_reg_we),
                              .uc2rb_desc_11_axuser_15_reg_we(uc2rb_desc_11_axuser_15_reg_we),
                              .uc2rb_desc_11_wuser_0_reg_we(uc2rb_desc_11_wuser_0_reg_we),
                              .uc2rb_desc_11_wuser_1_reg_we(uc2rb_desc_11_wuser_1_reg_we),
                              .uc2rb_desc_11_wuser_2_reg_we(uc2rb_desc_11_wuser_2_reg_we),
                              .uc2rb_desc_11_wuser_3_reg_we(uc2rb_desc_11_wuser_3_reg_we),
                              .uc2rb_desc_11_wuser_4_reg_we(uc2rb_desc_11_wuser_4_reg_we),
                              .uc2rb_desc_11_wuser_5_reg_we(uc2rb_desc_11_wuser_5_reg_we),
                              .uc2rb_desc_11_wuser_6_reg_we(uc2rb_desc_11_wuser_6_reg_we),
                              .uc2rb_desc_11_wuser_7_reg_we(uc2rb_desc_11_wuser_7_reg_we),
                              .uc2rb_desc_11_wuser_8_reg_we(uc2rb_desc_11_wuser_8_reg_we),
                              .uc2rb_desc_11_wuser_9_reg_we(uc2rb_desc_11_wuser_9_reg_we),
                              .uc2rb_desc_11_wuser_10_reg_we(uc2rb_desc_11_wuser_10_reg_we),
                              .uc2rb_desc_11_wuser_11_reg_we(uc2rb_desc_11_wuser_11_reg_we),
                              .uc2rb_desc_11_wuser_12_reg_we(uc2rb_desc_11_wuser_12_reg_we),
                              .uc2rb_desc_11_wuser_13_reg_we(uc2rb_desc_11_wuser_13_reg_we),
                              .uc2rb_desc_11_wuser_14_reg_we(uc2rb_desc_11_wuser_14_reg_we),
                              .uc2rb_desc_11_wuser_15_reg_we(uc2rb_desc_11_wuser_15_reg_we),
                              .uc2rb_desc_12_txn_type_reg_we(uc2rb_desc_12_txn_type_reg_we),
                              .uc2rb_desc_12_size_reg_we(uc2rb_desc_12_size_reg_we),
                              .uc2rb_desc_12_data_offset_reg_we(uc2rb_desc_12_data_offset_reg_we),
                              .uc2rb_desc_12_axsize_reg_we(uc2rb_desc_12_axsize_reg_we),
                              .uc2rb_desc_12_attr_reg_we(uc2rb_desc_12_attr_reg_we),
                              .uc2rb_desc_12_axaddr_0_reg_we(uc2rb_desc_12_axaddr_0_reg_we),
                              .uc2rb_desc_12_axaddr_1_reg_we(uc2rb_desc_12_axaddr_1_reg_we),
                              .uc2rb_desc_12_axaddr_2_reg_we(uc2rb_desc_12_axaddr_2_reg_we),
                              .uc2rb_desc_12_axaddr_3_reg_we(uc2rb_desc_12_axaddr_3_reg_we),
                              .uc2rb_desc_12_axid_0_reg_we(uc2rb_desc_12_axid_0_reg_we),
                              .uc2rb_desc_12_axid_1_reg_we(uc2rb_desc_12_axid_1_reg_we),
                              .uc2rb_desc_12_axid_2_reg_we(uc2rb_desc_12_axid_2_reg_we),
                              .uc2rb_desc_12_axid_3_reg_we(uc2rb_desc_12_axid_3_reg_we),
                              .uc2rb_desc_12_axuser_0_reg_we(uc2rb_desc_12_axuser_0_reg_we),
                              .uc2rb_desc_12_axuser_1_reg_we(uc2rb_desc_12_axuser_1_reg_we),
                              .uc2rb_desc_12_axuser_2_reg_we(uc2rb_desc_12_axuser_2_reg_we),
                              .uc2rb_desc_12_axuser_3_reg_we(uc2rb_desc_12_axuser_3_reg_we),
                              .uc2rb_desc_12_axuser_4_reg_we(uc2rb_desc_12_axuser_4_reg_we),
                              .uc2rb_desc_12_axuser_5_reg_we(uc2rb_desc_12_axuser_5_reg_we),
                              .uc2rb_desc_12_axuser_6_reg_we(uc2rb_desc_12_axuser_6_reg_we),
                              .uc2rb_desc_12_axuser_7_reg_we(uc2rb_desc_12_axuser_7_reg_we),
                              .uc2rb_desc_12_axuser_8_reg_we(uc2rb_desc_12_axuser_8_reg_we),
                              .uc2rb_desc_12_axuser_9_reg_we(uc2rb_desc_12_axuser_9_reg_we),
                              .uc2rb_desc_12_axuser_10_reg_we(uc2rb_desc_12_axuser_10_reg_we),
                              .uc2rb_desc_12_axuser_11_reg_we(uc2rb_desc_12_axuser_11_reg_we),
                              .uc2rb_desc_12_axuser_12_reg_we(uc2rb_desc_12_axuser_12_reg_we),
                              .uc2rb_desc_12_axuser_13_reg_we(uc2rb_desc_12_axuser_13_reg_we),
                              .uc2rb_desc_12_axuser_14_reg_we(uc2rb_desc_12_axuser_14_reg_we),
                              .uc2rb_desc_12_axuser_15_reg_we(uc2rb_desc_12_axuser_15_reg_we),
                              .uc2rb_desc_12_wuser_0_reg_we(uc2rb_desc_12_wuser_0_reg_we),
                              .uc2rb_desc_12_wuser_1_reg_we(uc2rb_desc_12_wuser_1_reg_we),
                              .uc2rb_desc_12_wuser_2_reg_we(uc2rb_desc_12_wuser_2_reg_we),
                              .uc2rb_desc_12_wuser_3_reg_we(uc2rb_desc_12_wuser_3_reg_we),
                              .uc2rb_desc_12_wuser_4_reg_we(uc2rb_desc_12_wuser_4_reg_we),
                              .uc2rb_desc_12_wuser_5_reg_we(uc2rb_desc_12_wuser_5_reg_we),
                              .uc2rb_desc_12_wuser_6_reg_we(uc2rb_desc_12_wuser_6_reg_we),
                              .uc2rb_desc_12_wuser_7_reg_we(uc2rb_desc_12_wuser_7_reg_we),
                              .uc2rb_desc_12_wuser_8_reg_we(uc2rb_desc_12_wuser_8_reg_we),
                              .uc2rb_desc_12_wuser_9_reg_we(uc2rb_desc_12_wuser_9_reg_we),
                              .uc2rb_desc_12_wuser_10_reg_we(uc2rb_desc_12_wuser_10_reg_we),
                              .uc2rb_desc_12_wuser_11_reg_we(uc2rb_desc_12_wuser_11_reg_we),
                              .uc2rb_desc_12_wuser_12_reg_we(uc2rb_desc_12_wuser_12_reg_we),
                              .uc2rb_desc_12_wuser_13_reg_we(uc2rb_desc_12_wuser_13_reg_we),
                              .uc2rb_desc_12_wuser_14_reg_we(uc2rb_desc_12_wuser_14_reg_we),
                              .uc2rb_desc_12_wuser_15_reg_we(uc2rb_desc_12_wuser_15_reg_we),
                              .uc2rb_desc_13_txn_type_reg_we(uc2rb_desc_13_txn_type_reg_we),
                              .uc2rb_desc_13_size_reg_we(uc2rb_desc_13_size_reg_we),
                              .uc2rb_desc_13_data_offset_reg_we(uc2rb_desc_13_data_offset_reg_we),
                              .uc2rb_desc_13_axsize_reg_we(uc2rb_desc_13_axsize_reg_we),
                              .uc2rb_desc_13_attr_reg_we(uc2rb_desc_13_attr_reg_we),
                              .uc2rb_desc_13_axaddr_0_reg_we(uc2rb_desc_13_axaddr_0_reg_we),
                              .uc2rb_desc_13_axaddr_1_reg_we(uc2rb_desc_13_axaddr_1_reg_we),
                              .uc2rb_desc_13_axaddr_2_reg_we(uc2rb_desc_13_axaddr_2_reg_we),
                              .uc2rb_desc_13_axaddr_3_reg_we(uc2rb_desc_13_axaddr_3_reg_we),
                              .uc2rb_desc_13_axid_0_reg_we(uc2rb_desc_13_axid_0_reg_we),
                              .uc2rb_desc_13_axid_1_reg_we(uc2rb_desc_13_axid_1_reg_we),
                              .uc2rb_desc_13_axid_2_reg_we(uc2rb_desc_13_axid_2_reg_we),
                              .uc2rb_desc_13_axid_3_reg_we(uc2rb_desc_13_axid_3_reg_we),
                              .uc2rb_desc_13_axuser_0_reg_we(uc2rb_desc_13_axuser_0_reg_we),
                              .uc2rb_desc_13_axuser_1_reg_we(uc2rb_desc_13_axuser_1_reg_we),
                              .uc2rb_desc_13_axuser_2_reg_we(uc2rb_desc_13_axuser_2_reg_we),
                              .uc2rb_desc_13_axuser_3_reg_we(uc2rb_desc_13_axuser_3_reg_we),
                              .uc2rb_desc_13_axuser_4_reg_we(uc2rb_desc_13_axuser_4_reg_we),
                              .uc2rb_desc_13_axuser_5_reg_we(uc2rb_desc_13_axuser_5_reg_we),
                              .uc2rb_desc_13_axuser_6_reg_we(uc2rb_desc_13_axuser_6_reg_we),
                              .uc2rb_desc_13_axuser_7_reg_we(uc2rb_desc_13_axuser_7_reg_we),
                              .uc2rb_desc_13_axuser_8_reg_we(uc2rb_desc_13_axuser_8_reg_we),
                              .uc2rb_desc_13_axuser_9_reg_we(uc2rb_desc_13_axuser_9_reg_we),
                              .uc2rb_desc_13_axuser_10_reg_we(uc2rb_desc_13_axuser_10_reg_we),
                              .uc2rb_desc_13_axuser_11_reg_we(uc2rb_desc_13_axuser_11_reg_we),
                              .uc2rb_desc_13_axuser_12_reg_we(uc2rb_desc_13_axuser_12_reg_we),
                              .uc2rb_desc_13_axuser_13_reg_we(uc2rb_desc_13_axuser_13_reg_we),
                              .uc2rb_desc_13_axuser_14_reg_we(uc2rb_desc_13_axuser_14_reg_we),
                              .uc2rb_desc_13_axuser_15_reg_we(uc2rb_desc_13_axuser_15_reg_we),
                              .uc2rb_desc_13_wuser_0_reg_we(uc2rb_desc_13_wuser_0_reg_we),
                              .uc2rb_desc_13_wuser_1_reg_we(uc2rb_desc_13_wuser_1_reg_we),
                              .uc2rb_desc_13_wuser_2_reg_we(uc2rb_desc_13_wuser_2_reg_we),
                              .uc2rb_desc_13_wuser_3_reg_we(uc2rb_desc_13_wuser_3_reg_we),
                              .uc2rb_desc_13_wuser_4_reg_we(uc2rb_desc_13_wuser_4_reg_we),
                              .uc2rb_desc_13_wuser_5_reg_we(uc2rb_desc_13_wuser_5_reg_we),
                              .uc2rb_desc_13_wuser_6_reg_we(uc2rb_desc_13_wuser_6_reg_we),
                              .uc2rb_desc_13_wuser_7_reg_we(uc2rb_desc_13_wuser_7_reg_we),
                              .uc2rb_desc_13_wuser_8_reg_we(uc2rb_desc_13_wuser_8_reg_we),
                              .uc2rb_desc_13_wuser_9_reg_we(uc2rb_desc_13_wuser_9_reg_we),
                              .uc2rb_desc_13_wuser_10_reg_we(uc2rb_desc_13_wuser_10_reg_we),
                              .uc2rb_desc_13_wuser_11_reg_we(uc2rb_desc_13_wuser_11_reg_we),
                              .uc2rb_desc_13_wuser_12_reg_we(uc2rb_desc_13_wuser_12_reg_we),
                              .uc2rb_desc_13_wuser_13_reg_we(uc2rb_desc_13_wuser_13_reg_we),
                              .uc2rb_desc_13_wuser_14_reg_we(uc2rb_desc_13_wuser_14_reg_we),
                              .uc2rb_desc_13_wuser_15_reg_we(uc2rb_desc_13_wuser_15_reg_we),
                              .uc2rb_desc_14_txn_type_reg_we(uc2rb_desc_14_txn_type_reg_we),
                              .uc2rb_desc_14_size_reg_we(uc2rb_desc_14_size_reg_we),
                              .uc2rb_desc_14_data_offset_reg_we(uc2rb_desc_14_data_offset_reg_we),
                              .uc2rb_desc_14_axsize_reg_we(uc2rb_desc_14_axsize_reg_we),
                              .uc2rb_desc_14_attr_reg_we(uc2rb_desc_14_attr_reg_we),
                              .uc2rb_desc_14_axaddr_0_reg_we(uc2rb_desc_14_axaddr_0_reg_we),
                              .uc2rb_desc_14_axaddr_1_reg_we(uc2rb_desc_14_axaddr_1_reg_we),
                              .uc2rb_desc_14_axaddr_2_reg_we(uc2rb_desc_14_axaddr_2_reg_we),
                              .uc2rb_desc_14_axaddr_3_reg_we(uc2rb_desc_14_axaddr_3_reg_we),
                              .uc2rb_desc_14_axid_0_reg_we(uc2rb_desc_14_axid_0_reg_we),
                              .uc2rb_desc_14_axid_1_reg_we(uc2rb_desc_14_axid_1_reg_we),
                              .uc2rb_desc_14_axid_2_reg_we(uc2rb_desc_14_axid_2_reg_we),
                              .uc2rb_desc_14_axid_3_reg_we(uc2rb_desc_14_axid_3_reg_we),
                              .uc2rb_desc_14_axuser_0_reg_we(uc2rb_desc_14_axuser_0_reg_we),
                              .uc2rb_desc_14_axuser_1_reg_we(uc2rb_desc_14_axuser_1_reg_we),
                              .uc2rb_desc_14_axuser_2_reg_we(uc2rb_desc_14_axuser_2_reg_we),
                              .uc2rb_desc_14_axuser_3_reg_we(uc2rb_desc_14_axuser_3_reg_we),
                              .uc2rb_desc_14_axuser_4_reg_we(uc2rb_desc_14_axuser_4_reg_we),
                              .uc2rb_desc_14_axuser_5_reg_we(uc2rb_desc_14_axuser_5_reg_we),
                              .uc2rb_desc_14_axuser_6_reg_we(uc2rb_desc_14_axuser_6_reg_we),
                              .uc2rb_desc_14_axuser_7_reg_we(uc2rb_desc_14_axuser_7_reg_we),
                              .uc2rb_desc_14_axuser_8_reg_we(uc2rb_desc_14_axuser_8_reg_we),
                              .uc2rb_desc_14_axuser_9_reg_we(uc2rb_desc_14_axuser_9_reg_we),
                              .uc2rb_desc_14_axuser_10_reg_we(uc2rb_desc_14_axuser_10_reg_we),
                              .uc2rb_desc_14_axuser_11_reg_we(uc2rb_desc_14_axuser_11_reg_we),
                              .uc2rb_desc_14_axuser_12_reg_we(uc2rb_desc_14_axuser_12_reg_we),
                              .uc2rb_desc_14_axuser_13_reg_we(uc2rb_desc_14_axuser_13_reg_we),
                              .uc2rb_desc_14_axuser_14_reg_we(uc2rb_desc_14_axuser_14_reg_we),
                              .uc2rb_desc_14_axuser_15_reg_we(uc2rb_desc_14_axuser_15_reg_we),
                              .uc2rb_desc_14_wuser_0_reg_we(uc2rb_desc_14_wuser_0_reg_we),
                              .uc2rb_desc_14_wuser_1_reg_we(uc2rb_desc_14_wuser_1_reg_we),
                              .uc2rb_desc_14_wuser_2_reg_we(uc2rb_desc_14_wuser_2_reg_we),
                              .uc2rb_desc_14_wuser_3_reg_we(uc2rb_desc_14_wuser_3_reg_we),
                              .uc2rb_desc_14_wuser_4_reg_we(uc2rb_desc_14_wuser_4_reg_we),
                              .uc2rb_desc_14_wuser_5_reg_we(uc2rb_desc_14_wuser_5_reg_we),
                              .uc2rb_desc_14_wuser_6_reg_we(uc2rb_desc_14_wuser_6_reg_we),
                              .uc2rb_desc_14_wuser_7_reg_we(uc2rb_desc_14_wuser_7_reg_we),
                              .uc2rb_desc_14_wuser_8_reg_we(uc2rb_desc_14_wuser_8_reg_we),
                              .uc2rb_desc_14_wuser_9_reg_we(uc2rb_desc_14_wuser_9_reg_we),
                              .uc2rb_desc_14_wuser_10_reg_we(uc2rb_desc_14_wuser_10_reg_we),
                              .uc2rb_desc_14_wuser_11_reg_we(uc2rb_desc_14_wuser_11_reg_we),
                              .uc2rb_desc_14_wuser_12_reg_we(uc2rb_desc_14_wuser_12_reg_we),
                              .uc2rb_desc_14_wuser_13_reg_we(uc2rb_desc_14_wuser_13_reg_we),
                              .uc2rb_desc_14_wuser_14_reg_we(uc2rb_desc_14_wuser_14_reg_we),
                              .uc2rb_desc_14_wuser_15_reg_we(uc2rb_desc_14_wuser_15_reg_we),
                              .uc2rb_desc_15_txn_type_reg_we(uc2rb_desc_15_txn_type_reg_we),
                              .uc2rb_desc_15_size_reg_we(uc2rb_desc_15_size_reg_we),
                              .uc2rb_desc_15_data_offset_reg_we(uc2rb_desc_15_data_offset_reg_we),
                              .uc2rb_desc_15_axsize_reg_we(uc2rb_desc_15_axsize_reg_we),
                              .uc2rb_desc_15_attr_reg_we(uc2rb_desc_15_attr_reg_we),
                              .uc2rb_desc_15_axaddr_0_reg_we(uc2rb_desc_15_axaddr_0_reg_we),
                              .uc2rb_desc_15_axaddr_1_reg_we(uc2rb_desc_15_axaddr_1_reg_we),
                              .uc2rb_desc_15_axaddr_2_reg_we(uc2rb_desc_15_axaddr_2_reg_we),
                              .uc2rb_desc_15_axaddr_3_reg_we(uc2rb_desc_15_axaddr_3_reg_we),
                              .uc2rb_desc_15_axid_0_reg_we(uc2rb_desc_15_axid_0_reg_we),
                              .uc2rb_desc_15_axid_1_reg_we(uc2rb_desc_15_axid_1_reg_we),
                              .uc2rb_desc_15_axid_2_reg_we(uc2rb_desc_15_axid_2_reg_we),
                              .uc2rb_desc_15_axid_3_reg_we(uc2rb_desc_15_axid_3_reg_we),
                              .uc2rb_desc_15_axuser_0_reg_we(uc2rb_desc_15_axuser_0_reg_we),
                              .uc2rb_desc_15_axuser_1_reg_we(uc2rb_desc_15_axuser_1_reg_we),
                              .uc2rb_desc_15_axuser_2_reg_we(uc2rb_desc_15_axuser_2_reg_we),
                              .uc2rb_desc_15_axuser_3_reg_we(uc2rb_desc_15_axuser_3_reg_we),
                              .uc2rb_desc_15_axuser_4_reg_we(uc2rb_desc_15_axuser_4_reg_we),
                              .uc2rb_desc_15_axuser_5_reg_we(uc2rb_desc_15_axuser_5_reg_we),
                              .uc2rb_desc_15_axuser_6_reg_we(uc2rb_desc_15_axuser_6_reg_we),
                              .uc2rb_desc_15_axuser_7_reg_we(uc2rb_desc_15_axuser_7_reg_we),
                              .uc2rb_desc_15_axuser_8_reg_we(uc2rb_desc_15_axuser_8_reg_we),
                              .uc2rb_desc_15_axuser_9_reg_we(uc2rb_desc_15_axuser_9_reg_we),
                              .uc2rb_desc_15_axuser_10_reg_we(uc2rb_desc_15_axuser_10_reg_we),
                              .uc2rb_desc_15_axuser_11_reg_we(uc2rb_desc_15_axuser_11_reg_we),
                              .uc2rb_desc_15_axuser_12_reg_we(uc2rb_desc_15_axuser_12_reg_we),
                              .uc2rb_desc_15_axuser_13_reg_we(uc2rb_desc_15_axuser_13_reg_we),
                              .uc2rb_desc_15_axuser_14_reg_we(uc2rb_desc_15_axuser_14_reg_we),
                              .uc2rb_desc_15_axuser_15_reg_we(uc2rb_desc_15_axuser_15_reg_we),
                              .uc2rb_desc_15_wuser_0_reg_we(uc2rb_desc_15_wuser_0_reg_we),
                              .uc2rb_desc_15_wuser_1_reg_we(uc2rb_desc_15_wuser_1_reg_we),
                              .uc2rb_desc_15_wuser_2_reg_we(uc2rb_desc_15_wuser_2_reg_we),
                              .uc2rb_desc_15_wuser_3_reg_we(uc2rb_desc_15_wuser_3_reg_we),
                              .uc2rb_desc_15_wuser_4_reg_we(uc2rb_desc_15_wuser_4_reg_we),
                              .uc2rb_desc_15_wuser_5_reg_we(uc2rb_desc_15_wuser_5_reg_we),
                              .uc2rb_desc_15_wuser_6_reg_we(uc2rb_desc_15_wuser_6_reg_we),
                              .uc2rb_desc_15_wuser_7_reg_we(uc2rb_desc_15_wuser_7_reg_we),
                              .uc2rb_desc_15_wuser_8_reg_we(uc2rb_desc_15_wuser_8_reg_we),
                              .uc2rb_desc_15_wuser_9_reg_we(uc2rb_desc_15_wuser_9_reg_we),
                              .uc2rb_desc_15_wuser_10_reg_we(uc2rb_desc_15_wuser_10_reg_we),
                              .uc2rb_desc_15_wuser_11_reg_we(uc2rb_desc_15_wuser_11_reg_we),
                              .uc2rb_desc_15_wuser_12_reg_we(uc2rb_desc_15_wuser_12_reg_we),
                              .uc2rb_desc_15_wuser_13_reg_we(uc2rb_desc_15_wuser_13_reg_we),
                              .uc2rb_desc_15_wuser_14_reg_we(uc2rb_desc_15_wuser_14_reg_we),
                              .uc2rb_desc_15_wuser_15_reg_we(uc2rb_desc_15_wuser_15_reg_we),
   
							  .ih2rb_c2h_intr_status_0_reg     (ih2rb_c2h_intr_status_0_reg   ), 
							  .ih2rb_c2h_intr_status_1_reg     (ih2rb_c2h_intr_status_1_reg   ),
							  .ih2rb_intr_c2h_toggle_status_0_reg     (ih2rb_intr_c2h_toggle_status_0_reg   ), 
							  .ih2rb_intr_c2h_toggle_status_1_reg     (ih2rb_intr_c2h_toggle_status_1_reg   ), 
							  .ih2rb_c2h_gpio_0_reg     (ih2rb_c2h_gpio_0_reg   ),
							  .ih2rb_c2h_gpio_1_reg     (ih2rb_c2h_gpio_1_reg   ),
							  .ih2rb_c2h_gpio_2_reg     (ih2rb_c2h_gpio_2_reg   ),
							  .ih2rb_c2h_gpio_3_reg     (ih2rb_c2h_gpio_3_reg   ),
							  .ih2rb_c2h_gpio_4_reg     (ih2rb_c2h_gpio_4_reg   ),
							  .ih2rb_c2h_gpio_5_reg     (ih2rb_c2h_gpio_5_reg   ),
							  .ih2rb_c2h_gpio_6_reg     (ih2rb_c2h_gpio_6_reg   ),
							  .ih2rb_c2h_gpio_7_reg     (ih2rb_c2h_gpio_7_reg   ), 
							  .ih2rb_c2h_intr_status_0_reg_we  (ih2rb_c2h_intr_status_0_reg_we), 
							  .ih2rb_c2h_intr_status_1_reg_we  (ih2rb_c2h_intr_status_1_reg_we),
							  .ih2rb_intr_c2h_toggle_status_0_reg_we  (ih2rb_intr_c2h_toggle_status_0_reg_we), 
							  .ih2rb_intr_c2h_toggle_status_1_reg_we  (ih2rb_intr_c2h_toggle_status_1_reg_we), 
							  .ih2rb_c2h_gpio_0_reg_we  (ih2rb_c2h_gpio_0_reg_we),
							  .ih2rb_c2h_gpio_1_reg_we  (ih2rb_c2h_gpio_1_reg_we),
							  .ih2rb_c2h_gpio_2_reg_we  (ih2rb_c2h_gpio_2_reg_we),
							  .ih2rb_c2h_gpio_3_reg_we  (ih2rb_c2h_gpio_3_reg_we),
							  .ih2rb_c2h_gpio_4_reg_we  (ih2rb_c2h_gpio_4_reg_we),
							  .ih2rb_c2h_gpio_5_reg_we  (ih2rb_c2h_gpio_5_reg_we),
							  .ih2rb_c2h_gpio_6_reg_we  (ih2rb_c2h_gpio_6_reg_we),
							  .ih2rb_c2h_gpio_7_reg_we  (ih2rb_c2h_gpio_7_reg_we)
);
   host_master_s #(
                            .M_AXI_ADDR_WIDTH       (M_AXI_ADDR_WIDTH     ),  
                            .M_AXI_DATA_WIDTH       (M_AXI_DATA_WIDTH     ),  
                            .M_AXI_ID_WIDTH         (M_AXI_ID_WIDTH       ),  
                            .M_AXI_USER_WIDTH       (M_AXI_USER_WIDTH     ),  
                            .RAM_SIZE               (RAM_SIZE             ),  
                            .S_AXI_USR_DATA_WIDTH   (S_AXI_USR_DATA_WIDTH ),  
                            .MAX_DESC               (MAX_DESC             )  

     )

   host_control_slave_inst 
         (
          .axi_aclk                (axi_aclk),
          .axi_aresetn     (rst_n),
		  // Outputs
		  .hm2uc_done           (hm2uc_done),
		  .hm2rb_rd_addr        (hm2rb_rd_addr),
		  .hm2rb_wr_we          (hm2rb_wr_we),
		  .hm2rb_wr_bwe         (hm2rb_wr_bwe),
		  .hm2rb_wr_addr        (hm2rb_wr_addr),
		  .hm2rb_wr_data_in     (hm2rb_wr_data),
		  .hm2rb_wr_wstrb_in    (), //NC
		  .hm2rb_intr_error_status_reg_we(hm2rb_intr_error_status_reg_we),
          .hm2rb_intr_error_status_reg(hm2rb_intr_error_status_reg),
		  .rb2hm_intr_error_status_reg({31'h0,intr_error_status_reg[1]}),
		  .rb2hm_intr_error_clear_reg({31'h0,intr_error_clear_reg[1]}),

          // From RB-to HM
          
          .desc_0_txn_type_reg(desc_0_txn_type_reg),
          .desc_0_size_reg(desc_0_size_reg),
          .desc_0_data_offset_reg(desc_0_data_offset_reg),
          .desc_0_data_host_addr_0_reg(desc_0_data_host_addr_0_reg),
          .desc_0_data_host_addr_1_reg(desc_0_data_host_addr_1_reg),
          .desc_0_data_host_addr_2_reg(desc_0_data_host_addr_2_reg),
          .desc_0_data_host_addr_3_reg(desc_0_data_host_addr_3_reg),
          .desc_0_wstrb_host_addr_0_reg(desc_0_wstrb_host_addr_0_reg),
          .desc_0_wstrb_host_addr_1_reg(desc_0_wstrb_host_addr_1_reg),
          .desc_0_wstrb_host_addr_2_reg(desc_0_wstrb_host_addr_2_reg),
          .desc_0_wstrb_host_addr_3_reg(desc_0_wstrb_host_addr_3_reg),
          
          .desc_1_txn_type_reg(desc_1_txn_type_reg),
          .desc_1_size_reg(desc_1_size_reg),
          .desc_1_data_offset_reg(desc_1_data_offset_reg),
          .desc_1_data_host_addr_0_reg(desc_1_data_host_addr_0_reg),
          .desc_1_data_host_addr_1_reg(desc_1_data_host_addr_1_reg),
          .desc_1_data_host_addr_2_reg(desc_1_data_host_addr_2_reg),
          .desc_1_data_host_addr_3_reg(desc_1_data_host_addr_3_reg),
          .desc_1_wstrb_host_addr_0_reg(desc_1_wstrb_host_addr_0_reg),
          .desc_1_wstrb_host_addr_1_reg(desc_1_wstrb_host_addr_1_reg),
          .desc_1_wstrb_host_addr_2_reg(desc_1_wstrb_host_addr_2_reg),
          .desc_1_wstrb_host_addr_3_reg(desc_1_wstrb_host_addr_3_reg),
          
          .desc_2_txn_type_reg(desc_2_txn_type_reg),
          .desc_2_size_reg(desc_2_size_reg),
          .desc_2_data_offset_reg(desc_2_data_offset_reg),
          .desc_2_data_host_addr_0_reg(desc_2_data_host_addr_0_reg),
          .desc_2_data_host_addr_1_reg(desc_2_data_host_addr_1_reg),
          .desc_2_data_host_addr_2_reg(desc_2_data_host_addr_2_reg),
          .desc_2_data_host_addr_3_reg(desc_2_data_host_addr_3_reg),
          .desc_2_wstrb_host_addr_0_reg(desc_2_wstrb_host_addr_0_reg),
          .desc_2_wstrb_host_addr_1_reg(desc_2_wstrb_host_addr_1_reg),
          .desc_2_wstrb_host_addr_2_reg(desc_2_wstrb_host_addr_2_reg),
          .desc_2_wstrb_host_addr_3_reg(desc_2_wstrb_host_addr_3_reg),
          
          .desc_3_txn_type_reg(desc_3_txn_type_reg),
          .desc_3_size_reg(desc_3_size_reg),
          .desc_3_data_offset_reg(desc_3_data_offset_reg),
          .desc_3_data_host_addr_0_reg(desc_3_data_host_addr_0_reg),
          .desc_3_data_host_addr_1_reg(desc_3_data_host_addr_1_reg),
          .desc_3_data_host_addr_2_reg(desc_3_data_host_addr_2_reg),
          .desc_3_data_host_addr_3_reg(desc_3_data_host_addr_3_reg),
          .desc_3_wstrb_host_addr_0_reg(desc_3_wstrb_host_addr_0_reg),
          .desc_3_wstrb_host_addr_1_reg(desc_3_wstrb_host_addr_1_reg),
          .desc_3_wstrb_host_addr_2_reg(desc_3_wstrb_host_addr_2_reg),
          .desc_3_wstrb_host_addr_3_reg(desc_3_wstrb_host_addr_3_reg),
          
          .desc_4_txn_type_reg(desc_4_txn_type_reg),
          .desc_4_size_reg(desc_4_size_reg),
          .desc_4_data_offset_reg(desc_4_data_offset_reg),
          .desc_4_data_host_addr_0_reg(desc_4_data_host_addr_0_reg),
          .desc_4_data_host_addr_1_reg(desc_4_data_host_addr_1_reg),
          .desc_4_data_host_addr_2_reg(desc_4_data_host_addr_2_reg),
          .desc_4_data_host_addr_3_reg(desc_4_data_host_addr_3_reg),
          .desc_4_wstrb_host_addr_0_reg(desc_4_wstrb_host_addr_0_reg),
          .desc_4_wstrb_host_addr_1_reg(desc_4_wstrb_host_addr_1_reg),
          .desc_4_wstrb_host_addr_2_reg(desc_4_wstrb_host_addr_2_reg),
          .desc_4_wstrb_host_addr_3_reg(desc_4_wstrb_host_addr_3_reg),
          
          .desc_5_txn_type_reg(desc_5_txn_type_reg),
          .desc_5_size_reg(desc_5_size_reg),
          .desc_5_data_offset_reg(desc_5_data_offset_reg),
          .desc_5_data_host_addr_0_reg(desc_5_data_host_addr_0_reg),
          .desc_5_data_host_addr_1_reg(desc_5_data_host_addr_1_reg),
          .desc_5_data_host_addr_2_reg(desc_5_data_host_addr_2_reg),
          .desc_5_data_host_addr_3_reg(desc_5_data_host_addr_3_reg),
          .desc_5_wstrb_host_addr_0_reg(desc_5_wstrb_host_addr_0_reg),
          .desc_5_wstrb_host_addr_1_reg(desc_5_wstrb_host_addr_1_reg),
          .desc_5_wstrb_host_addr_2_reg(desc_5_wstrb_host_addr_2_reg),
          .desc_5_wstrb_host_addr_3_reg(desc_5_wstrb_host_addr_3_reg),
          
          
          .desc_6_txn_type_reg(desc_6_txn_type_reg),
          .desc_6_size_reg(desc_6_size_reg),
          .desc_6_data_offset_reg(desc_6_data_offset_reg),
          .desc_6_data_host_addr_0_reg(desc_6_data_host_addr_0_reg),
          .desc_6_data_host_addr_1_reg(desc_6_data_host_addr_1_reg),
          .desc_6_data_host_addr_2_reg(desc_6_data_host_addr_2_reg),
          .desc_6_data_host_addr_3_reg(desc_6_data_host_addr_3_reg),
          .desc_6_wstrb_host_addr_0_reg(desc_6_wstrb_host_addr_0_reg),
          .desc_6_wstrb_host_addr_1_reg(desc_6_wstrb_host_addr_1_reg),
          .desc_6_wstrb_host_addr_2_reg(desc_6_wstrb_host_addr_2_reg),
          .desc_6_wstrb_host_addr_3_reg(desc_6_wstrb_host_addr_3_reg),
          
          
          .desc_7_txn_type_reg(desc_7_txn_type_reg),
          .desc_7_size_reg(desc_7_size_reg),
          .desc_7_data_offset_reg(desc_7_data_offset_reg),
          .desc_7_data_host_addr_0_reg(desc_7_data_host_addr_0_reg),
          .desc_7_data_host_addr_1_reg(desc_7_data_host_addr_1_reg),
          .desc_7_data_host_addr_2_reg(desc_7_data_host_addr_2_reg),
          .desc_7_data_host_addr_3_reg(desc_7_data_host_addr_3_reg),
          .desc_7_wstrb_host_addr_0_reg(desc_7_wstrb_host_addr_0_reg),
          .desc_7_wstrb_host_addr_1_reg(desc_7_wstrb_host_addr_1_reg),
          .desc_7_wstrb_host_addr_2_reg(desc_7_wstrb_host_addr_2_reg),
          .desc_7_wstrb_host_addr_3_reg(desc_7_wstrb_host_addr_3_reg),
          
          .desc_8_txn_type_reg(desc_8_txn_type_reg),
          .desc_8_size_reg(desc_8_size_reg),
          .desc_8_data_offset_reg(desc_8_data_offset_reg),
          .desc_8_data_host_addr_0_reg(desc_8_data_host_addr_0_reg),
          .desc_8_data_host_addr_1_reg(desc_8_data_host_addr_1_reg),
          .desc_8_data_host_addr_2_reg(desc_8_data_host_addr_2_reg),
          .desc_8_data_host_addr_3_reg(desc_8_data_host_addr_3_reg),
          .desc_8_wstrb_host_addr_0_reg(desc_8_wstrb_host_addr_0_reg),
          .desc_8_wstrb_host_addr_1_reg(desc_8_wstrb_host_addr_1_reg),
          .desc_8_wstrb_host_addr_2_reg(desc_8_wstrb_host_addr_2_reg),
          .desc_8_wstrb_host_addr_3_reg(desc_8_wstrb_host_addr_3_reg),
          
          .desc_9_txn_type_reg(desc_9_txn_type_reg),
          .desc_9_size_reg(desc_9_size_reg),
          .desc_9_data_offset_reg(desc_9_data_offset_reg),
          .desc_9_data_host_addr_0_reg(desc_9_data_host_addr_0_reg),
          .desc_9_data_host_addr_1_reg(desc_9_data_host_addr_1_reg),
          .desc_9_data_host_addr_2_reg(desc_9_data_host_addr_2_reg),
          .desc_9_data_host_addr_3_reg(desc_9_data_host_addr_3_reg),
          .desc_9_wstrb_host_addr_0_reg(desc_9_wstrb_host_addr_0_reg),
          .desc_9_wstrb_host_addr_1_reg(desc_9_wstrb_host_addr_1_reg),
          .desc_9_wstrb_host_addr_2_reg(desc_9_wstrb_host_addr_2_reg),
          .desc_9_wstrb_host_addr_3_reg(desc_9_wstrb_host_addr_3_reg),
          
          .desc_10_txn_type_reg(desc_10_txn_type_reg),
          .desc_10_size_reg(desc_10_size_reg),
          .desc_10_data_offset_reg(desc_10_data_offset_reg),
          .desc_10_data_host_addr_0_reg(desc_10_data_host_addr_0_reg),
          .desc_10_data_host_addr_1_reg(desc_10_data_host_addr_1_reg),
          .desc_10_data_host_addr_2_reg(desc_10_data_host_addr_2_reg),
          .desc_10_data_host_addr_3_reg(desc_10_data_host_addr_3_reg),
          .desc_10_wstrb_host_addr_0_reg(desc_10_wstrb_host_addr_0_reg),
          .desc_10_wstrb_host_addr_1_reg(desc_10_wstrb_host_addr_1_reg),
          .desc_10_wstrb_host_addr_2_reg(desc_10_wstrb_host_addr_2_reg),
          .desc_10_wstrb_host_addr_3_reg(desc_10_wstrb_host_addr_3_reg),
          
          .desc_11_txn_type_reg(desc_11_txn_type_reg),
          .desc_11_size_reg(desc_11_size_reg),
          .desc_11_data_offset_reg(desc_11_data_offset_reg),
          .desc_11_data_host_addr_0_reg(desc_11_data_host_addr_0_reg),
          .desc_11_data_host_addr_1_reg(desc_11_data_host_addr_1_reg),
          .desc_11_data_host_addr_2_reg(desc_11_data_host_addr_2_reg),
          .desc_11_data_host_addr_3_reg(desc_11_data_host_addr_3_reg),
          .desc_11_wstrb_host_addr_0_reg(desc_11_wstrb_host_addr_0_reg),
          .desc_11_wstrb_host_addr_1_reg(desc_11_wstrb_host_addr_1_reg),
          .desc_11_wstrb_host_addr_2_reg(desc_11_wstrb_host_addr_2_reg),
          .desc_11_wstrb_host_addr_3_reg(desc_11_wstrb_host_addr_3_reg),
          
          
          .desc_12_txn_type_reg(desc_12_txn_type_reg),
          .desc_12_size_reg(desc_12_size_reg),
          .desc_12_data_offset_reg(desc_12_data_offset_reg),
          .desc_12_data_host_addr_0_reg(desc_12_data_host_addr_0_reg),
          .desc_12_data_host_addr_1_reg(desc_12_data_host_addr_1_reg),
          .desc_12_data_host_addr_2_reg(desc_12_data_host_addr_2_reg),
          .desc_12_data_host_addr_3_reg(desc_12_data_host_addr_3_reg),
          .desc_12_wstrb_host_addr_0_reg(desc_12_wstrb_host_addr_0_reg),
          .desc_12_wstrb_host_addr_1_reg(desc_12_wstrb_host_addr_1_reg),
          .desc_12_wstrb_host_addr_2_reg(desc_12_wstrb_host_addr_2_reg),
          .desc_12_wstrb_host_addr_3_reg(desc_12_wstrb_host_addr_3_reg),
          
          
          .desc_13_txn_type_reg(desc_13_txn_type_reg),
          .desc_13_size_reg(desc_13_size_reg),
          .desc_13_data_offset_reg(desc_13_data_offset_reg),
          .desc_13_data_host_addr_0_reg(desc_13_data_host_addr_0_reg),
          .desc_13_data_host_addr_1_reg(desc_13_data_host_addr_1_reg),
          .desc_13_data_host_addr_2_reg(desc_13_data_host_addr_2_reg),
          .desc_13_data_host_addr_3_reg(desc_13_data_host_addr_3_reg),
          .desc_13_wstrb_host_addr_0_reg(desc_13_wstrb_host_addr_0_reg),
          .desc_13_wstrb_host_addr_1_reg(desc_13_wstrb_host_addr_1_reg),
          .desc_13_wstrb_host_addr_2_reg(desc_13_wstrb_host_addr_2_reg),
          .desc_13_wstrb_host_addr_3_reg(desc_13_wstrb_host_addr_3_reg),
          
          .desc_14_txn_type_reg(desc_14_txn_type_reg),
          .desc_14_size_reg(desc_14_size_reg),
          .desc_14_data_offset_reg(desc_14_data_offset_reg),
          .desc_14_data_host_addr_0_reg(desc_14_data_host_addr_0_reg),
          .desc_14_data_host_addr_1_reg(desc_14_data_host_addr_1_reg),
          .desc_14_data_host_addr_2_reg(desc_14_data_host_addr_2_reg),
          .desc_14_data_host_addr_3_reg(desc_14_data_host_addr_3_reg),
          .desc_14_wstrb_host_addr_0_reg(desc_14_wstrb_host_addr_0_reg),
          .desc_14_wstrb_host_addr_1_reg(desc_14_wstrb_host_addr_1_reg),
          .desc_14_wstrb_host_addr_2_reg(desc_14_wstrb_host_addr_2_reg),
          .desc_14_wstrb_host_addr_3_reg(desc_14_wstrb_host_addr_3_reg),
          
          
          .desc_15_txn_type_reg(desc_15_txn_type_reg),
          .desc_15_size_reg(desc_15_size_reg),
          .desc_15_data_offset_reg(desc_15_data_offset_reg),
          .desc_15_data_host_addr_0_reg(desc_15_data_host_addr_0_reg),
          .desc_15_data_host_addr_1_reg(desc_15_data_host_addr_1_reg),
          .desc_15_data_host_addr_2_reg(desc_15_data_host_addr_2_reg),
          .desc_15_data_host_addr_3_reg(desc_15_data_host_addr_3_reg),
          .desc_15_wstrb_host_addr_0_reg(desc_15_wstrb_host_addr_0_reg),
          .desc_15_wstrb_host_addr_1_reg(desc_15_wstrb_host_addr_1_reg),
          .desc_15_wstrb_host_addr_2_reg(desc_15_wstrb_host_addr_2_reg),
          .desc_15_wstrb_host_addr_3_reg(desc_15_wstrb_host_addr_3_reg),


		  // M-AXI 
		  .m_axi_awid       (m_axi_awid    ), 
		  .m_axi_awaddr     (m_axi_awaddr  ), 
		  .m_axi_awlen      (m_axi_awlen   ), 
		  .m_axi_awsize     (m_axi_awsize  ), 
		  .m_axi_awburst    (m_axi_awburst ), 
		  .m_axi_awlock     (m_axi_awlock  ), 
		  .m_axi_awcache    (m_axi_awcache ), 
		  .m_axi_awprot     (m_axi_awprot  ), 
		  .m_axi_awqos      (m_axi_awqos   ), 
		  .m_axi_awregion   (m_axi_awregion), 
		  .m_axi_awuser     (m_axi_awuser  ), 
		  .m_axi_awvalid    (m_axi_awvalid ), 
		  .m_axi_awready    (m_axi_awready ), 
		  .m_axi_wdata      (m_axi_wdata   ), 
		  .m_axi_wstrb      (m_axi_wstrb   ), 
		  .m_axi_wlast      (m_axi_wlast   ), 
		  .m_axi_wuser      (m_axi_wuser   ), 
		  .m_axi_wvalid     (m_axi_wvalid  ), 
		  .m_axi_wready     (m_axi_wready  ), 
		  .m_axi_bid        (m_axi_bid     ), 
		  .m_axi_bresp      (m_axi_bresp   ), 
		  .m_axi_buser      (m_axi_buser   ), 
		  .m_axi_bvalid     (m_axi_bvalid  ), 
		  .m_axi_bready     (m_axi_bready  ), 
		  .m_axi_arid       (m_axi_arid    ), 
		  .m_axi_araddr     (m_axi_araddr  ), 
		  .m_axi_arlen      (m_axi_arlen   ), 
		  .m_axi_arsize     (m_axi_arsize  ), 
		  .m_axi_arburst    (m_axi_arburst ), 
		  .m_axi_arlock     (m_axi_arlock  ), 
		  .m_axi_arcache    (m_axi_arcache ), 
		  .m_axi_arprot     (m_axi_arprot  ), 
		  .m_axi_arqos      (m_axi_arqos   ), 
		  .m_axi_arregion   (m_axi_arregion), 
		  .m_axi_aruser     (m_axi_aruser  ), 
		  .m_axi_arvalid    (m_axi_arvalid ), 
		  .m_axi_arready    (m_axi_arready ), 
		  .m_axi_rid        (m_axi_rid     ), 
		  .m_axi_rdata      (m_axi_rdata   ), 
		  .m_axi_rresp      (m_axi_rresp   ), 
		  .m_axi_rlast      (m_axi_rlast   ), 
		  .m_axi_ruser      (m_axi_ruser   ), 
		  .m_axi_rvalid     (m_axi_rvalid  ), 
		  .m_axi_rready     (m_axi_rready  ), 


		  // Inputs
		  .version_reg          (version_reg),
		  .bridge_type_reg      (bridge_type_reg),
		  .axi_max_desc_reg     (axi_max_desc_reg),
		  
		  .uc2hm_trig           (uc2hm_trig),
		  .rb2hm_rd_dout        (rb2hm_rd_data),
          .rb2hm_rd_wstrb       (rb2hm_rd_wstrb));

   
   
   intr_handler_slave #(
                        .M_AXI_ADDR_WIDTH  (M_AXI_ADDR_WIDTH), 
                        .M_AXI_DATA_WIDTH  (M_AXI_DATA_WIDTH), 
                        .M_AXI_ID_WIDTH    (M_AXI_ID_WIDTH  ), 
                        .M_AXI_USER_WIDTH  (M_AXI_USER_WIDTH), 
                        .S_AXI_USR_DATA_WIDTH (S_AXI_USR_DATA_WIDTH),
                        .RAM_SIZE          (RAM_SIZE        ), 
                        .MAX_DESC          (MAX_DESC        ) 
) 
   intr_handler_slave_inst 
	 (
	  .axi_aclk                       (axi_aclk                      ), 
	  .axi_aresetn                    (rst_n                         ), 
	  .irq_out                        (irq_out                       ), 
	  .irq_ack                        (irq_ack                       ), 
	  .h2c_intr_out                   (h2c_intr_out                  ),
	  .h2c_gpio_out                   (h2c_gpio_out                  ),
	  .c2h_intr_in                    (c2h_intr_in                   ), 
	  .c2h_gpio_in                    (c2h_gpio_in                   ), 
	  .ih2rb_c2h_intr_status_0_reg    (ih2rb_c2h_intr_status_0_reg   ), 
	  .ih2rb_c2h_intr_status_1_reg    (ih2rb_c2h_intr_status_1_reg   ),
	  .ih2rb_intr_c2h_toggle_status_0_reg    (ih2rb_intr_c2h_toggle_status_0_reg   ), 
	  .ih2rb_intr_c2h_toggle_status_1_reg    (ih2rb_intr_c2h_toggle_status_1_reg   ),
	  .intr_c2h_toggle_clear_0_reg           (intr_c2h_toggle_clear_0_reg          ),
	  .intr_c2h_toggle_clear_1_reg           (intr_c2h_toggle_clear_1_reg          ),
	  .ih2rb_c2h_gpio_0_reg     (ih2rb_c2h_gpio_0_reg   ),
      .ih2rb_c2h_gpio_1_reg     (ih2rb_c2h_gpio_1_reg   ),
      .ih2rb_c2h_gpio_2_reg     (ih2rb_c2h_gpio_2_reg   ),
      .ih2rb_c2h_gpio_3_reg     (ih2rb_c2h_gpio_3_reg   ),
      .ih2rb_c2h_gpio_4_reg     (ih2rb_c2h_gpio_4_reg   ),
      .ih2rb_c2h_gpio_5_reg     (ih2rb_c2h_gpio_5_reg   ),
      .ih2rb_c2h_gpio_6_reg     (ih2rb_c2h_gpio_6_reg   ),
      .ih2rb_c2h_gpio_7_reg     (ih2rb_c2h_gpio_7_reg   ), 
	  .ih2rb_c2h_intr_status_0_reg_we (ih2rb_c2h_intr_status_0_reg_we), 
	  .ih2rb_c2h_intr_status_1_reg_we (ih2rb_c2h_intr_status_1_reg_we),
	  .ih2rb_intr_c2h_toggle_status_0_reg_we (ih2rb_intr_c2h_toggle_status_0_reg_we), 
	  .ih2rb_intr_c2h_toggle_status_1_reg_we (ih2rb_intr_c2h_toggle_status_1_reg_we), 
	  .ih2rb_c2h_gpio_0_reg_we  (ih2rb_c2h_gpio_0_reg_we),
      .ih2rb_c2h_gpio_1_reg_we  (ih2rb_c2h_gpio_1_reg_we),
	  .ih2rb_c2h_gpio_2_reg_we  (ih2rb_c2h_gpio_2_reg_we),
      .ih2rb_c2h_gpio_3_reg_we  (ih2rb_c2h_gpio_3_reg_we),
      .ih2rb_c2h_gpio_4_reg_we  (ih2rb_c2h_gpio_4_reg_we),
      .ih2rb_c2h_gpio_5_reg_we  (ih2rb_c2h_gpio_5_reg_we),
      .ih2rb_c2h_gpio_6_reg_we  (ih2rb_c2h_gpio_6_reg_we),
      .ih2rb_c2h_gpio_7_reg_we  (ih2rb_c2h_gpio_7_reg_we),
	  .version_reg                    (version_reg                   ), 
	  .bridge_type_reg                (bridge_type_reg               ), 
	  .mode_select_reg                (mode_select_reg               ), 
	  .reset_reg                      (reset_reg                     ), 
	  .h2c_intr_0_reg                 (h2c_intr_0_reg                ), 
	  .h2c_intr_1_reg                 (h2c_intr_1_reg                ),
	  .h2c_intr_2_reg                 (h2c_intr_2_reg                ), 
	  .h2c_intr_3_reg                 (h2c_intr_3_reg                ), 
	  .c2h_intr_status_0_reg          (c2h_intr_status_0_reg         ), 
	  .c2h_intr_status_1_reg          (c2h_intr_status_1_reg         ),
  	  .intr_c2h_toggle_status_0_reg   (intr_c2h_toggle_status_0_reg  ), 
	  .intr_c2h_toggle_status_1_reg   (intr_c2h_toggle_status_1_reg  ),
  	  .intr_c2h_toggle_enable_0_reg   (intr_c2h_toggle_enable_0_reg  ), 
	  .intr_c2h_toggle_enable_1_reg   (intr_c2h_toggle_enable_1_reg  ), 
	  .c2h_gpio_0_reg          (c2h_gpio_0_reg         ), 
	  .c2h_gpio_1_reg          (c2h_gpio_1_reg         ), 
	  .c2h_gpio_2_reg          (c2h_gpio_2_reg         ), 
	  .c2h_gpio_3_reg          (c2h_gpio_3_reg         ), 
	  .c2h_gpio_4_reg          (c2h_gpio_4_reg         ), 
	  .c2h_gpio_5_reg          (c2h_gpio_5_reg         ), 
	  .c2h_gpio_6_reg          (c2h_gpio_6_reg         ), 
	  .c2h_gpio_7_reg          (c2h_gpio_7_reg         ), 
	  .c2h_gpio_8_reg          (c2h_gpio_8_reg         ), 
	  .c2h_gpio_9_reg          (c2h_gpio_9_reg         ), 
	  .c2h_gpio_10_reg         (c2h_gpio_10_reg        ), 
	  .c2h_gpio_11_reg         (c2h_gpio_11_reg        ), 
	  .c2h_gpio_12_reg         (c2h_gpio_12_reg        ), 
	  .c2h_gpio_13_reg         (c2h_gpio_13_reg        ), 
	  .c2h_gpio_14_reg         (c2h_gpio_14_reg        ), 
	  .c2h_gpio_15_reg         (c2h_gpio_15_reg        ),
	  .h2c_gpio_0_reg          (h2c_gpio_0_reg         ), 
	  .h2c_gpio_1_reg          (h2c_gpio_1_reg         ), 
	  .h2c_gpio_2_reg          (h2c_gpio_2_reg         ), 
	  .h2c_gpio_3_reg          (h2c_gpio_3_reg         ), 
	  .h2c_gpio_4_reg          (h2c_gpio_4_reg         ), 
	  .h2c_gpio_5_reg          (h2c_gpio_5_reg         ), 
	  .h2c_gpio_6_reg          (h2c_gpio_6_reg         ), 
	  .h2c_gpio_7_reg          (h2c_gpio_7_reg         ), 
	  .axi_bridge_config_reg          (axi_bridge_config_reg         ), 
	  .axi_max_desc_reg               (axi_max_desc_reg              ), 
	  .intr_status_reg                (intr_status_reg               ), 
	  .intr_error_status_reg          (intr_error_status_reg         ), 
	  .intr_error_clear_reg           (intr_error_clear_reg          ), 
	  .intr_error_enable_reg          (intr_error_enable_reg         ), 
	  .ownership_reg                  (ownership_reg                 ), 
	  .ownership_flip_reg             (ownership_flip_reg            ), 
	  .status_resp_reg                (status_resp_reg               ), 
	  .intr_txn_avail_status_reg      (intr_txn_avail_status_reg     ), 
	  .intr_txn_avail_clear_reg       (intr_txn_avail_clear_reg      ), 
	  .intr_txn_avail_enable_reg      (intr_txn_avail_enable_reg     ),
	  .intr_comp_status_reg           (intr_comp_status_reg          ), 
	  .intr_comp_clear_reg            (intr_comp_clear_reg           ), 
	  .intr_comp_enable_reg           (intr_comp_enable_reg          ));



  endmodule 

// Local Variables:
// verilog-library-directories:("./")
// End:


