/*
 * Copyright (c) 2019 Xilinx Inc.
 * Written by Meera Bagdai. 
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy 
 * of this software and associated documentation files (the 'Software'), to deal 
 * in the Software without restriction, including without limitation the rights 
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
 * copies of the Software, and to permit persons to whom the Software is 
 * furnished to do so, subject to the following conditions: 
 * 
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED 'AS IS', WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 * 
 * Description: 
 *   This module is replica of user_slave_control module but it converts
 *   all registers into the internal fields as int_<reg>_<field> . Only these fields 
 *   are used in further hierarchy rather than registers.
 *
 *
 */

`include "defines_common.vh"

module user_slave_control_field #(

         parameter EN_INTFS_AXI4                                        =  1 
        ,parameter EN_INTFS_AXI4LITE                                    =  0 
        ,parameter EN_INTFS_AXI3                                        =  0 
                        
        ,parameter ADDR_WIDTH                                           = 64    
        ,parameter DATA_WIDTH                                           = 128
        ,parameter ID_WIDTH                                             = 16  
        ,parameter AWUSER_WIDTH                                         = 32    
        ,parameter WUSER_WIDTH                                          = 32    
        ,parameter BUSER_WIDTH                                          = 32    
        ,parameter ARUSER_WIDTH                                         = 32    
        ,parameter RUSER_WIDTH                                          = 32    
        ,parameter RAM_SIZE                                             = 16384  
        ,parameter MAX_DESC                                             = 16                   
        ,parameter FORCE_RESP_ORDER                                     = 1

)(

        //Clock and reset
         input 	     	                                                axi_aclk		
        ,input 	     	                                                axi_aresetn		
 		
        //S_AXI_USR
        ,input [ID_WIDTH-1:0]                                           s_axi_usr_awid
        ,input [ADDR_WIDTH-1:0]                                         s_axi_usr_awaddr
        ,input [7:0]                                                    s_axi_usr_awlen
        ,input [2:0]                                                    s_axi_usr_awsize
        ,input [1:0]                                                    s_axi_usr_awburst
        ,input [1:0]                                                    s_axi_usr_awlock
        ,input [3:0]                                                    s_axi_usr_awcache
        ,input [2:0]                                                    s_axi_usr_awprot
        ,input [3:0]                                                    s_axi_usr_awqos
        ,input [3:0]                                                    s_axi_usr_awregion 
        ,input [AWUSER_WIDTH-1:0]                                       s_axi_usr_awuser
        ,input                                                          s_axi_usr_awvalid
        ,output                                                         s_axi_usr_awready
        ,input [DATA_WIDTH-1:0]                                         s_axi_usr_wdata
        ,input [(DATA_WIDTH/8)-1:0]                                     s_axi_usr_wstrb
        ,input                                                          s_axi_usr_wlast
        ,input [ID_WIDTH-1:0]                                           s_axi_usr_wid
        ,input [WUSER_WIDTH-1:0]                                        s_axi_usr_wuser
        ,input                                                          s_axi_usr_wvalid
        ,output                                                         s_axi_usr_wready
        ,output [ID_WIDTH-1:0]                                          s_axi_usr_bid
        ,output [1:0]                                                   s_axi_usr_bresp
        ,output [BUSER_WIDTH-1:0]                                       s_axi_usr_buser
        ,output                                                         s_axi_usr_bvalid
        ,input                                                          s_axi_usr_bready
        ,input [ID_WIDTH-1:0]                                           s_axi_usr_arid
        ,input [ADDR_WIDTH-1:0]                                         s_axi_usr_araddr
        ,input [7:0]                                                    s_axi_usr_arlen
        ,input [2:0]                                                    s_axi_usr_arsize
        ,input [1:0]                                                    s_axi_usr_arburst
        ,input [1:0]                                                    s_axi_usr_arlock
        ,input [3:0]                                                    s_axi_usr_arcache
        ,input [2:0]                                                    s_axi_usr_arprot
        ,input [3:0]                                                    s_axi_usr_arqos
        ,input [3:0]                                                    s_axi_usr_arregion 
        ,input [ARUSER_WIDTH-1:0]                                       s_axi_usr_aruser
        ,input                                                          s_axi_usr_arvalid
        ,output                                                         s_axi_usr_arready
        ,output [ID_WIDTH-1:0]                                          s_axi_usr_rid
        ,output [DATA_WIDTH-1:0]                                        s_axi_usr_rdata
        ,output [1:0]                                                   s_axi_usr_rresp
        ,output                                                         s_axi_usr_rlast
        ,output [RUSER_WIDTH-1:0]                                       s_axi_usr_ruser
        ,output                                                         s_axi_usr_rvalid
        ,input                                                          s_axi_usr_rready

        ,input  [31:0]                                                  version_reg	
        ,input  [31:0]                                                  bridge_type_reg	
        ,input  [31:0]                                                  mode_select_reg	
        ,input  [31:0]                                                  reset_reg	
        ,input  [31:0]                                                  intr_h2c_0_reg	
        ,input  [31:0]                                                  intr_h2c_1_reg	
        ,input  [31:0]                                                  intr_c2h_0_status_reg	
        ,input  [31:0]                                                  intr_c2h_1_status_reg	
        ,input  [31:0]                                                  c2h_gpio_0_status_reg	
        ,input  [31:0]                                                  c2h_gpio_1_status_reg	
        ,input  [31:0]                                                  c2h_gpio_2_status_reg	
        ,input  [31:0]                                                  c2h_gpio_3_status_reg	
        ,input  [31:0]                                                  c2h_gpio_4_status_reg	
        ,input  [31:0]                                                  c2h_gpio_5_status_reg	
        ,input  [31:0]                                                  c2h_gpio_6_status_reg	
        ,input  [31:0]                                                  c2h_gpio_7_status_reg	
        ,input  [31:0]                                                  c2h_gpio_8_status_reg	
        ,input  [31:0]                                                  c2h_gpio_9_status_reg	
        ,input  [31:0]                                                  c2h_gpio_10_status_reg	
        ,input  [31:0]                                                  c2h_gpio_11_status_reg	
        ,input  [31:0]                                                  c2h_gpio_12_status_reg	
        ,input  [31:0]                                                  c2h_gpio_13_status_reg	
        ,input  [31:0]                                                  c2h_gpio_14_status_reg	
        ,input  [31:0]                                                  c2h_gpio_15_status_reg	
        ,input  [31:0]                                                  axi_bridge_config_reg	
        ,input  [31:0]                                                  axi_max_desc_reg	
        ,input  [31:0]                                                  intr_status_reg	
        ,input  [31:0]                                                  intr_error_status_reg	
        ,input  [31:0]                                                  intr_error_clear_reg	
        ,input  [31:0]                                                  intr_error_enable_reg	
        ,input  [31:0]                                                  addr_in_0_reg	
        ,input  [31:0]                                                  addr_in_1_reg	
        ,input  [31:0]                                                  addr_in_2_reg	
        ,input  [31:0]                                                  addr_in_3_reg	
        ,input  [31:0]                                                  trans_mask_0_reg	
        ,input  [31:0]                                                  trans_mask_1_reg	
        ,input  [31:0]                                                  trans_mask_2_reg	
        ,input  [31:0]                                                  trans_mask_3_reg	
        ,input  [31:0]                                                  trans_addr_0_reg	
        ,input  [31:0]                                                  trans_addr_1_reg	
        ,input  [31:0]                                                  trans_addr_2_reg	
        ,input  [31:0]                                                  trans_addr_3_reg	
        ,input  [31:0]                                                  ownership_reg	
        ,input  [31:0]                                                  ownership_flip_reg	
        ,input  [31:0]                                                  status_resp_reg	
        ,input  [31:0]                                                  intr_txn_avail_status_reg	
        ,input  [31:0]                                                  intr_txn_avail_clear_reg	
        ,input  [31:0]                                                  intr_txn_avail_enable_reg	
        ,input  [31:0]                                                  intr_comp_status_reg	
        ,input  [31:0]                                                  intr_comp_clear_reg	
        ,input  [31:0]                                                  intr_comp_enable_reg	
        ,input  [31:0]                                                  status_resp_comp_reg	
        ,input  [31:0]                                                  status_busy_reg	
        ,input  [31:0]                                                  resp_fifo_free_level_reg	
        ,input  [31:0]                                                  resp_order_reg
        ,input  [31:0]                                                  desc_0_txn_type_reg	
        ,input  [31:0]                                                  desc_0_size_reg	
        ,input  [31:0]                                                  desc_0_data_offset_reg	
        ,input  [31:0]                                                  desc_0_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_0_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_0_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_0_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_0_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_0_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_0_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_0_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_0_axsize_reg	
        ,input  [31:0]                                                  desc_0_attr_reg	
        ,input  [31:0]                                                  desc_0_axaddr_0_reg	
        ,input  [31:0]                                                  desc_0_axaddr_1_reg	
        ,input  [31:0]                                                  desc_0_axaddr_2_reg	
        ,input  [31:0]                                                  desc_0_axaddr_3_reg	
        ,input  [31:0]                                                  desc_0_axid_0_reg	
        ,input  [31:0]                                                  desc_0_axid_1_reg	
        ,input  [31:0]                                                  desc_0_axid_2_reg	
        ,input  [31:0]                                                  desc_0_axid_3_reg	
        ,input  [31:0]                                                  desc_0_axuser_0_reg	
        ,input  [31:0]                                                  desc_0_axuser_1_reg	
        ,input  [31:0]                                                  desc_0_axuser_2_reg	
        ,input  [31:0]                                                  desc_0_axuser_3_reg	
        ,input  [31:0]                                                  desc_0_axuser_4_reg	
        ,input  [31:0]                                                  desc_0_axuser_5_reg	
        ,input  [31:0]                                                  desc_0_axuser_6_reg	
        ,input  [31:0]                                                  desc_0_axuser_7_reg	
        ,input  [31:0]                                                  desc_0_axuser_8_reg	
        ,input  [31:0]                                                  desc_0_axuser_9_reg	
        ,input  [31:0]                                                  desc_0_axuser_10_reg	
        ,input  [31:0]                                                  desc_0_axuser_11_reg	
        ,input  [31:0]                                                  desc_0_axuser_12_reg	
        ,input  [31:0]                                                  desc_0_axuser_13_reg	
        ,input  [31:0]                                                  desc_0_axuser_14_reg	
        ,input  [31:0]                                                  desc_0_axuser_15_reg	
        ,input  [31:0]                                                  desc_0_xuser_0_reg	
        ,input  [31:0]                                                  desc_0_xuser_1_reg	
        ,input  [31:0]                                                  desc_0_xuser_2_reg	
        ,input  [31:0]                                                  desc_0_xuser_3_reg	
        ,input  [31:0]                                                  desc_0_xuser_4_reg	
        ,input  [31:0]                                                  desc_0_xuser_5_reg	
        ,input  [31:0]                                                  desc_0_xuser_6_reg	
        ,input  [31:0]                                                  desc_0_xuser_7_reg	
        ,input  [31:0]                                                  desc_0_xuser_8_reg	
        ,input  [31:0]                                                  desc_0_xuser_9_reg	
        ,input  [31:0]                                                  desc_0_xuser_10_reg	
        ,input  [31:0]                                                  desc_0_xuser_11_reg	
        ,input  [31:0]                                                  desc_0_xuser_12_reg	
        ,input  [31:0]                                                  desc_0_xuser_13_reg	
        ,input  [31:0]                                                  desc_0_xuser_14_reg	
        ,input  [31:0]                                                  desc_0_xuser_15_reg	
        ,input  [31:0]                                                  desc_0_wuser_0_reg	
        ,input  [31:0]                                                  desc_0_wuser_1_reg	
        ,input  [31:0]                                                  desc_0_wuser_2_reg	
        ,input  [31:0]                                                  desc_0_wuser_3_reg	
        ,input  [31:0]                                                  desc_0_wuser_4_reg	
        ,input  [31:0]                                                  desc_0_wuser_5_reg	
        ,input  [31:0]                                                  desc_0_wuser_6_reg	
        ,input  [31:0]                                                  desc_0_wuser_7_reg	
        ,input  [31:0]                                                  desc_0_wuser_8_reg	
        ,input  [31:0]                                                  desc_0_wuser_9_reg	
        ,input  [31:0]                                                  desc_0_wuser_10_reg	
        ,input  [31:0]                                                  desc_0_wuser_11_reg	
        ,input  [31:0]                                                  desc_0_wuser_12_reg	
        ,input  [31:0]                                                  desc_0_wuser_13_reg	
        ,input  [31:0]                                                  desc_0_wuser_14_reg	
        ,input  [31:0]                                                  desc_0_wuser_15_reg	
        ,input  [31:0]                                                  desc_1_txn_type_reg	
        ,input  [31:0]                                                  desc_1_size_reg	
        ,input  [31:0]                                                  desc_1_data_offset_reg	
        ,input  [31:0]                                                  desc_1_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_1_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_1_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_1_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_1_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_1_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_1_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_1_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_1_axsize_reg	
        ,input  [31:0]                                                  desc_1_attr_reg	
        ,input  [31:0]                                                  desc_1_axaddr_0_reg	
        ,input  [31:0]                                                  desc_1_axaddr_1_reg	
        ,input  [31:0]                                                  desc_1_axaddr_2_reg	
        ,input  [31:0]                                                  desc_1_axaddr_3_reg	
        ,input  [31:0]                                                  desc_1_axid_0_reg	
        ,input  [31:0]                                                  desc_1_axid_1_reg	
        ,input  [31:0]                                                  desc_1_axid_2_reg	
        ,input  [31:0]                                                  desc_1_axid_3_reg	
        ,input  [31:0]                                                  desc_1_axuser_0_reg	
        ,input  [31:0]                                                  desc_1_axuser_1_reg	
        ,input  [31:0]                                                  desc_1_axuser_2_reg	
        ,input  [31:0]                                                  desc_1_axuser_3_reg	
        ,input  [31:0]                                                  desc_1_axuser_4_reg	
        ,input  [31:0]                                                  desc_1_axuser_5_reg	
        ,input  [31:0]                                                  desc_1_axuser_6_reg	
        ,input  [31:0]                                                  desc_1_axuser_7_reg	
        ,input  [31:0]                                                  desc_1_axuser_8_reg	
        ,input  [31:0]                                                  desc_1_axuser_9_reg	
        ,input  [31:0]                                                  desc_1_axuser_10_reg	
        ,input  [31:0]                                                  desc_1_axuser_11_reg	
        ,input  [31:0]                                                  desc_1_axuser_12_reg	
        ,input  [31:0]                                                  desc_1_axuser_13_reg	
        ,input  [31:0]                                                  desc_1_axuser_14_reg	
        ,input  [31:0]                                                  desc_1_axuser_15_reg	
        ,input  [31:0]                                                  desc_1_xuser_0_reg	
        ,input  [31:0]                                                  desc_1_xuser_1_reg	
        ,input  [31:0]                                                  desc_1_xuser_2_reg	
        ,input  [31:0]                                                  desc_1_xuser_3_reg	
        ,input  [31:0]                                                  desc_1_xuser_4_reg	
        ,input  [31:0]                                                  desc_1_xuser_5_reg	
        ,input  [31:0]                                                  desc_1_xuser_6_reg	
        ,input  [31:0]                                                  desc_1_xuser_7_reg	
        ,input  [31:0]                                                  desc_1_xuser_8_reg	
        ,input  [31:0]                                                  desc_1_xuser_9_reg	
        ,input  [31:0]                                                  desc_1_xuser_10_reg	
        ,input  [31:0]                                                  desc_1_xuser_11_reg	
        ,input  [31:0]                                                  desc_1_xuser_12_reg	
        ,input  [31:0]                                                  desc_1_xuser_13_reg	
        ,input  [31:0]                                                  desc_1_xuser_14_reg	
        ,input  [31:0]                                                  desc_1_xuser_15_reg	
        ,input  [31:0]                                                  desc_1_wuser_0_reg	
        ,input  [31:0]                                                  desc_1_wuser_1_reg	
        ,input  [31:0]                                                  desc_1_wuser_2_reg	
        ,input  [31:0]                                                  desc_1_wuser_3_reg	
        ,input  [31:0]                                                  desc_1_wuser_4_reg	
        ,input  [31:0]                                                  desc_1_wuser_5_reg	
        ,input  [31:0]                                                  desc_1_wuser_6_reg	
        ,input  [31:0]                                                  desc_1_wuser_7_reg	
        ,input  [31:0]                                                  desc_1_wuser_8_reg	
        ,input  [31:0]                                                  desc_1_wuser_9_reg	
        ,input  [31:0]                                                  desc_1_wuser_10_reg	
        ,input  [31:0]                                                  desc_1_wuser_11_reg	
        ,input  [31:0]                                                  desc_1_wuser_12_reg	
        ,input  [31:0]                                                  desc_1_wuser_13_reg	
        ,input  [31:0]                                                  desc_1_wuser_14_reg	
        ,input  [31:0]                                                  desc_1_wuser_15_reg	
        ,input  [31:0]                                                  desc_2_txn_type_reg	
        ,input  [31:0]                                                  desc_2_size_reg	
        ,input  [31:0]                                                  desc_2_data_offset_reg	
        ,input  [31:0]                                                  desc_2_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_2_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_2_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_2_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_2_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_2_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_2_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_2_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_2_axsize_reg	
        ,input  [31:0]                                                  desc_2_attr_reg	
        ,input  [31:0]                                                  desc_2_axaddr_0_reg	
        ,input  [31:0]                                                  desc_2_axaddr_1_reg	
        ,input  [31:0]                                                  desc_2_axaddr_2_reg	
        ,input  [31:0]                                                  desc_2_axaddr_3_reg	
        ,input  [31:0]                                                  desc_2_axid_0_reg	
        ,input  [31:0]                                                  desc_2_axid_1_reg	
        ,input  [31:0]                                                  desc_2_axid_2_reg	
        ,input  [31:0]                                                  desc_2_axid_3_reg	
        ,input  [31:0]                                                  desc_2_axuser_0_reg	
        ,input  [31:0]                                                  desc_2_axuser_1_reg	
        ,input  [31:0]                                                  desc_2_axuser_2_reg	
        ,input  [31:0]                                                  desc_2_axuser_3_reg	
        ,input  [31:0]                                                  desc_2_axuser_4_reg	
        ,input  [31:0]                                                  desc_2_axuser_5_reg	
        ,input  [31:0]                                                  desc_2_axuser_6_reg	
        ,input  [31:0]                                                  desc_2_axuser_7_reg	
        ,input  [31:0]                                                  desc_2_axuser_8_reg	
        ,input  [31:0]                                                  desc_2_axuser_9_reg	
        ,input  [31:0]                                                  desc_2_axuser_10_reg	
        ,input  [31:0]                                                  desc_2_axuser_11_reg	
        ,input  [31:0]                                                  desc_2_axuser_12_reg	
        ,input  [31:0]                                                  desc_2_axuser_13_reg	
        ,input  [31:0]                                                  desc_2_axuser_14_reg	
        ,input  [31:0]                                                  desc_2_axuser_15_reg	
        ,input  [31:0]                                                  desc_2_xuser_0_reg	
        ,input  [31:0]                                                  desc_2_xuser_1_reg	
        ,input  [31:0]                                                  desc_2_xuser_2_reg	
        ,input  [31:0]                                                  desc_2_xuser_3_reg	
        ,input  [31:0]                                                  desc_2_xuser_4_reg	
        ,input  [31:0]                                                  desc_2_xuser_5_reg	
        ,input  [31:0]                                                  desc_2_xuser_6_reg	
        ,input  [31:0]                                                  desc_2_xuser_7_reg	
        ,input  [31:0]                                                  desc_2_xuser_8_reg	
        ,input  [31:0]                                                  desc_2_xuser_9_reg	
        ,input  [31:0]                                                  desc_2_xuser_10_reg	
        ,input  [31:0]                                                  desc_2_xuser_11_reg	
        ,input  [31:0]                                                  desc_2_xuser_12_reg	
        ,input  [31:0]                                                  desc_2_xuser_13_reg	
        ,input  [31:0]                                                  desc_2_xuser_14_reg	
        ,input  [31:0]                                                  desc_2_xuser_15_reg	
        ,input  [31:0]                                                  desc_2_wuser_0_reg	
        ,input  [31:0]                                                  desc_2_wuser_1_reg	
        ,input  [31:0]                                                  desc_2_wuser_2_reg	
        ,input  [31:0]                                                  desc_2_wuser_3_reg	
        ,input  [31:0]                                                  desc_2_wuser_4_reg	
        ,input  [31:0]                                                  desc_2_wuser_5_reg	
        ,input  [31:0]                                                  desc_2_wuser_6_reg	
        ,input  [31:0]                                                  desc_2_wuser_7_reg	
        ,input  [31:0]                                                  desc_2_wuser_8_reg	
        ,input  [31:0]                                                  desc_2_wuser_9_reg	
        ,input  [31:0]                                                  desc_2_wuser_10_reg	
        ,input  [31:0]                                                  desc_2_wuser_11_reg	
        ,input  [31:0]                                                  desc_2_wuser_12_reg	
        ,input  [31:0]                                                  desc_2_wuser_13_reg	
        ,input  [31:0]                                                  desc_2_wuser_14_reg	
        ,input  [31:0]                                                  desc_2_wuser_15_reg	
        ,input  [31:0]                                                  desc_3_txn_type_reg	
        ,input  [31:0]                                                  desc_3_size_reg	
        ,input  [31:0]                                                  desc_3_data_offset_reg	
        ,input  [31:0]                                                  desc_3_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_3_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_3_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_3_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_3_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_3_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_3_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_3_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_3_axsize_reg	
        ,input  [31:0]                                                  desc_3_attr_reg	
        ,input  [31:0]                                                  desc_3_axaddr_0_reg	
        ,input  [31:0]                                                  desc_3_axaddr_1_reg	
        ,input  [31:0]                                                  desc_3_axaddr_2_reg	
        ,input  [31:0]                                                  desc_3_axaddr_3_reg	
        ,input  [31:0]                                                  desc_3_axid_0_reg	
        ,input  [31:0]                                                  desc_3_axid_1_reg	
        ,input  [31:0]                                                  desc_3_axid_2_reg	
        ,input  [31:0]                                                  desc_3_axid_3_reg	
        ,input  [31:0]                                                  desc_3_axuser_0_reg	
        ,input  [31:0]                                                  desc_3_axuser_1_reg	
        ,input  [31:0]                                                  desc_3_axuser_2_reg	
        ,input  [31:0]                                                  desc_3_axuser_3_reg	
        ,input  [31:0]                                                  desc_3_axuser_4_reg	
        ,input  [31:0]                                                  desc_3_axuser_5_reg	
        ,input  [31:0]                                                  desc_3_axuser_6_reg	
        ,input  [31:0]                                                  desc_3_axuser_7_reg	
        ,input  [31:0]                                                  desc_3_axuser_8_reg	
        ,input  [31:0]                                                  desc_3_axuser_9_reg	
        ,input  [31:0]                                                  desc_3_axuser_10_reg	
        ,input  [31:0]                                                  desc_3_axuser_11_reg	
        ,input  [31:0]                                                  desc_3_axuser_12_reg	
        ,input  [31:0]                                                  desc_3_axuser_13_reg	
        ,input  [31:0]                                                  desc_3_axuser_14_reg	
        ,input  [31:0]                                                  desc_3_axuser_15_reg	
        ,input  [31:0]                                                  desc_3_xuser_0_reg	
        ,input  [31:0]                                                  desc_3_xuser_1_reg	
        ,input  [31:0]                                                  desc_3_xuser_2_reg	
        ,input  [31:0]                                                  desc_3_xuser_3_reg	
        ,input  [31:0]                                                  desc_3_xuser_4_reg	
        ,input  [31:0]                                                  desc_3_xuser_5_reg	
        ,input  [31:0]                                                  desc_3_xuser_6_reg	
        ,input  [31:0]                                                  desc_3_xuser_7_reg	
        ,input  [31:0]                                                  desc_3_xuser_8_reg	
        ,input  [31:0]                                                  desc_3_xuser_9_reg	
        ,input  [31:0]                                                  desc_3_xuser_10_reg	
        ,input  [31:0]                                                  desc_3_xuser_11_reg	
        ,input  [31:0]                                                  desc_3_xuser_12_reg	
        ,input  [31:0]                                                  desc_3_xuser_13_reg	
        ,input  [31:0]                                                  desc_3_xuser_14_reg	
        ,input  [31:0]                                                  desc_3_xuser_15_reg	
        ,input  [31:0]                                                  desc_3_wuser_0_reg	
        ,input  [31:0]                                                  desc_3_wuser_1_reg	
        ,input  [31:0]                                                  desc_3_wuser_2_reg	
        ,input  [31:0]                                                  desc_3_wuser_3_reg	
        ,input  [31:0]                                                  desc_3_wuser_4_reg	
        ,input  [31:0]                                                  desc_3_wuser_5_reg	
        ,input  [31:0]                                                  desc_3_wuser_6_reg	
        ,input  [31:0]                                                  desc_3_wuser_7_reg	
        ,input  [31:0]                                                  desc_3_wuser_8_reg	
        ,input  [31:0]                                                  desc_3_wuser_9_reg	
        ,input  [31:0]                                                  desc_3_wuser_10_reg	
        ,input  [31:0]                                                  desc_3_wuser_11_reg	
        ,input  [31:0]                                                  desc_3_wuser_12_reg	
        ,input  [31:0]                                                  desc_3_wuser_13_reg	
        ,input  [31:0]                                                  desc_3_wuser_14_reg	
        ,input  [31:0]                                                  desc_3_wuser_15_reg	
        ,input  [31:0]                                                  desc_4_txn_type_reg	
        ,input  [31:0]                                                  desc_4_size_reg	
        ,input  [31:0]                                                  desc_4_data_offset_reg	
        ,input  [31:0]                                                  desc_4_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_4_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_4_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_4_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_4_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_4_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_4_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_4_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_4_axsize_reg	
        ,input  [31:0]                                                  desc_4_attr_reg	
        ,input  [31:0]                                                  desc_4_axaddr_0_reg	
        ,input  [31:0]                                                  desc_4_axaddr_1_reg	
        ,input  [31:0]                                                  desc_4_axaddr_2_reg	
        ,input  [31:0]                                                  desc_4_axaddr_3_reg	
        ,input  [31:0]                                                  desc_4_axid_0_reg	
        ,input  [31:0]                                                  desc_4_axid_1_reg	
        ,input  [31:0]                                                  desc_4_axid_2_reg	
        ,input  [31:0]                                                  desc_4_axid_3_reg	
        ,input  [31:0]                                                  desc_4_axuser_0_reg	
        ,input  [31:0]                                                  desc_4_axuser_1_reg	
        ,input  [31:0]                                                  desc_4_axuser_2_reg	
        ,input  [31:0]                                                  desc_4_axuser_3_reg	
        ,input  [31:0]                                                  desc_4_axuser_4_reg	
        ,input  [31:0]                                                  desc_4_axuser_5_reg	
        ,input  [31:0]                                                  desc_4_axuser_6_reg	
        ,input  [31:0]                                                  desc_4_axuser_7_reg	
        ,input  [31:0]                                                  desc_4_axuser_8_reg	
        ,input  [31:0]                                                  desc_4_axuser_9_reg	
        ,input  [31:0]                                                  desc_4_axuser_10_reg	
        ,input  [31:0]                                                  desc_4_axuser_11_reg	
        ,input  [31:0]                                                  desc_4_axuser_12_reg	
        ,input  [31:0]                                                  desc_4_axuser_13_reg	
        ,input  [31:0]                                                  desc_4_axuser_14_reg	
        ,input  [31:0]                                                  desc_4_axuser_15_reg	
        ,input  [31:0]                                                  desc_4_xuser_0_reg	
        ,input  [31:0]                                                  desc_4_xuser_1_reg	
        ,input  [31:0]                                                  desc_4_xuser_2_reg	
        ,input  [31:0]                                                  desc_4_xuser_3_reg	
        ,input  [31:0]                                                  desc_4_xuser_4_reg	
        ,input  [31:0]                                                  desc_4_xuser_5_reg	
        ,input  [31:0]                                                  desc_4_xuser_6_reg	
        ,input  [31:0]                                                  desc_4_xuser_7_reg	
        ,input  [31:0]                                                  desc_4_xuser_8_reg	
        ,input  [31:0]                                                  desc_4_xuser_9_reg	
        ,input  [31:0]                                                  desc_4_xuser_10_reg	
        ,input  [31:0]                                                  desc_4_xuser_11_reg	
        ,input  [31:0]                                                  desc_4_xuser_12_reg	
        ,input  [31:0]                                                  desc_4_xuser_13_reg	
        ,input  [31:0]                                                  desc_4_xuser_14_reg	
        ,input  [31:0]                                                  desc_4_xuser_15_reg	
        ,input  [31:0]                                                  desc_4_wuser_0_reg	
        ,input  [31:0]                                                  desc_4_wuser_1_reg	
        ,input  [31:0]                                                  desc_4_wuser_2_reg	
        ,input  [31:0]                                                  desc_4_wuser_3_reg	
        ,input  [31:0]                                                  desc_4_wuser_4_reg	
        ,input  [31:0]                                                  desc_4_wuser_5_reg	
        ,input  [31:0]                                                  desc_4_wuser_6_reg	
        ,input  [31:0]                                                  desc_4_wuser_7_reg	
        ,input  [31:0]                                                  desc_4_wuser_8_reg	
        ,input  [31:0]                                                  desc_4_wuser_9_reg	
        ,input  [31:0]                                                  desc_4_wuser_10_reg	
        ,input  [31:0]                                                  desc_4_wuser_11_reg	
        ,input  [31:0]                                                  desc_4_wuser_12_reg	
        ,input  [31:0]                                                  desc_4_wuser_13_reg	
        ,input  [31:0]                                                  desc_4_wuser_14_reg	
        ,input  [31:0]                                                  desc_4_wuser_15_reg	
        ,input  [31:0]                                                  desc_5_txn_type_reg	
        ,input  [31:0]                                                  desc_5_size_reg	
        ,input  [31:0]                                                  desc_5_data_offset_reg	
        ,input  [31:0]                                                  desc_5_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_5_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_5_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_5_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_5_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_5_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_5_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_5_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_5_axsize_reg	
        ,input  [31:0]                                                  desc_5_attr_reg	
        ,input  [31:0]                                                  desc_5_axaddr_0_reg	
        ,input  [31:0]                                                  desc_5_axaddr_1_reg	
        ,input  [31:0]                                                  desc_5_axaddr_2_reg	
        ,input  [31:0]                                                  desc_5_axaddr_3_reg	
        ,input  [31:0]                                                  desc_5_axid_0_reg	
        ,input  [31:0]                                                  desc_5_axid_1_reg	
        ,input  [31:0]                                                  desc_5_axid_2_reg	
        ,input  [31:0]                                                  desc_5_axid_3_reg	
        ,input  [31:0]                                                  desc_5_axuser_0_reg	
        ,input  [31:0]                                                  desc_5_axuser_1_reg	
        ,input  [31:0]                                                  desc_5_axuser_2_reg	
        ,input  [31:0]                                                  desc_5_axuser_3_reg	
        ,input  [31:0]                                                  desc_5_axuser_4_reg	
        ,input  [31:0]                                                  desc_5_axuser_5_reg	
        ,input  [31:0]                                                  desc_5_axuser_6_reg	
        ,input  [31:0]                                                  desc_5_axuser_7_reg	
        ,input  [31:0]                                                  desc_5_axuser_8_reg	
        ,input  [31:0]                                                  desc_5_axuser_9_reg	
        ,input  [31:0]                                                  desc_5_axuser_10_reg	
        ,input  [31:0]                                                  desc_5_axuser_11_reg	
        ,input  [31:0]                                                  desc_5_axuser_12_reg	
        ,input  [31:0]                                                  desc_5_axuser_13_reg	
        ,input  [31:0]                                                  desc_5_axuser_14_reg	
        ,input  [31:0]                                                  desc_5_axuser_15_reg	
        ,input  [31:0]                                                  desc_5_xuser_0_reg	
        ,input  [31:0]                                                  desc_5_xuser_1_reg	
        ,input  [31:0]                                                  desc_5_xuser_2_reg	
        ,input  [31:0]                                                  desc_5_xuser_3_reg	
        ,input  [31:0]                                                  desc_5_xuser_4_reg	
        ,input  [31:0]                                                  desc_5_xuser_5_reg	
        ,input  [31:0]                                                  desc_5_xuser_6_reg	
        ,input  [31:0]                                                  desc_5_xuser_7_reg	
        ,input  [31:0]                                                  desc_5_xuser_8_reg	
        ,input  [31:0]                                                  desc_5_xuser_9_reg	
        ,input  [31:0]                                                  desc_5_xuser_10_reg	
        ,input  [31:0]                                                  desc_5_xuser_11_reg	
        ,input  [31:0]                                                  desc_5_xuser_12_reg	
        ,input  [31:0]                                                  desc_5_xuser_13_reg	
        ,input  [31:0]                                                  desc_5_xuser_14_reg	
        ,input  [31:0]                                                  desc_5_xuser_15_reg	
        ,input  [31:0]                                                  desc_5_wuser_0_reg	
        ,input  [31:0]                                                  desc_5_wuser_1_reg	
        ,input  [31:0]                                                  desc_5_wuser_2_reg	
        ,input  [31:0]                                                  desc_5_wuser_3_reg	
        ,input  [31:0]                                                  desc_5_wuser_4_reg	
        ,input  [31:0]                                                  desc_5_wuser_5_reg	
        ,input  [31:0]                                                  desc_5_wuser_6_reg	
        ,input  [31:0]                                                  desc_5_wuser_7_reg	
        ,input  [31:0]                                                  desc_5_wuser_8_reg	
        ,input  [31:0]                                                  desc_5_wuser_9_reg	
        ,input  [31:0]                                                  desc_5_wuser_10_reg	
        ,input  [31:0]                                                  desc_5_wuser_11_reg	
        ,input  [31:0]                                                  desc_5_wuser_12_reg	
        ,input  [31:0]                                                  desc_5_wuser_13_reg	
        ,input  [31:0]                                                  desc_5_wuser_14_reg	
        ,input  [31:0]                                                  desc_5_wuser_15_reg	
        ,input  [31:0]                                                  desc_6_txn_type_reg	
        ,input  [31:0]                                                  desc_6_size_reg	
        ,input  [31:0]                                                  desc_6_data_offset_reg	
        ,input  [31:0]                                                  desc_6_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_6_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_6_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_6_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_6_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_6_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_6_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_6_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_6_axsize_reg	
        ,input  [31:0]                                                  desc_6_attr_reg	
        ,input  [31:0]                                                  desc_6_axaddr_0_reg	
        ,input  [31:0]                                                  desc_6_axaddr_1_reg	
        ,input  [31:0]                                                  desc_6_axaddr_2_reg	
        ,input  [31:0]                                                  desc_6_axaddr_3_reg	
        ,input  [31:0]                                                  desc_6_axid_0_reg	
        ,input  [31:0]                                                  desc_6_axid_1_reg	
        ,input  [31:0]                                                  desc_6_axid_2_reg	
        ,input  [31:0]                                                  desc_6_axid_3_reg	
        ,input  [31:0]                                                  desc_6_axuser_0_reg	
        ,input  [31:0]                                                  desc_6_axuser_1_reg	
        ,input  [31:0]                                                  desc_6_axuser_2_reg	
        ,input  [31:0]                                                  desc_6_axuser_3_reg	
        ,input  [31:0]                                                  desc_6_axuser_4_reg	
        ,input  [31:0]                                                  desc_6_axuser_5_reg	
        ,input  [31:0]                                                  desc_6_axuser_6_reg	
        ,input  [31:0]                                                  desc_6_axuser_7_reg	
        ,input  [31:0]                                                  desc_6_axuser_8_reg	
        ,input  [31:0]                                                  desc_6_axuser_9_reg	
        ,input  [31:0]                                                  desc_6_axuser_10_reg	
        ,input  [31:0]                                                  desc_6_axuser_11_reg	
        ,input  [31:0]                                                  desc_6_axuser_12_reg	
        ,input  [31:0]                                                  desc_6_axuser_13_reg	
        ,input  [31:0]                                                  desc_6_axuser_14_reg	
        ,input  [31:0]                                                  desc_6_axuser_15_reg	
        ,input  [31:0]                                                  desc_6_xuser_0_reg	
        ,input  [31:0]                                                  desc_6_xuser_1_reg	
        ,input  [31:0]                                                  desc_6_xuser_2_reg	
        ,input  [31:0]                                                  desc_6_xuser_3_reg	
        ,input  [31:0]                                                  desc_6_xuser_4_reg	
        ,input  [31:0]                                                  desc_6_xuser_5_reg	
        ,input  [31:0]                                                  desc_6_xuser_6_reg	
        ,input  [31:0]                                                  desc_6_xuser_7_reg	
        ,input  [31:0]                                                  desc_6_xuser_8_reg	
        ,input  [31:0]                                                  desc_6_xuser_9_reg	
        ,input  [31:0]                                                  desc_6_xuser_10_reg	
        ,input  [31:0]                                                  desc_6_xuser_11_reg	
        ,input  [31:0]                                                  desc_6_xuser_12_reg	
        ,input  [31:0]                                                  desc_6_xuser_13_reg	
        ,input  [31:0]                                                  desc_6_xuser_14_reg	
        ,input  [31:0]                                                  desc_6_xuser_15_reg	
        ,input  [31:0]                                                  desc_6_wuser_0_reg	
        ,input  [31:0]                                                  desc_6_wuser_1_reg	
        ,input  [31:0]                                                  desc_6_wuser_2_reg	
        ,input  [31:0]                                                  desc_6_wuser_3_reg	
        ,input  [31:0]                                                  desc_6_wuser_4_reg	
        ,input  [31:0]                                                  desc_6_wuser_5_reg	
        ,input  [31:0]                                                  desc_6_wuser_6_reg	
        ,input  [31:0]                                                  desc_6_wuser_7_reg	
        ,input  [31:0]                                                  desc_6_wuser_8_reg	
        ,input  [31:0]                                                  desc_6_wuser_9_reg	
        ,input  [31:0]                                                  desc_6_wuser_10_reg	
        ,input  [31:0]                                                  desc_6_wuser_11_reg	
        ,input  [31:0]                                                  desc_6_wuser_12_reg	
        ,input  [31:0]                                                  desc_6_wuser_13_reg	
        ,input  [31:0]                                                  desc_6_wuser_14_reg	
        ,input  [31:0]                                                  desc_6_wuser_15_reg	
        ,input  [31:0]                                                  desc_7_txn_type_reg	
        ,input  [31:0]                                                  desc_7_size_reg	
        ,input  [31:0]                                                  desc_7_data_offset_reg	
        ,input  [31:0]                                                  desc_7_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_7_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_7_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_7_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_7_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_7_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_7_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_7_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_7_axsize_reg	
        ,input  [31:0]                                                  desc_7_attr_reg	
        ,input  [31:0]                                                  desc_7_axaddr_0_reg	
        ,input  [31:0]                                                  desc_7_axaddr_1_reg	
        ,input  [31:0]                                                  desc_7_axaddr_2_reg	
        ,input  [31:0]                                                  desc_7_axaddr_3_reg	
        ,input  [31:0]                                                  desc_7_axid_0_reg	
        ,input  [31:0]                                                  desc_7_axid_1_reg	
        ,input  [31:0]                                                  desc_7_axid_2_reg	
        ,input  [31:0]                                                  desc_7_axid_3_reg	
        ,input  [31:0]                                                  desc_7_axuser_0_reg	
        ,input  [31:0]                                                  desc_7_axuser_1_reg	
        ,input  [31:0]                                                  desc_7_axuser_2_reg	
        ,input  [31:0]                                                  desc_7_axuser_3_reg	
        ,input  [31:0]                                                  desc_7_axuser_4_reg	
        ,input  [31:0]                                                  desc_7_axuser_5_reg	
        ,input  [31:0]                                                  desc_7_axuser_6_reg	
        ,input  [31:0]                                                  desc_7_axuser_7_reg	
        ,input  [31:0]                                                  desc_7_axuser_8_reg	
        ,input  [31:0]                                                  desc_7_axuser_9_reg	
        ,input  [31:0]                                                  desc_7_axuser_10_reg	
        ,input  [31:0]                                                  desc_7_axuser_11_reg	
        ,input  [31:0]                                                  desc_7_axuser_12_reg	
        ,input  [31:0]                                                  desc_7_axuser_13_reg	
        ,input  [31:0]                                                  desc_7_axuser_14_reg	
        ,input  [31:0]                                                  desc_7_axuser_15_reg	
        ,input  [31:0]                                                  desc_7_xuser_0_reg	
        ,input  [31:0]                                                  desc_7_xuser_1_reg	
        ,input  [31:0]                                                  desc_7_xuser_2_reg	
        ,input  [31:0]                                                  desc_7_xuser_3_reg	
        ,input  [31:0]                                                  desc_7_xuser_4_reg	
        ,input  [31:0]                                                  desc_7_xuser_5_reg	
        ,input  [31:0]                                                  desc_7_xuser_6_reg	
        ,input  [31:0]                                                  desc_7_xuser_7_reg	
        ,input  [31:0]                                                  desc_7_xuser_8_reg	
        ,input  [31:0]                                                  desc_7_xuser_9_reg	
        ,input  [31:0]                                                  desc_7_xuser_10_reg	
        ,input  [31:0]                                                  desc_7_xuser_11_reg	
        ,input  [31:0]                                                  desc_7_xuser_12_reg	
        ,input  [31:0]                                                  desc_7_xuser_13_reg	
        ,input  [31:0]                                                  desc_7_xuser_14_reg	
        ,input  [31:0]                                                  desc_7_xuser_15_reg	
        ,input  [31:0]                                                  desc_7_wuser_0_reg	
        ,input  [31:0]                                                  desc_7_wuser_1_reg	
        ,input  [31:0]                                                  desc_7_wuser_2_reg	
        ,input  [31:0]                                                  desc_7_wuser_3_reg	
        ,input  [31:0]                                                  desc_7_wuser_4_reg	
        ,input  [31:0]                                                  desc_7_wuser_5_reg	
        ,input  [31:0]                                                  desc_7_wuser_6_reg	
        ,input  [31:0]                                                  desc_7_wuser_7_reg	
        ,input  [31:0]                                                  desc_7_wuser_8_reg	
        ,input  [31:0]                                                  desc_7_wuser_9_reg	
        ,input  [31:0]                                                  desc_7_wuser_10_reg	
        ,input  [31:0]                                                  desc_7_wuser_11_reg	
        ,input  [31:0]                                                  desc_7_wuser_12_reg	
        ,input  [31:0]                                                  desc_7_wuser_13_reg	
        ,input  [31:0]                                                  desc_7_wuser_14_reg	
        ,input  [31:0]                                                  desc_7_wuser_15_reg	
        ,input  [31:0]                                                  desc_8_txn_type_reg	
        ,input  [31:0]                                                  desc_8_size_reg	
        ,input  [31:0]                                                  desc_8_data_offset_reg	
        ,input  [31:0]                                                  desc_8_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_8_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_8_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_8_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_8_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_8_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_8_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_8_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_8_axsize_reg	
        ,input  [31:0]                                                  desc_8_attr_reg	
        ,input  [31:0]                                                  desc_8_axaddr_0_reg	
        ,input  [31:0]                                                  desc_8_axaddr_1_reg	
        ,input  [31:0]                                                  desc_8_axaddr_2_reg	
        ,input  [31:0]                                                  desc_8_axaddr_3_reg	
        ,input  [31:0]                                                  desc_8_axid_0_reg	
        ,input  [31:0]                                                  desc_8_axid_1_reg	
        ,input  [31:0]                                                  desc_8_axid_2_reg	
        ,input  [31:0]                                                  desc_8_axid_3_reg	
        ,input  [31:0]                                                  desc_8_axuser_0_reg	
        ,input  [31:0]                                                  desc_8_axuser_1_reg	
        ,input  [31:0]                                                  desc_8_axuser_2_reg	
        ,input  [31:0]                                                  desc_8_axuser_3_reg	
        ,input  [31:0]                                                  desc_8_axuser_4_reg	
        ,input  [31:0]                                                  desc_8_axuser_5_reg	
        ,input  [31:0]                                                  desc_8_axuser_6_reg	
        ,input  [31:0]                                                  desc_8_axuser_7_reg	
        ,input  [31:0]                                                  desc_8_axuser_8_reg	
        ,input  [31:0]                                                  desc_8_axuser_9_reg	
        ,input  [31:0]                                                  desc_8_axuser_10_reg	
        ,input  [31:0]                                                  desc_8_axuser_11_reg	
        ,input  [31:0]                                                  desc_8_axuser_12_reg	
        ,input  [31:0]                                                  desc_8_axuser_13_reg	
        ,input  [31:0]                                                  desc_8_axuser_14_reg	
        ,input  [31:0]                                                  desc_8_axuser_15_reg	
        ,input  [31:0]                                                  desc_8_xuser_0_reg	
        ,input  [31:0]                                                  desc_8_xuser_1_reg	
        ,input  [31:0]                                                  desc_8_xuser_2_reg	
        ,input  [31:0]                                                  desc_8_xuser_3_reg	
        ,input  [31:0]                                                  desc_8_xuser_4_reg	
        ,input  [31:0]                                                  desc_8_xuser_5_reg	
        ,input  [31:0]                                                  desc_8_xuser_6_reg	
        ,input  [31:0]                                                  desc_8_xuser_7_reg	
        ,input  [31:0]                                                  desc_8_xuser_8_reg	
        ,input  [31:0]                                                  desc_8_xuser_9_reg	
        ,input  [31:0]                                                  desc_8_xuser_10_reg	
        ,input  [31:0]                                                  desc_8_xuser_11_reg	
        ,input  [31:0]                                                  desc_8_xuser_12_reg	
        ,input  [31:0]                                                  desc_8_xuser_13_reg	
        ,input  [31:0]                                                  desc_8_xuser_14_reg	
        ,input  [31:0]                                                  desc_8_xuser_15_reg	
        ,input  [31:0]                                                  desc_8_wuser_0_reg	
        ,input  [31:0]                                                  desc_8_wuser_1_reg	
        ,input  [31:0]                                                  desc_8_wuser_2_reg	
        ,input  [31:0]                                                  desc_8_wuser_3_reg	
        ,input  [31:0]                                                  desc_8_wuser_4_reg	
        ,input  [31:0]                                                  desc_8_wuser_5_reg	
        ,input  [31:0]                                                  desc_8_wuser_6_reg	
        ,input  [31:0]                                                  desc_8_wuser_7_reg	
        ,input  [31:0]                                                  desc_8_wuser_8_reg	
        ,input  [31:0]                                                  desc_8_wuser_9_reg	
        ,input  [31:0]                                                  desc_8_wuser_10_reg	
        ,input  [31:0]                                                  desc_8_wuser_11_reg	
        ,input  [31:0]                                                  desc_8_wuser_12_reg	
        ,input  [31:0]                                                  desc_8_wuser_13_reg	
        ,input  [31:0]                                                  desc_8_wuser_14_reg	
        ,input  [31:0]                                                  desc_8_wuser_15_reg	
        ,input  [31:0]                                                  desc_9_txn_type_reg	
        ,input  [31:0]                                                  desc_9_size_reg	
        ,input  [31:0]                                                  desc_9_data_offset_reg	
        ,input  [31:0]                                                  desc_9_data_host_addr_0_reg	
        ,input  [31:0]                                                  desc_9_data_host_addr_1_reg	
        ,input  [31:0]                                                  desc_9_data_host_addr_2_reg	
        ,input  [31:0]                                                  desc_9_data_host_addr_3_reg	
        ,input  [31:0]                                                  desc_9_wstrb_host_addr_0_reg	
        ,input  [31:0]                                                  desc_9_wstrb_host_addr_1_reg	
        ,input  [31:0]                                                  desc_9_wstrb_host_addr_2_reg	
        ,input  [31:0]                                                  desc_9_wstrb_host_addr_3_reg	
        ,input  [31:0]                                                  desc_9_axsize_reg	
        ,input  [31:0]                                                  desc_9_attr_reg	
        ,input  [31:0]                                                  desc_9_axaddr_0_reg	
        ,input  [31:0]                                                  desc_9_axaddr_1_reg	
        ,input  [31:0]                                                  desc_9_axaddr_2_reg	
        ,input  [31:0]                                                  desc_9_axaddr_3_reg	
        ,input  [31:0]                                                  desc_9_axid_0_reg	
        ,input  [31:0]                                                  desc_9_axid_1_reg	
        ,input  [31:0]                                                  desc_9_axid_2_reg	
        ,input  [31:0]                                                  desc_9_axid_3_reg	
        ,input  [31:0]                                                  desc_9_axuser_0_reg	
        ,input  [31:0]                                                  desc_9_axuser_1_reg	
        ,input  [31:0]                                                  desc_9_axuser_2_reg	
        ,input  [31:0]                                                  desc_9_axuser_3_reg	
        ,input  [31:0]                                                  desc_9_axuser_4_reg	
        ,input  [31:0]                                                  desc_9_axuser_5_reg	
        ,input  [31:0]                                                  desc_9_axuser_6_reg	
        ,input  [31:0]                                                  desc_9_axuser_7_reg	
        ,input  [31:0]                                                  desc_9_axuser_8_reg	
        ,input  [31:0]                                                  desc_9_axuser_9_reg	
        ,input  [31:0]                                                  desc_9_axuser_10_reg	
        ,input  [31:0]                                                  desc_9_axuser_11_reg	
        ,input  [31:0]                                                  desc_9_axuser_12_reg	
        ,input  [31:0]                                                  desc_9_axuser_13_reg	
        ,input  [31:0]                                                  desc_9_axuser_14_reg	
        ,input  [31:0]                                                  desc_9_axuser_15_reg	
        ,input  [31:0]                                                  desc_9_xuser_0_reg	
        ,input  [31:0]                                                  desc_9_xuser_1_reg	
        ,input  [31:0]                                                  desc_9_xuser_2_reg	
        ,input  [31:0]                                                  desc_9_xuser_3_reg	
        ,input  [31:0]                                                  desc_9_xuser_4_reg	
        ,input  [31:0]                                                  desc_9_xuser_5_reg	
        ,input  [31:0]                                                  desc_9_xuser_6_reg	
        ,input  [31:0]                                                  desc_9_xuser_7_reg	
        ,input  [31:0]                                                  desc_9_xuser_8_reg	
        ,input  [31:0]                                                  desc_9_xuser_9_reg	
        ,input  [31:0]                                                  desc_9_xuser_10_reg	
        ,input  [31:0]                                                  desc_9_xuser_11_reg	
        ,input  [31:0]                                                  desc_9_xuser_12_reg	
        ,input  [31:0]                                                  desc_9_xuser_13_reg	
        ,input  [31:0]                                                  desc_9_xuser_14_reg	
        ,input  [31:0]                                                  desc_9_xuser_15_reg	
        ,input  [31:0]                                                  desc_9_wuser_0_reg	
        ,input  [31:0]                                                  desc_9_wuser_1_reg	
        ,input  [31:0]                                                  desc_9_wuser_2_reg	
        ,input  [31:0]                                                  desc_9_wuser_3_reg	
        ,input  [31:0]                                                  desc_9_wuser_4_reg	
        ,input  [31:0]                                                  desc_9_wuser_5_reg	
        ,input  [31:0]                                                  desc_9_wuser_6_reg	
        ,input  [31:0]                                                  desc_9_wuser_7_reg	
        ,input  [31:0]                                                  desc_9_wuser_8_reg	
        ,input  [31:0]                                                  desc_9_wuser_9_reg	
        ,input  [31:0]                                                  desc_9_wuser_10_reg	
        ,input  [31:0]                                                  desc_9_wuser_11_reg	
        ,input  [31:0]                                                  desc_9_wuser_12_reg	
        ,input  [31:0]                                                  desc_9_wuser_13_reg	
        ,input  [31:0]                                                  desc_9_wuser_14_reg	
        ,input  [31:0]                                                  desc_9_wuser_15_reg	
        ,input  [31:0]                                                  desc_10_txn_type_reg			
        ,input  [31:0]                                                  desc_10_size_reg			
        ,input  [31:0]                                                  desc_10_data_offset_reg			
        ,input  [31:0]                                                  desc_10_data_host_addr_0_reg			
        ,input  [31:0]                                                  desc_10_data_host_addr_1_reg			
        ,input  [31:0]                                                  desc_10_data_host_addr_2_reg			
        ,input  [31:0]                                                  desc_10_data_host_addr_3_reg			
        ,input  [31:0]                                                  desc_10_wstrb_host_addr_0_reg			
        ,input  [31:0]                                                  desc_10_wstrb_host_addr_1_reg			
        ,input  [31:0]                                                  desc_10_wstrb_host_addr_2_reg			
        ,input  [31:0]                                                  desc_10_wstrb_host_addr_3_reg			
        ,input  [31:0]                                                  desc_10_axsize_reg			
        ,input  [31:0]                                                  desc_10_attr_reg			
        ,input  [31:0]                                                  desc_10_axaddr_0_reg			
        ,input  [31:0]                                                  desc_10_axaddr_1_reg			
        ,input  [31:0]                                                  desc_10_axaddr_2_reg			
        ,input  [31:0]                                                  desc_10_axaddr_3_reg			
        ,input  [31:0]                                                  desc_10_axid_0_reg			
        ,input  [31:0]                                                  desc_10_axid_1_reg			
        ,input  [31:0]                                                  desc_10_axid_2_reg			
        ,input  [31:0]                                                  desc_10_axid_3_reg			
        ,input  [31:0]                                                  desc_10_axuser_0_reg			
        ,input  [31:0]                                                  desc_10_axuser_1_reg			
        ,input  [31:0]                                                  desc_10_axuser_2_reg			
        ,input  [31:0]                                                  desc_10_axuser_3_reg			
        ,input  [31:0]                                                  desc_10_axuser_4_reg			
        ,input  [31:0]                                                  desc_10_axuser_5_reg			
        ,input  [31:0]                                                  desc_10_axuser_6_reg			
        ,input  [31:0]                                                  desc_10_axuser_7_reg			
        ,input  [31:0]                                                  desc_10_axuser_8_reg			
        ,input  [31:0]                                                  desc_10_axuser_9_reg			
        ,input  [31:0]                                                  desc_10_axuser_10_reg			
        ,input  [31:0]                                                  desc_10_axuser_11_reg			
        ,input  [31:0]                                                  desc_10_axuser_12_reg			
        ,input  [31:0]                                                  desc_10_axuser_13_reg			
        ,input  [31:0]                                                  desc_10_axuser_14_reg			
        ,input  [31:0]                                                  desc_10_axuser_15_reg			
        ,input  [31:0]                                                  desc_10_xuser_0_reg			
        ,input  [31:0]                                                  desc_10_xuser_1_reg			
        ,input  [31:0]                                                  desc_10_xuser_2_reg			
        ,input  [31:0]                                                  desc_10_xuser_3_reg			
        ,input  [31:0]                                                  desc_10_xuser_4_reg			
        ,input  [31:0]                                                  desc_10_xuser_5_reg			
        ,input  [31:0]                                                  desc_10_xuser_6_reg			
        ,input  [31:0]                                                  desc_10_xuser_7_reg			
        ,input  [31:0]                                                  desc_10_xuser_8_reg			
        ,input  [31:0]                                                  desc_10_xuser_9_reg			
        ,input  [31:0]                                                  desc_10_xuser_10_reg			
        ,input  [31:0]                                                  desc_10_xuser_11_reg			
        ,input  [31:0]                                                  desc_10_xuser_12_reg			
        ,input  [31:0]                                                  desc_10_xuser_13_reg			
        ,input  [31:0]                                                  desc_10_xuser_14_reg			
        ,input  [31:0]                                                  desc_10_xuser_15_reg			
        ,input  [31:0]                                                  desc_10_wuser_0_reg			
        ,input  [31:0]                                                  desc_10_wuser_1_reg			
        ,input  [31:0]                                                  desc_10_wuser_2_reg			
        ,input  [31:0]                                                  desc_10_wuser_3_reg			
        ,input  [31:0]                                                  desc_10_wuser_4_reg			
        ,input  [31:0]                                                  desc_10_wuser_5_reg			
        ,input  [31:0]                                                  desc_10_wuser_6_reg			
        ,input  [31:0]                                                  desc_10_wuser_7_reg			
        ,input  [31:0]                                                  desc_10_wuser_8_reg			
        ,input  [31:0]                                                  desc_10_wuser_9_reg			
        ,input  [31:0]                                                  desc_10_wuser_10_reg			
        ,input  [31:0]                                                  desc_10_wuser_11_reg			
        ,input  [31:0]                                                  desc_10_wuser_12_reg			
        ,input  [31:0]                                                  desc_10_wuser_13_reg			
        ,input  [31:0]                                                  desc_10_wuser_14_reg			
        ,input  [31:0]                                                  desc_10_wuser_15_reg			
        ,input  [31:0]                                                  desc_11_txn_type_reg			
        ,input  [31:0]                                                  desc_11_size_reg			
        ,input  [31:0]                                                  desc_11_data_offset_reg			
        ,input  [31:0]                                                  desc_11_data_host_addr_0_reg			
        ,input  [31:0]                                                  desc_11_data_host_addr_1_reg			
        ,input  [31:0]                                                  desc_11_data_host_addr_2_reg			
        ,input  [31:0]                                                  desc_11_data_host_addr_3_reg			
        ,input  [31:0]                                                  desc_11_wstrb_host_addr_0_reg			
        ,input  [31:0]                                                  desc_11_wstrb_host_addr_1_reg			
        ,input  [31:0]                                                  desc_11_wstrb_host_addr_2_reg			
        ,input  [31:0]                                                  desc_11_wstrb_host_addr_3_reg			
        ,input  [31:0]                                                  desc_11_axsize_reg			
        ,input  [31:0]                                                  desc_11_attr_reg			
        ,input  [31:0]                                                  desc_11_axaddr_0_reg			
        ,input  [31:0]                                                  desc_11_axaddr_1_reg			
        ,input  [31:0]                                                  desc_11_axaddr_2_reg			
        ,input  [31:0]                                                  desc_11_axaddr_3_reg			
        ,input  [31:0]                                                  desc_11_axid_0_reg			
        ,input  [31:0]                                                  desc_11_axid_1_reg			
        ,input  [31:0]                                                  desc_11_axid_2_reg			
        ,input  [31:0]                                                  desc_11_axid_3_reg			
        ,input  [31:0]                                                  desc_11_axuser_0_reg			
        ,input  [31:0]                                                  desc_11_axuser_1_reg			
        ,input  [31:0]                                                  desc_11_axuser_2_reg			
        ,input  [31:0]                                                  desc_11_axuser_3_reg			
        ,input  [31:0]                                                  desc_11_axuser_4_reg			
        ,input  [31:0]                                                  desc_11_axuser_5_reg			
        ,input  [31:0]                                                  desc_11_axuser_6_reg			
        ,input  [31:0]                                                  desc_11_axuser_7_reg			
        ,input  [31:0]                                                  desc_11_axuser_8_reg			
        ,input  [31:0]                                                  desc_11_axuser_9_reg			
        ,input  [31:0]                                                  desc_11_axuser_10_reg			
        ,input  [31:0]                                                  desc_11_axuser_11_reg			
        ,input  [31:0]                                                  desc_11_axuser_12_reg			
        ,input  [31:0]                                                  desc_11_axuser_13_reg			
        ,input  [31:0]                                                  desc_11_axuser_14_reg			
        ,input  [31:0]                                                  desc_11_axuser_15_reg			
        ,input  [31:0]                                                  desc_11_xuser_0_reg			
        ,input  [31:0]                                                  desc_11_xuser_1_reg			
        ,input  [31:0]                                                  desc_11_xuser_2_reg			
        ,input  [31:0]                                                  desc_11_xuser_3_reg			
        ,input  [31:0]                                                  desc_11_xuser_4_reg			
        ,input  [31:0]                                                  desc_11_xuser_5_reg			
        ,input  [31:0]                                                  desc_11_xuser_6_reg			
        ,input  [31:0]                                                  desc_11_xuser_7_reg			
        ,input  [31:0]                                                  desc_11_xuser_8_reg			
        ,input  [31:0]                                                  desc_11_xuser_9_reg			
        ,input  [31:0]                                                  desc_11_xuser_10_reg			
        ,input  [31:0]                                                  desc_11_xuser_11_reg			
        ,input  [31:0]                                                  desc_11_xuser_12_reg			
        ,input  [31:0]                                                  desc_11_xuser_13_reg			
        ,input  [31:0]                                                  desc_11_xuser_14_reg			
        ,input  [31:0]                                                  desc_11_xuser_15_reg			
        ,input  [31:0]                                                  desc_11_wuser_0_reg			
        ,input  [31:0]                                                  desc_11_wuser_1_reg			
        ,input  [31:0]                                                  desc_11_wuser_2_reg			
        ,input  [31:0]                                                  desc_11_wuser_3_reg			
        ,input  [31:0]                                                  desc_11_wuser_4_reg			
        ,input  [31:0]                                                  desc_11_wuser_5_reg			
        ,input  [31:0]                                                  desc_11_wuser_6_reg			
        ,input  [31:0]                                                  desc_11_wuser_7_reg			
        ,input  [31:0]                                                  desc_11_wuser_8_reg			
        ,input  [31:0]                                                  desc_11_wuser_9_reg			
        ,input  [31:0]                                                  desc_11_wuser_10_reg			
        ,input  [31:0]                                                  desc_11_wuser_11_reg			
        ,input  [31:0]                                                  desc_11_wuser_12_reg			
        ,input  [31:0]                                                  desc_11_wuser_13_reg			
        ,input  [31:0]                                                  desc_11_wuser_14_reg			
        ,input  [31:0]                                                  desc_11_wuser_15_reg			
        ,input  [31:0]                                                  desc_12_txn_type_reg			
        ,input  [31:0]                                                  desc_12_size_reg			
        ,input  [31:0]                                                  desc_12_data_offset_reg			
        ,input  [31:0]                                                  desc_12_data_host_addr_0_reg			
        ,input  [31:0]                                                  desc_12_data_host_addr_1_reg			
        ,input  [31:0]                                                  desc_12_data_host_addr_2_reg			
        ,input  [31:0]                                                  desc_12_data_host_addr_3_reg			
        ,input  [31:0]                                                  desc_12_wstrb_host_addr_0_reg			
        ,input  [31:0]                                                  desc_12_wstrb_host_addr_1_reg			
        ,input  [31:0]                                                  desc_12_wstrb_host_addr_2_reg			
        ,input  [31:0]                                                  desc_12_wstrb_host_addr_3_reg			
        ,input  [31:0]                                                  desc_12_axsize_reg			
        ,input  [31:0]                                                  desc_12_attr_reg			
        ,input  [31:0]                                                  desc_12_axaddr_0_reg			
        ,input  [31:0]                                                  desc_12_axaddr_1_reg			
        ,input  [31:0]                                                  desc_12_axaddr_2_reg			
        ,input  [31:0]                                                  desc_12_axaddr_3_reg			
        ,input  [31:0]                                                  desc_12_axid_0_reg			
        ,input  [31:0]                                                  desc_12_axid_1_reg			
        ,input  [31:0]                                                  desc_12_axid_2_reg			
        ,input  [31:0]                                                  desc_12_axid_3_reg			
        ,input  [31:0]                                                  desc_12_axuser_0_reg			
        ,input  [31:0]                                                  desc_12_axuser_1_reg			
        ,input  [31:0]                                                  desc_12_axuser_2_reg			
        ,input  [31:0]                                                  desc_12_axuser_3_reg			
        ,input  [31:0]                                                  desc_12_axuser_4_reg			
        ,input  [31:0]                                                  desc_12_axuser_5_reg			
        ,input  [31:0]                                                  desc_12_axuser_6_reg			
        ,input  [31:0]                                                  desc_12_axuser_7_reg			
        ,input  [31:0]                                                  desc_12_axuser_8_reg			
        ,input  [31:0]                                                  desc_12_axuser_9_reg			
        ,input  [31:0]                                                  desc_12_axuser_10_reg			
        ,input  [31:0]                                                  desc_12_axuser_11_reg			
        ,input  [31:0]                                                  desc_12_axuser_12_reg			
        ,input  [31:0]                                                  desc_12_axuser_13_reg			
        ,input  [31:0]                                                  desc_12_axuser_14_reg			
        ,input  [31:0]                                                  desc_12_axuser_15_reg			
        ,input  [31:0]                                                  desc_12_xuser_0_reg			
        ,input  [31:0]                                                  desc_12_xuser_1_reg			
        ,input  [31:0]                                                  desc_12_xuser_2_reg			
        ,input  [31:0]                                                  desc_12_xuser_3_reg			
        ,input  [31:0]                                                  desc_12_xuser_4_reg			
        ,input  [31:0]                                                  desc_12_xuser_5_reg			
        ,input  [31:0]                                                  desc_12_xuser_6_reg			
        ,input  [31:0]                                                  desc_12_xuser_7_reg			
        ,input  [31:0]                                                  desc_12_xuser_8_reg			
        ,input  [31:0]                                                  desc_12_xuser_9_reg			
        ,input  [31:0]                                                  desc_12_xuser_10_reg			
        ,input  [31:0]                                                  desc_12_xuser_11_reg			
        ,input  [31:0]                                                  desc_12_xuser_12_reg			
        ,input  [31:0]                                                  desc_12_xuser_13_reg			
        ,input  [31:0]                                                  desc_12_xuser_14_reg			
        ,input  [31:0]                                                  desc_12_xuser_15_reg			
        ,input  [31:0]                                                  desc_12_wuser_0_reg			
        ,input  [31:0]                                                  desc_12_wuser_1_reg			
        ,input  [31:0]                                                  desc_12_wuser_2_reg			
        ,input  [31:0]                                                  desc_12_wuser_3_reg			
        ,input  [31:0]                                                  desc_12_wuser_4_reg			
        ,input  [31:0]                                                  desc_12_wuser_5_reg			
        ,input  [31:0]                                                  desc_12_wuser_6_reg			
        ,input  [31:0]                                                  desc_12_wuser_7_reg			
        ,input  [31:0]                                                  desc_12_wuser_8_reg			
        ,input  [31:0]                                                  desc_12_wuser_9_reg			
        ,input  [31:0]                                                  desc_12_wuser_10_reg			
        ,input  [31:0]                                                  desc_12_wuser_11_reg			
        ,input  [31:0]                                                  desc_12_wuser_12_reg			
        ,input  [31:0]                                                  desc_12_wuser_13_reg			
        ,input  [31:0]                                                  desc_12_wuser_14_reg			
        ,input  [31:0]                                                  desc_12_wuser_15_reg			
        ,input  [31:0]                                                  desc_13_txn_type_reg			
        ,input  [31:0]                                                  desc_13_size_reg			
        ,input  [31:0]                                                  desc_13_data_offset_reg			
        ,input  [31:0]                                                  desc_13_data_host_addr_0_reg			
        ,input  [31:0]                                                  desc_13_data_host_addr_1_reg			
        ,input  [31:0]                                                  desc_13_data_host_addr_2_reg			
        ,input  [31:0]                                                  desc_13_data_host_addr_3_reg			
        ,input  [31:0]                                                  desc_13_wstrb_host_addr_0_reg			
        ,input  [31:0]                                                  desc_13_wstrb_host_addr_1_reg			
        ,input  [31:0]                                                  desc_13_wstrb_host_addr_2_reg			
        ,input  [31:0]                                                  desc_13_wstrb_host_addr_3_reg			
        ,input  [31:0]                                                  desc_13_axsize_reg			
        ,input  [31:0]                                                  desc_13_attr_reg			
        ,input  [31:0]                                                  desc_13_axaddr_0_reg			
        ,input  [31:0]                                                  desc_13_axaddr_1_reg			
        ,input  [31:0]                                                  desc_13_axaddr_2_reg			
        ,input  [31:0]                                                  desc_13_axaddr_3_reg			
        ,input  [31:0]                                                  desc_13_axid_0_reg			
        ,input  [31:0]                                                  desc_13_axid_1_reg			
        ,input  [31:0]                                                  desc_13_axid_2_reg			
        ,input  [31:0]                                                  desc_13_axid_3_reg			
        ,input  [31:0]                                                  desc_13_axuser_0_reg			
        ,input  [31:0]                                                  desc_13_axuser_1_reg			
        ,input  [31:0]                                                  desc_13_axuser_2_reg			
        ,input  [31:0]                                                  desc_13_axuser_3_reg			
        ,input  [31:0]                                                  desc_13_axuser_4_reg			
        ,input  [31:0]                                                  desc_13_axuser_5_reg			
        ,input  [31:0]                                                  desc_13_axuser_6_reg			
        ,input  [31:0]                                                  desc_13_axuser_7_reg			
        ,input  [31:0]                                                  desc_13_axuser_8_reg			
        ,input  [31:0]                                                  desc_13_axuser_9_reg			
        ,input  [31:0]                                                  desc_13_axuser_10_reg			
        ,input  [31:0]                                                  desc_13_axuser_11_reg			
        ,input  [31:0]                                                  desc_13_axuser_12_reg			
        ,input  [31:0]                                                  desc_13_axuser_13_reg			
        ,input  [31:0]                                                  desc_13_axuser_14_reg			
        ,input  [31:0]                                                  desc_13_axuser_15_reg			
        ,input  [31:0]                                                  desc_13_xuser_0_reg			
        ,input  [31:0]                                                  desc_13_xuser_1_reg			
        ,input  [31:0]                                                  desc_13_xuser_2_reg			
        ,input  [31:0]                                                  desc_13_xuser_3_reg			
        ,input  [31:0]                                                  desc_13_xuser_4_reg			
        ,input  [31:0]                                                  desc_13_xuser_5_reg			
        ,input  [31:0]                                                  desc_13_xuser_6_reg			
        ,input  [31:0]                                                  desc_13_xuser_7_reg			
        ,input  [31:0]                                                  desc_13_xuser_8_reg			
        ,input  [31:0]                                                  desc_13_xuser_9_reg			
        ,input  [31:0]                                                  desc_13_xuser_10_reg			
        ,input  [31:0]                                                  desc_13_xuser_11_reg			
        ,input  [31:0]                                                  desc_13_xuser_12_reg			
        ,input  [31:0]                                                  desc_13_xuser_13_reg			
        ,input  [31:0]                                                  desc_13_xuser_14_reg			
        ,input  [31:0]                                                  desc_13_xuser_15_reg			
        ,input  [31:0]                                                  desc_13_wuser_0_reg			
        ,input  [31:0]                                                  desc_13_wuser_1_reg			
        ,input  [31:0]                                                  desc_13_wuser_2_reg			
        ,input  [31:0]                                                  desc_13_wuser_3_reg			
        ,input  [31:0]                                                  desc_13_wuser_4_reg			
        ,input  [31:0]                                                  desc_13_wuser_5_reg			
        ,input  [31:0]                                                  desc_13_wuser_6_reg			
        ,input  [31:0]                                                  desc_13_wuser_7_reg			
        ,input  [31:0]                                                  desc_13_wuser_8_reg			
        ,input  [31:0]                                                  desc_13_wuser_9_reg			
        ,input  [31:0]                                                  desc_13_wuser_10_reg			
        ,input  [31:0]                                                  desc_13_wuser_11_reg			
        ,input  [31:0]                                                  desc_13_wuser_12_reg			
        ,input  [31:0]                                                  desc_13_wuser_13_reg			
        ,input  [31:0]                                                  desc_13_wuser_14_reg			
        ,input  [31:0]                                                  desc_13_wuser_15_reg			
        ,input  [31:0]                                                  desc_14_txn_type_reg			
        ,input  [31:0]                                                  desc_14_size_reg			
        ,input  [31:0]                                                  desc_14_data_offset_reg			
        ,input  [31:0]                                                  desc_14_data_host_addr_0_reg			
        ,input  [31:0]                                                  desc_14_data_host_addr_1_reg			
        ,input  [31:0]                                                  desc_14_data_host_addr_2_reg			
        ,input  [31:0]                                                  desc_14_data_host_addr_3_reg			
        ,input  [31:0]                                                  desc_14_wstrb_host_addr_0_reg			
        ,input  [31:0]                                                  desc_14_wstrb_host_addr_1_reg			
        ,input  [31:0]                                                  desc_14_wstrb_host_addr_2_reg			
        ,input  [31:0]                                                  desc_14_wstrb_host_addr_3_reg			
        ,input  [31:0]                                                  desc_14_axsize_reg			
        ,input  [31:0]                                                  desc_14_attr_reg			
        ,input  [31:0]                                                  desc_14_axaddr_0_reg			
        ,input  [31:0]                                                  desc_14_axaddr_1_reg			
        ,input  [31:0]                                                  desc_14_axaddr_2_reg			
        ,input  [31:0]                                                  desc_14_axaddr_3_reg			
        ,input  [31:0]                                                  desc_14_axid_0_reg			
        ,input  [31:0]                                                  desc_14_axid_1_reg			
        ,input  [31:0]                                                  desc_14_axid_2_reg			
        ,input  [31:0]                                                  desc_14_axid_3_reg			
        ,input  [31:0]                                                  desc_14_axuser_0_reg			
        ,input  [31:0]                                                  desc_14_axuser_1_reg			
        ,input  [31:0]                                                  desc_14_axuser_2_reg			
        ,input  [31:0]                                                  desc_14_axuser_3_reg			
        ,input  [31:0]                                                  desc_14_axuser_4_reg			
        ,input  [31:0]                                                  desc_14_axuser_5_reg			
        ,input  [31:0]                                                  desc_14_axuser_6_reg			
        ,input  [31:0]                                                  desc_14_axuser_7_reg			
        ,input  [31:0]                                                  desc_14_axuser_8_reg			
        ,input  [31:0]                                                  desc_14_axuser_9_reg			
        ,input  [31:0]                                                  desc_14_axuser_10_reg			
        ,input  [31:0]                                                  desc_14_axuser_11_reg			
        ,input  [31:0]                                                  desc_14_axuser_12_reg			
        ,input  [31:0]                                                  desc_14_axuser_13_reg			
        ,input  [31:0]                                                  desc_14_axuser_14_reg			
        ,input  [31:0]                                                  desc_14_axuser_15_reg			
        ,input  [31:0]                                                  desc_14_xuser_0_reg			
        ,input  [31:0]                                                  desc_14_xuser_1_reg			
        ,input  [31:0]                                                  desc_14_xuser_2_reg			
        ,input  [31:0]                                                  desc_14_xuser_3_reg			
        ,input  [31:0]                                                  desc_14_xuser_4_reg			
        ,input  [31:0]                                                  desc_14_xuser_5_reg			
        ,input  [31:0]                                                  desc_14_xuser_6_reg			
        ,input  [31:0]                                                  desc_14_xuser_7_reg			
        ,input  [31:0]                                                  desc_14_xuser_8_reg			
        ,input  [31:0]                                                  desc_14_xuser_9_reg			
        ,input  [31:0]                                                  desc_14_xuser_10_reg			
        ,input  [31:0]                                                  desc_14_xuser_11_reg			
        ,input  [31:0]                                                  desc_14_xuser_12_reg			
        ,input  [31:0]                                                  desc_14_xuser_13_reg			
        ,input  [31:0]                                                  desc_14_xuser_14_reg			
        ,input  [31:0]                                                  desc_14_xuser_15_reg			
        ,input  [31:0]                                                  desc_14_wuser_0_reg			
        ,input  [31:0]                                                  desc_14_wuser_1_reg			
        ,input  [31:0]                                                  desc_14_wuser_2_reg			
        ,input  [31:0]                                                  desc_14_wuser_3_reg			
        ,input  [31:0]                                                  desc_14_wuser_4_reg			
        ,input  [31:0]                                                  desc_14_wuser_5_reg			
        ,input  [31:0]                                                  desc_14_wuser_6_reg			
        ,input  [31:0]                                                  desc_14_wuser_7_reg			
        ,input  [31:0]                                                  desc_14_wuser_8_reg			
        ,input  [31:0]                                                  desc_14_wuser_9_reg			
        ,input  [31:0]                                                  desc_14_wuser_10_reg			
        ,input  [31:0]                                                  desc_14_wuser_11_reg			
        ,input  [31:0]                                                  desc_14_wuser_12_reg			
        ,input  [31:0]                                                  desc_14_wuser_13_reg			
        ,input  [31:0]                                                  desc_14_wuser_14_reg			
        ,input  [31:0]                                                  desc_14_wuser_15_reg			
        ,input  [31:0]                                                  desc_15_txn_type_reg			
        ,input  [31:0]                                                  desc_15_size_reg			
        ,input  [31:0]                                                  desc_15_data_offset_reg			
        ,input  [31:0]                                                  desc_15_data_host_addr_0_reg			
        ,input  [31:0]                                                  desc_15_data_host_addr_1_reg			
        ,input  [31:0]                                                  desc_15_data_host_addr_2_reg			
        ,input  [31:0]                                                  desc_15_data_host_addr_3_reg			
        ,input  [31:0]                                                  desc_15_wstrb_host_addr_0_reg			
        ,input  [31:0]                                                  desc_15_wstrb_host_addr_1_reg			
        ,input  [31:0]                                                  desc_15_wstrb_host_addr_2_reg			
        ,input  [31:0]                                                  desc_15_wstrb_host_addr_3_reg			
        ,input  [31:0]                                                  desc_15_axsize_reg			
        ,input  [31:0]                                                  desc_15_attr_reg			
        ,input  [31:0]                                                  desc_15_axaddr_0_reg			
        ,input  [31:0]                                                  desc_15_axaddr_1_reg			
        ,input  [31:0]                                                  desc_15_axaddr_2_reg			
        ,input  [31:0]                                                  desc_15_axaddr_3_reg			
        ,input  [31:0]                                                  desc_15_axid_0_reg			
        ,input  [31:0]                                                  desc_15_axid_1_reg			
        ,input  [31:0]                                                  desc_15_axid_2_reg			
        ,input  [31:0]                                                  desc_15_axid_3_reg			
        ,input  [31:0]                                                  desc_15_axuser_0_reg			
        ,input  [31:0]                                                  desc_15_axuser_1_reg			
        ,input  [31:0]                                                  desc_15_axuser_2_reg			
        ,input  [31:0]                                                  desc_15_axuser_3_reg			
        ,input  [31:0]                                                  desc_15_axuser_4_reg			
        ,input  [31:0]                                                  desc_15_axuser_5_reg			
        ,input  [31:0]                                                  desc_15_axuser_6_reg			
        ,input  [31:0]                                                  desc_15_axuser_7_reg			
        ,input  [31:0]                                                  desc_15_axuser_8_reg			
        ,input  [31:0]                                                  desc_15_axuser_9_reg			
        ,input  [31:0]                                                  desc_15_axuser_10_reg			
        ,input  [31:0]                                                  desc_15_axuser_11_reg			
        ,input  [31:0]                                                  desc_15_axuser_12_reg			
        ,input  [31:0]                                                  desc_15_axuser_13_reg			
        ,input  [31:0]                                                  desc_15_axuser_14_reg			
        ,input  [31:0]                                                  desc_15_axuser_15_reg			
        ,input  [31:0]                                                  desc_15_xuser_0_reg			
        ,input  [31:0]                                                  desc_15_xuser_1_reg			
        ,input  [31:0]                                                  desc_15_xuser_2_reg			
        ,input  [31:0]                                                  desc_15_xuser_3_reg			
        ,input  [31:0]                                                  desc_15_xuser_4_reg			
        ,input  [31:0]                                                  desc_15_xuser_5_reg			
        ,input  [31:0]                                                  desc_15_xuser_6_reg			
        ,input  [31:0]                                                  desc_15_xuser_7_reg			
        ,input  [31:0]                                                  desc_15_xuser_8_reg			
        ,input  [31:0]                                                  desc_15_xuser_9_reg			
        ,input  [31:0]                                                  desc_15_xuser_10_reg			
        ,input  [31:0]                                                  desc_15_xuser_11_reg			
        ,input  [31:0]                                                  desc_15_xuser_12_reg			
        ,input  [31:0]                                                  desc_15_xuser_13_reg			
        ,input  [31:0]                                                  desc_15_xuser_14_reg			
        ,input  [31:0]                                                  desc_15_xuser_15_reg			
        ,input  [31:0]                                                  desc_15_wuser_0_reg			
        ,input  [31:0]                                                  desc_15_wuser_1_reg			
        ,input  [31:0]                                                  desc_15_wuser_2_reg			
        ,input  [31:0]                                                  desc_15_wuser_3_reg			
        ,input  [31:0]                                                  desc_15_wuser_4_reg			
        ,input  [31:0]                                                  desc_15_wuser_5_reg			
        ,input  [31:0]                                                  desc_15_wuser_6_reg			
        ,input  [31:0]                                                  desc_15_wuser_7_reg			
        ,input  [31:0]                                                  desc_15_wuser_8_reg			
        ,input  [31:0]                                                  desc_15_wuser_9_reg			
        ,input  [31:0]                                                  desc_15_wuser_10_reg			
        ,input  [31:0]                                                  desc_15_wuser_11_reg			
        ,input  [31:0]                                                  desc_15_wuser_12_reg			
        ,input  [31:0]                                                  desc_15_wuser_13_reg			
        ,input  [31:0]                                                  desc_15_wuser_14_reg			
        ,input  [31:0]                                                  desc_15_wuser_15_reg
        			
        ,output [31:0]                                                  uc2rb_intr_error_status_reg				
        ,output [31:0]                                                  uc2rb_ownership_reg				
        ,output [31:0]                                                  uc2rb_intr_txn_avail_status_reg				
        ,output [31:0]                                                  uc2rb_intr_comp_status_reg				
        ,output [31:0]                                                  uc2rb_status_busy_reg				
        ,output [31:0]                                                  uc2rb_resp_fifo_free_level_reg				
        ,output [31:0]                                                  uc2rb_desc_0_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_0_size_reg				
        ,output [31:0]                                                  uc2rb_desc_0_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_0_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_1_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_1_size_reg				
        ,output [31:0]                                                  uc2rb_desc_1_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_1_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_2_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_2_size_reg				
        ,output [31:0]                                                  uc2rb_desc_2_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_2_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_3_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_3_size_reg				
        ,output [31:0]                                                  uc2rb_desc_3_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_3_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_4_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_4_size_reg				
        ,output [31:0]                                                  uc2rb_desc_4_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_4_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_5_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_5_size_reg				
        ,output [31:0]                                                  uc2rb_desc_5_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_5_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_6_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_6_size_reg				
        ,output [31:0]                                                  uc2rb_desc_6_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_6_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_7_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_7_size_reg				
        ,output [31:0]                                                  uc2rb_desc_7_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_7_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_8_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_8_size_reg				
        ,output [31:0]                                                  uc2rb_desc_8_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_8_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_9_txn_type_reg				
        ,output [31:0]                                                  uc2rb_desc_9_size_reg				
        ,output [31:0]                                                  uc2rb_desc_9_data_offset_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axsize_reg				
        ,output [31:0]                                                  uc2rb_desc_9_attr_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_0_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_1_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_2_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_3_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axid_0_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axid_1_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axid_2_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axid_3_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_0_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_1_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_2_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_3_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_4_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_5_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_6_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_7_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_8_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_9_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_10_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_11_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_12_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_13_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_14_reg				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_15_reg				
        ,output [31:0]                                                  uc2rb_desc_10_txn_type_reg						
        ,output [31:0]                                                  uc2rb_desc_10_size_reg						
        ,output [31:0]                                                  uc2rb_desc_10_data_offset_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axsize_reg						
        ,output [31:0]                                                  uc2rb_desc_10_attr_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_0_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_1_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_2_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_3_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axid_0_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axid_1_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axid_2_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axid_3_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_11_txn_type_reg						
        ,output [31:0]                                                  uc2rb_desc_11_size_reg						
        ,output [31:0]                                                  uc2rb_desc_11_data_offset_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axsize_reg						
        ,output [31:0]                                                  uc2rb_desc_11_attr_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_0_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_1_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_2_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_3_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axid_0_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axid_1_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axid_2_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axid_3_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_12_txn_type_reg						
        ,output [31:0]                                                  uc2rb_desc_12_size_reg						
        ,output [31:0]                                                  uc2rb_desc_12_data_offset_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axsize_reg						
        ,output [31:0]                                                  uc2rb_desc_12_attr_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_0_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_1_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_2_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_3_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axid_0_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axid_1_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axid_2_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axid_3_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_13_txn_type_reg						
        ,output [31:0]                                                  uc2rb_desc_13_size_reg						
        ,output [31:0]                                                  uc2rb_desc_13_data_offset_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axsize_reg						
        ,output [31:0]                                                  uc2rb_desc_13_attr_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_0_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_1_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_2_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_3_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axid_0_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axid_1_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axid_2_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axid_3_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_14_txn_type_reg						
        ,output [31:0]                                                  uc2rb_desc_14_size_reg						
        ,output [31:0]                                                  uc2rb_desc_14_data_offset_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axsize_reg						
        ,output [31:0]                                                  uc2rb_desc_14_attr_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_0_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_1_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_2_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_3_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axid_0_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axid_1_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axid_2_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axid_3_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_15_txn_type_reg						
        ,output [31:0]                                                  uc2rb_desc_15_size_reg						
        ,output [31:0]                                                  uc2rb_desc_15_data_offset_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axsize_reg						
        ,output [31:0]                                                  uc2rb_desc_15_attr_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_0_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_1_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_2_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_3_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axid_0_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axid_1_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axid_2_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axid_3_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_15_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_0_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_1_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_2_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_3_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_4_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_5_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_6_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_7_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_8_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_9_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_10_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_11_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_12_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_13_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_14_reg						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_15_reg						
        
        ,output [31:0]                                                  uc2rb_intr_error_status_reg_we				
        ,output [31:0]                                                  uc2rb_ownership_reg_we				
        ,output [31:0]                                                  uc2rb_intr_txn_avail_status_reg_we				
        ,output [31:0]                                                  uc2rb_intr_comp_status_reg_we				
        ,output [31:0]                                                  uc2rb_status_busy_reg_we				
        ,output [31:0]                                                  uc2rb_resp_fifo_free_level_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_0_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_1_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_2_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_3_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_4_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_5_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_6_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_7_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_8_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_txn_type_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_size_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_data_offset_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axsize_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_attr_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axaddr_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axid_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axid_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axid_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axid_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_axuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_0_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_1_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_2_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_3_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_4_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_5_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_6_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_7_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_8_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_9_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_10_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_11_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_12_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_13_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_14_reg_we				
        ,output [31:0]                                                  uc2rb_desc_9_wuser_15_reg_we				
        ,output [31:0]                                                  uc2rb_desc_10_txn_type_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_size_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_data_offset_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axsize_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_attr_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axaddr_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axid_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axid_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axid_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axid_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_axuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_10_wuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_txn_type_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_size_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_data_offset_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axsize_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_attr_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axaddr_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axid_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axid_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axid_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axid_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_axuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_11_wuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_txn_type_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_size_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_data_offset_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axsize_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_attr_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axaddr_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axid_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axid_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axid_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axid_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_axuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_12_wuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_txn_type_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_size_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_data_offset_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axsize_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_attr_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axaddr_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axid_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axid_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axid_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axid_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_axuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_13_wuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_txn_type_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_size_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_data_offset_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axsize_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_attr_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axaddr_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axid_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axid_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axid_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axid_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_axuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_14_wuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_txn_type_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_size_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_data_offset_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axsize_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_attr_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axaddr_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axid_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axid_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axid_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axid_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_axuser_15_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_0_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_1_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_2_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_3_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_4_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_5_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_6_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_7_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_8_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_9_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_10_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_11_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_12_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_13_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_14_reg_we						
        ,output [31:0]                                                  uc2rb_desc_15_wuser_15_reg_we						

        //RDATA_RAM signals
        ,output	[(`CLOG2((RAM_SIZE*8)/DATA_WIDTH))-1:0]                 uc2rb_rd_addr		
        ,input 	[DATA_WIDTH-1:0]                                        rb2uc_rd_data
        
        //WDATA_RAM and WSTRB_RAM signals				
        ,output	     	                                                uc2rb_wr_we		
        ,output	[(DATA_WIDTH/8)-1:0]                                    uc2rb_wr_bwe            //Generate all 1s always 	
        ,output	[(`CLOG2((RAM_SIZE*8)/DATA_WIDTH))-1:0]                 uc2rb_wr_addr		
        ,output	[DATA_WIDTH-1:0]                                        uc2rb_wr_data   		
        ,output	[(DATA_WIDTH/8)-1:0]                                    uc2rb_wr_wstrb   		
              		                                                	
        ,output	[MAX_DESC-1:0]                                          uc2hm_trig
        ,input 	[MAX_DESC-1:0]                                          hm2uc_done

  );
   
localparam DESC_IDX_WIDTH                                               = `CLOG2(MAX_DESC);
localparam RAM_OFFSET_WIDTH                                             = `CLOG2((RAM_SIZE*8)/DATA_WIDTH);

//Declare all fields ( <reg>_<field>_f )
wire	[7:0]				version_major_ver_f;
wire	[7:0]				version_minor_ver_f;
wire	[7:0]				bridge_type_type_f;
wire	[7:0]				axi_bridge_config_user_width_f;
wire	[7:0]				axi_bridge_config_id_width_f;
wire	[2:0]				axi_bridge_config_data_width_f;
wire	     				reset_dut_srst_3_f;
wire	     				reset_dut_srst_2_f;
wire	     				reset_dut_srst_1_f;
wire	     				reset_dut_srst_0_f;
wire	     				reset_srst_f;
wire	     				mode_select_imm_bresp_f;
wire	     				mode_select_mode_2_f;
wire	     				mode_select_mode_0_1_f;
wire	[MAX_DESC-1:0]			ownership_own_f;
wire	[MAX_DESC-1:0]			ownership_flip_flip_f;
wire	[MAX_DESC-1:0]			status_resp_comp_resp_comp_f;
wire	[31:0]				status_resp_resp_f;
wire	[MAX_DESC-1:0]			status_busy_busy_f;
wire	[DESC_IDX_WIDTH:0]              resp_fifo_free_level_level_f;
wire	     				intr_status_comp_f;
wire	     				intr_status_c2h_f;
wire	     				intr_status_error_f;
wire	     				intr_status_txn_avail_f;
wire	[MAX_DESC-1:0]			intr_txn_avail_status_avail_f;
wire	[MAX_DESC-1:0]			intr_txn_avail_clear_clr_avail_f;
wire	[MAX_DESC-1:0]			intr_txn_avail_enable_en_avail_f;
wire	[MAX_DESC-1:0]			intr_comp_status_comp_f;
wire	[MAX_DESC-1:0]			intr_comp_clear_clr_comp_f;
wire	[MAX_DESC-1:0]			intr_comp_enable_en_comp_f;
wire	     				intr_error_status_err_2_f;
wire	     				intr_error_status_err_1_f;
wire	     				intr_error_status_err_0_f;
wire	     				intr_error_clear_clr_err_2_f;
wire	     				intr_error_clear_clr_err_1_f;
wire	     				intr_error_clear_clr_err_0_f;
wire	     				intr_error_enable_en_err_2_f;
wire	     				intr_error_enable_en_err_1_f;
wire	     				intr_error_enable_en_err_0_f;
wire	[31:0]				intr_h2c_0_h2c_f;
wire	[31:0]				intr_h2c_1_h2c_f;
wire	[31:0]				intr_c2h_0_status_c2h_f;
wire	[31:0]				intr_c2h_1_status_c2h_f;
wire	[31:0]				c2h_gpio_0_status_gpio_f;
wire	[31:0]				c2h_gpio_1_status_gpio_f;
wire	[31:0]				c2h_gpio_2_status_gpio_f;
wire	[31:0]				c2h_gpio_3_status_gpio_f;
wire	[31:0]				c2h_gpio_4_status_gpio_f;
wire	[31:0]				c2h_gpio_5_status_gpio_f;
wire	[31:0]				c2h_gpio_6_status_gpio_f;
wire	[31:0]				c2h_gpio_7_status_gpio_f;
wire	[31:0]				c2h_gpio_8_status_gpio_f;
wire	[31:0]				c2h_gpio_9_status_gpio_f;
wire	[31:0]				c2h_gpio_10_status_gpio_f;
wire	[31:0]				c2h_gpio_11_status_gpio_f;
wire	[31:0]				c2h_gpio_12_status_gpio_f;
wire	[31:0]				c2h_gpio_13_status_gpio_f;
wire	[31:0]				c2h_gpio_14_status_gpio_f;
wire	[31:0]				c2h_gpio_15_status_gpio_f;
wire	[31:0]				addr_in_0_addr_f;
wire	[31:0]				addr_in_1_addr_f;
wire	[31:0]				addr_in_2_addr_f;
wire	[31:0]				addr_in_3_addr_f;
wire	[31:0]				trans_mask_0_addr_f;
wire	[31:0]				trans_mask_1_addr_f;
wire	[31:0]				trans_mask_2_addr_f;
wire	[31:0]				trans_mask_3_addr_f;
wire	[31:0]				trans_addr_0_addr_f;
wire	[31:0]				trans_addr_1_addr_f;
wire	[31:0]				trans_addr_2_addr_f;
wire	[31:0]				trans_addr_3_addr_f;
wire    [31:0]                          resp_order_field_f;

wire [0:0]	desc_0_txn_type_wr_strb_f;
wire [0:0]	desc_0_txn_type_wr_rd_f;
wire [3:0]	desc_0_attr_axregion_f;
wire [3:0]	desc_0_attr_axqos_f;
wire [2:0]	desc_0_attr_axprot_f;
wire [3:0]	desc_0_attr_axcache_f;
wire [1:0]	desc_0_attr_axlock_f;
wire [1:0]	desc_0_attr_axburst_f;
wire [31:0]	desc_0_axid_0_axid_f;
wire [31:0]	desc_0_axid_1_axid_f;
wire [31:0]	desc_0_axid_2_axid_f;
wire [31:0]	desc_0_axid_3_axid_f;
wire [31:0]	desc_0_axuser_0_axuser_f;
wire [31:0]	desc_0_axuser_1_axuser_f;
wire [31:0]	desc_0_axuser_2_axuser_f;
wire [31:0]	desc_0_axuser_3_axuser_f;
wire [31:0]	desc_0_axuser_4_axuser_f;
wire [31:0]	desc_0_axuser_5_axuser_f;
wire [31:0]	desc_0_axuser_6_axuser_f;
wire [31:0]	desc_0_axuser_7_axuser_f;
wire [31:0]	desc_0_axuser_8_axuser_f;
wire [31:0]	desc_0_axuser_9_axuser_f;
wire [31:0]	desc_0_axuser_10_axuser_f;
wire [31:0]	desc_0_axuser_11_axuser_f;
wire [31:0]	desc_0_axuser_12_axuser_f;
wire [31:0]	desc_0_axuser_13_axuser_f;
wire [31:0]	desc_0_axuser_14_axuser_f;
wire [31:0]	desc_0_axuser_15_axuser_f;
wire [15:0]	desc_0_size_txn_size_f;
wire [2:0]	desc_0_axsize_axsize_f;
wire [31:0]	desc_0_axaddr_0_addr_f;
wire [31:0]	desc_0_axaddr_1_addr_f;
wire [31:0]	desc_0_axaddr_2_addr_f;
wire [31:0]	desc_0_axaddr_3_addr_f;
wire [31:0]	desc_0_data_offset_addr_f;
wire [31:0]	desc_0_wuser_0_wuser_f;
wire [31:0]	desc_0_wuser_1_wuser_f;
wire [31:0]	desc_0_wuser_2_wuser_f;
wire [31:0]	desc_0_wuser_3_wuser_f;
wire [31:0]	desc_0_wuser_4_wuser_f;
wire [31:0]	desc_0_wuser_5_wuser_f;
wire [31:0]	desc_0_wuser_6_wuser_f;
wire [31:0]	desc_0_wuser_7_wuser_f;
wire [31:0]	desc_0_wuser_8_wuser_f;
wire [31:0]	desc_0_wuser_9_wuser_f;
wire [31:0]	desc_0_wuser_10_wuser_f;
wire [31:0]	desc_0_wuser_11_wuser_f;
wire [31:0]	desc_0_wuser_12_wuser_f;
wire [31:0]	desc_0_wuser_13_wuser_f;
wire [31:0]	desc_0_wuser_14_wuser_f;
wire [31:0]	desc_0_wuser_15_wuser_f;
wire [31:0]	desc_0_data_host_addr_0_addr_f;
wire [31:0]	desc_0_data_host_addr_1_addr_f;
wire [31:0]	desc_0_data_host_addr_2_addr_f;
wire [31:0]	desc_0_data_host_addr_3_addr_f;
wire [31:0]	desc_0_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_0_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_0_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_0_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_0_xuser_0_xuser_f;
wire [31:0]	desc_0_xuser_1_xuser_f;
wire [31:0]	desc_0_xuser_2_xuser_f;
wire [31:0]	desc_0_xuser_3_xuser_f;
wire [31:0]	desc_0_xuser_4_xuser_f;
wire [31:0]	desc_0_xuser_5_xuser_f;
wire [31:0]	desc_0_xuser_6_xuser_f;
wire [31:0]	desc_0_xuser_7_xuser_f;
wire [31:0]	desc_0_xuser_8_xuser_f;
wire [31:0]	desc_0_xuser_9_xuser_f;
wire [31:0]	desc_0_xuser_10_xuser_f;
wire [31:0]	desc_0_xuser_11_xuser_f;
wire [31:0]	desc_0_xuser_12_xuser_f;
wire [31:0]	desc_0_xuser_13_xuser_f;
wire [31:0]	desc_0_xuser_14_xuser_f;
wire [31:0]	desc_0_xuser_15_xuser_f;
wire [0:0]	desc_1_txn_type_wr_strb_f;
wire [0:0]	desc_1_txn_type_wr_rd_f;
wire [3:0]	desc_1_attr_axregion_f;
wire [3:0]	desc_1_attr_axqos_f;
wire [2:0]	desc_1_attr_axprot_f;
wire [3:0]	desc_1_attr_axcache_f;
wire [1:0]	desc_1_attr_axlock_f;
wire [1:0]	desc_1_attr_axburst_f;
wire [31:0]	desc_1_axid_0_axid_f;
wire [31:0]	desc_1_axid_1_axid_f;
wire [31:0]	desc_1_axid_2_axid_f;
wire [31:0]	desc_1_axid_3_axid_f;
wire [31:0]	desc_1_axuser_0_axuser_f;
wire [31:0]	desc_1_axuser_1_axuser_f;
wire [31:0]	desc_1_axuser_2_axuser_f;
wire [31:0]	desc_1_axuser_3_axuser_f;
wire [31:0]	desc_1_axuser_4_axuser_f;
wire [31:0]	desc_1_axuser_5_axuser_f;
wire [31:0]	desc_1_axuser_6_axuser_f;
wire [31:0]	desc_1_axuser_7_axuser_f;
wire [31:0]	desc_1_axuser_8_axuser_f;
wire [31:0]	desc_1_axuser_9_axuser_f;
wire [31:0]	desc_1_axuser_10_axuser_f;
wire [31:0]	desc_1_axuser_11_axuser_f;
wire [31:0]	desc_1_axuser_12_axuser_f;
wire [31:0]	desc_1_axuser_13_axuser_f;
wire [31:0]	desc_1_axuser_14_axuser_f;
wire [31:0]	desc_1_axuser_15_axuser_f;
wire [15:0]	desc_1_size_txn_size_f;
wire [2:0]	desc_1_axsize_axsize_f;
wire [31:0]	desc_1_axaddr_0_addr_f;
wire [31:0]	desc_1_axaddr_1_addr_f;
wire [31:0]	desc_1_axaddr_2_addr_f;
wire [31:0]	desc_1_axaddr_3_addr_f;
wire [31:0]	desc_1_data_offset_addr_f;
wire [31:0]	desc_1_wuser_0_wuser_f;
wire [31:0]	desc_1_wuser_1_wuser_f;
wire [31:0]	desc_1_wuser_2_wuser_f;
wire [31:0]	desc_1_wuser_3_wuser_f;
wire [31:0]	desc_1_wuser_4_wuser_f;
wire [31:0]	desc_1_wuser_5_wuser_f;
wire [31:0]	desc_1_wuser_6_wuser_f;
wire [31:0]	desc_1_wuser_7_wuser_f;
wire [31:0]	desc_1_wuser_8_wuser_f;
wire [31:0]	desc_1_wuser_9_wuser_f;
wire [31:0]	desc_1_wuser_10_wuser_f;
wire [31:0]	desc_1_wuser_11_wuser_f;
wire [31:0]	desc_1_wuser_12_wuser_f;
wire [31:0]	desc_1_wuser_13_wuser_f;
wire [31:0]	desc_1_wuser_14_wuser_f;
wire [31:0]	desc_1_wuser_15_wuser_f;
wire [31:0]	desc_1_data_host_addr_0_addr_f;
wire [31:0]	desc_1_data_host_addr_1_addr_f;
wire [31:0]	desc_1_data_host_addr_2_addr_f;
wire [31:0]	desc_1_data_host_addr_3_addr_f;
wire [31:0]	desc_1_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_1_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_1_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_1_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_1_xuser_0_xuser_f;
wire [31:0]	desc_1_xuser_1_xuser_f;
wire [31:0]	desc_1_xuser_2_xuser_f;
wire [31:0]	desc_1_xuser_3_xuser_f;
wire [31:0]	desc_1_xuser_4_xuser_f;
wire [31:0]	desc_1_xuser_5_xuser_f;
wire [31:0]	desc_1_xuser_6_xuser_f;
wire [31:0]	desc_1_xuser_7_xuser_f;
wire [31:0]	desc_1_xuser_8_xuser_f;
wire [31:0]	desc_1_xuser_9_xuser_f;
wire [31:0]	desc_1_xuser_10_xuser_f;
wire [31:0]	desc_1_xuser_11_xuser_f;
wire [31:0]	desc_1_xuser_12_xuser_f;
wire [31:0]	desc_1_xuser_13_xuser_f;
wire [31:0]	desc_1_xuser_14_xuser_f;
wire [31:0]	desc_1_xuser_15_xuser_f;
wire [0:0]	desc_2_txn_type_wr_strb_f;
wire [0:0]	desc_2_txn_type_wr_rd_f;
wire [3:0]	desc_2_attr_axregion_f;
wire [3:0]	desc_2_attr_axqos_f;
wire [2:0]	desc_2_attr_axprot_f;
wire [3:0]	desc_2_attr_axcache_f;
wire [1:0]	desc_2_attr_axlock_f;
wire [1:0]	desc_2_attr_axburst_f;
wire [31:0]	desc_2_axid_0_axid_f;
wire [31:0]	desc_2_axid_1_axid_f;
wire [31:0]	desc_2_axid_2_axid_f;
wire [31:0]	desc_2_axid_3_axid_f;
wire [31:0]	desc_2_axuser_0_axuser_f;
wire [31:0]	desc_2_axuser_1_axuser_f;
wire [31:0]	desc_2_axuser_2_axuser_f;
wire [31:0]	desc_2_axuser_3_axuser_f;
wire [31:0]	desc_2_axuser_4_axuser_f;
wire [31:0]	desc_2_axuser_5_axuser_f;
wire [31:0]	desc_2_axuser_6_axuser_f;
wire [31:0]	desc_2_axuser_7_axuser_f;
wire [31:0]	desc_2_axuser_8_axuser_f;
wire [31:0]	desc_2_axuser_9_axuser_f;
wire [31:0]	desc_2_axuser_10_axuser_f;
wire [31:0]	desc_2_axuser_11_axuser_f;
wire [31:0]	desc_2_axuser_12_axuser_f;
wire [31:0]	desc_2_axuser_13_axuser_f;
wire [31:0]	desc_2_axuser_14_axuser_f;
wire [31:0]	desc_2_axuser_15_axuser_f;
wire [15:0]	desc_2_size_txn_size_f;
wire [2:0]	desc_2_axsize_axsize_f;
wire [31:0]	desc_2_axaddr_0_addr_f;
wire [31:0]	desc_2_axaddr_1_addr_f;
wire [31:0]	desc_2_axaddr_2_addr_f;
wire [31:0]	desc_2_axaddr_3_addr_f;
wire [31:0]	desc_2_data_offset_addr_f;
wire [31:0]	desc_2_wuser_0_wuser_f;
wire [31:0]	desc_2_wuser_1_wuser_f;
wire [31:0]	desc_2_wuser_2_wuser_f;
wire [31:0]	desc_2_wuser_3_wuser_f;
wire [31:0]	desc_2_wuser_4_wuser_f;
wire [31:0]	desc_2_wuser_5_wuser_f;
wire [31:0]	desc_2_wuser_6_wuser_f;
wire [31:0]	desc_2_wuser_7_wuser_f;
wire [31:0]	desc_2_wuser_8_wuser_f;
wire [31:0]	desc_2_wuser_9_wuser_f;
wire [31:0]	desc_2_wuser_10_wuser_f;
wire [31:0]	desc_2_wuser_11_wuser_f;
wire [31:0]	desc_2_wuser_12_wuser_f;
wire [31:0]	desc_2_wuser_13_wuser_f;
wire [31:0]	desc_2_wuser_14_wuser_f;
wire [31:0]	desc_2_wuser_15_wuser_f;
wire [31:0]	desc_2_data_host_addr_0_addr_f;
wire [31:0]	desc_2_data_host_addr_1_addr_f;
wire [31:0]	desc_2_data_host_addr_2_addr_f;
wire [31:0]	desc_2_data_host_addr_3_addr_f;
wire [31:0]	desc_2_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_2_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_2_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_2_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_2_xuser_0_xuser_f;
wire [31:0]	desc_2_xuser_1_xuser_f;
wire [31:0]	desc_2_xuser_2_xuser_f;
wire [31:0]	desc_2_xuser_3_xuser_f;
wire [31:0]	desc_2_xuser_4_xuser_f;
wire [31:0]	desc_2_xuser_5_xuser_f;
wire [31:0]	desc_2_xuser_6_xuser_f;
wire [31:0]	desc_2_xuser_7_xuser_f;
wire [31:0]	desc_2_xuser_8_xuser_f;
wire [31:0]	desc_2_xuser_9_xuser_f;
wire [31:0]	desc_2_xuser_10_xuser_f;
wire [31:0]	desc_2_xuser_11_xuser_f;
wire [31:0]	desc_2_xuser_12_xuser_f;
wire [31:0]	desc_2_xuser_13_xuser_f;
wire [31:0]	desc_2_xuser_14_xuser_f;
wire [31:0]	desc_2_xuser_15_xuser_f;
wire [0:0]	desc_3_txn_type_wr_strb_f;
wire [0:0]	desc_3_txn_type_wr_rd_f;
wire [3:0]	desc_3_attr_axregion_f;
wire [3:0]	desc_3_attr_axqos_f;
wire [2:0]	desc_3_attr_axprot_f;
wire [3:0]	desc_3_attr_axcache_f;
wire [1:0]	desc_3_attr_axlock_f;
wire [1:0]	desc_3_attr_axburst_f;
wire [31:0]	desc_3_axid_0_axid_f;
wire [31:0]	desc_3_axid_1_axid_f;
wire [31:0]	desc_3_axid_2_axid_f;
wire [31:0]	desc_3_axid_3_axid_f;
wire [31:0]	desc_3_axuser_0_axuser_f;
wire [31:0]	desc_3_axuser_1_axuser_f;
wire [31:0]	desc_3_axuser_2_axuser_f;
wire [31:0]	desc_3_axuser_3_axuser_f;
wire [31:0]	desc_3_axuser_4_axuser_f;
wire [31:0]	desc_3_axuser_5_axuser_f;
wire [31:0]	desc_3_axuser_6_axuser_f;
wire [31:0]	desc_3_axuser_7_axuser_f;
wire [31:0]	desc_3_axuser_8_axuser_f;
wire [31:0]	desc_3_axuser_9_axuser_f;
wire [31:0]	desc_3_axuser_10_axuser_f;
wire [31:0]	desc_3_axuser_11_axuser_f;
wire [31:0]	desc_3_axuser_12_axuser_f;
wire [31:0]	desc_3_axuser_13_axuser_f;
wire [31:0]	desc_3_axuser_14_axuser_f;
wire [31:0]	desc_3_axuser_15_axuser_f;
wire [15:0]	desc_3_size_txn_size_f;
wire [2:0]	desc_3_axsize_axsize_f;
wire [31:0]	desc_3_axaddr_0_addr_f;
wire [31:0]	desc_3_axaddr_1_addr_f;
wire [31:0]	desc_3_axaddr_2_addr_f;
wire [31:0]	desc_3_axaddr_3_addr_f;
wire [31:0]	desc_3_data_offset_addr_f;
wire [31:0]	desc_3_wuser_0_wuser_f;
wire [31:0]	desc_3_wuser_1_wuser_f;
wire [31:0]	desc_3_wuser_2_wuser_f;
wire [31:0]	desc_3_wuser_3_wuser_f;
wire [31:0]	desc_3_wuser_4_wuser_f;
wire [31:0]	desc_3_wuser_5_wuser_f;
wire [31:0]	desc_3_wuser_6_wuser_f;
wire [31:0]	desc_3_wuser_7_wuser_f;
wire [31:0]	desc_3_wuser_8_wuser_f;
wire [31:0]	desc_3_wuser_9_wuser_f;
wire [31:0]	desc_3_wuser_10_wuser_f;
wire [31:0]	desc_3_wuser_11_wuser_f;
wire [31:0]	desc_3_wuser_12_wuser_f;
wire [31:0]	desc_3_wuser_13_wuser_f;
wire [31:0]	desc_3_wuser_14_wuser_f;
wire [31:0]	desc_3_wuser_15_wuser_f;
wire [31:0]	desc_3_data_host_addr_0_addr_f;
wire [31:0]	desc_3_data_host_addr_1_addr_f;
wire [31:0]	desc_3_data_host_addr_2_addr_f;
wire [31:0]	desc_3_data_host_addr_3_addr_f;
wire [31:0]	desc_3_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_3_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_3_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_3_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_3_xuser_0_xuser_f;
wire [31:0]	desc_3_xuser_1_xuser_f;
wire [31:0]	desc_3_xuser_2_xuser_f;
wire [31:0]	desc_3_xuser_3_xuser_f;
wire [31:0]	desc_3_xuser_4_xuser_f;
wire [31:0]	desc_3_xuser_5_xuser_f;
wire [31:0]	desc_3_xuser_6_xuser_f;
wire [31:0]	desc_3_xuser_7_xuser_f;
wire [31:0]	desc_3_xuser_8_xuser_f;
wire [31:0]	desc_3_xuser_9_xuser_f;
wire [31:0]	desc_3_xuser_10_xuser_f;
wire [31:0]	desc_3_xuser_11_xuser_f;
wire [31:0]	desc_3_xuser_12_xuser_f;
wire [31:0]	desc_3_xuser_13_xuser_f;
wire [31:0]	desc_3_xuser_14_xuser_f;
wire [31:0]	desc_3_xuser_15_xuser_f;
wire [0:0]	desc_4_txn_type_wr_strb_f;
wire [0:0]	desc_4_txn_type_wr_rd_f;
wire [3:0]	desc_4_attr_axregion_f;
wire [3:0]	desc_4_attr_axqos_f;
wire [2:0]	desc_4_attr_axprot_f;
wire [3:0]	desc_4_attr_axcache_f;
wire [1:0]	desc_4_attr_axlock_f;
wire [1:0]	desc_4_attr_axburst_f;
wire [31:0]	desc_4_axid_0_axid_f;
wire [31:0]	desc_4_axid_1_axid_f;
wire [31:0]	desc_4_axid_2_axid_f;
wire [31:0]	desc_4_axid_3_axid_f;
wire [31:0]	desc_4_axuser_0_axuser_f;
wire [31:0]	desc_4_axuser_1_axuser_f;
wire [31:0]	desc_4_axuser_2_axuser_f;
wire [31:0]	desc_4_axuser_3_axuser_f;
wire [31:0]	desc_4_axuser_4_axuser_f;
wire [31:0]	desc_4_axuser_5_axuser_f;
wire [31:0]	desc_4_axuser_6_axuser_f;
wire [31:0]	desc_4_axuser_7_axuser_f;
wire [31:0]	desc_4_axuser_8_axuser_f;
wire [31:0]	desc_4_axuser_9_axuser_f;
wire [31:0]	desc_4_axuser_10_axuser_f;
wire [31:0]	desc_4_axuser_11_axuser_f;
wire [31:0]	desc_4_axuser_12_axuser_f;
wire [31:0]	desc_4_axuser_13_axuser_f;
wire [31:0]	desc_4_axuser_14_axuser_f;
wire [31:0]	desc_4_axuser_15_axuser_f;
wire [15:0]	desc_4_size_txn_size_f;
wire [2:0]	desc_4_axsize_axsize_f;
wire [31:0]	desc_4_axaddr_0_addr_f;
wire [31:0]	desc_4_axaddr_1_addr_f;
wire [31:0]	desc_4_axaddr_2_addr_f;
wire [31:0]	desc_4_axaddr_3_addr_f;
wire [31:0]	desc_4_data_offset_addr_f;
wire [31:0]	desc_4_wuser_0_wuser_f;
wire [31:0]	desc_4_wuser_1_wuser_f;
wire [31:0]	desc_4_wuser_2_wuser_f;
wire [31:0]	desc_4_wuser_3_wuser_f;
wire [31:0]	desc_4_wuser_4_wuser_f;
wire [31:0]	desc_4_wuser_5_wuser_f;
wire [31:0]	desc_4_wuser_6_wuser_f;
wire [31:0]	desc_4_wuser_7_wuser_f;
wire [31:0]	desc_4_wuser_8_wuser_f;
wire [31:0]	desc_4_wuser_9_wuser_f;
wire [31:0]	desc_4_wuser_10_wuser_f;
wire [31:0]	desc_4_wuser_11_wuser_f;
wire [31:0]	desc_4_wuser_12_wuser_f;
wire [31:0]	desc_4_wuser_13_wuser_f;
wire [31:0]	desc_4_wuser_14_wuser_f;
wire [31:0]	desc_4_wuser_15_wuser_f;
wire [31:0]	desc_4_data_host_addr_0_addr_f;
wire [31:0]	desc_4_data_host_addr_1_addr_f;
wire [31:0]	desc_4_data_host_addr_2_addr_f;
wire [31:0]	desc_4_data_host_addr_3_addr_f;
wire [31:0]	desc_4_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_4_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_4_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_4_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_4_xuser_0_xuser_f;
wire [31:0]	desc_4_xuser_1_xuser_f;
wire [31:0]	desc_4_xuser_2_xuser_f;
wire [31:0]	desc_4_xuser_3_xuser_f;
wire [31:0]	desc_4_xuser_4_xuser_f;
wire [31:0]	desc_4_xuser_5_xuser_f;
wire [31:0]	desc_4_xuser_6_xuser_f;
wire [31:0]	desc_4_xuser_7_xuser_f;
wire [31:0]	desc_4_xuser_8_xuser_f;
wire [31:0]	desc_4_xuser_9_xuser_f;
wire [31:0]	desc_4_xuser_10_xuser_f;
wire [31:0]	desc_4_xuser_11_xuser_f;
wire [31:0]	desc_4_xuser_12_xuser_f;
wire [31:0]	desc_4_xuser_13_xuser_f;
wire [31:0]	desc_4_xuser_14_xuser_f;
wire [31:0]	desc_4_xuser_15_xuser_f;
wire [0:0]	desc_5_txn_type_wr_strb_f;
wire [0:0]	desc_5_txn_type_wr_rd_f;
wire [3:0]	desc_5_attr_axregion_f;
wire [3:0]	desc_5_attr_axqos_f;
wire [2:0]	desc_5_attr_axprot_f;
wire [3:0]	desc_5_attr_axcache_f;
wire [1:0]	desc_5_attr_axlock_f;
wire [1:0]	desc_5_attr_axburst_f;
wire [31:0]	desc_5_axid_0_axid_f;
wire [31:0]	desc_5_axid_1_axid_f;
wire [31:0]	desc_5_axid_2_axid_f;
wire [31:0]	desc_5_axid_3_axid_f;
wire [31:0]	desc_5_axuser_0_axuser_f;
wire [31:0]	desc_5_axuser_1_axuser_f;
wire [31:0]	desc_5_axuser_2_axuser_f;
wire [31:0]	desc_5_axuser_3_axuser_f;
wire [31:0]	desc_5_axuser_4_axuser_f;
wire [31:0]	desc_5_axuser_5_axuser_f;
wire [31:0]	desc_5_axuser_6_axuser_f;
wire [31:0]	desc_5_axuser_7_axuser_f;
wire [31:0]	desc_5_axuser_8_axuser_f;
wire [31:0]	desc_5_axuser_9_axuser_f;
wire [31:0]	desc_5_axuser_10_axuser_f;
wire [31:0]	desc_5_axuser_11_axuser_f;
wire [31:0]	desc_5_axuser_12_axuser_f;
wire [31:0]	desc_5_axuser_13_axuser_f;
wire [31:0]	desc_5_axuser_14_axuser_f;
wire [31:0]	desc_5_axuser_15_axuser_f;
wire [15:0]	desc_5_size_txn_size_f;
wire [2:0]	desc_5_axsize_axsize_f;
wire [31:0]	desc_5_axaddr_0_addr_f;
wire [31:0]	desc_5_axaddr_1_addr_f;
wire [31:0]	desc_5_axaddr_2_addr_f;
wire [31:0]	desc_5_axaddr_3_addr_f;
wire [31:0]	desc_5_data_offset_addr_f;
wire [31:0]	desc_5_wuser_0_wuser_f;
wire [31:0]	desc_5_wuser_1_wuser_f;
wire [31:0]	desc_5_wuser_2_wuser_f;
wire [31:0]	desc_5_wuser_3_wuser_f;
wire [31:0]	desc_5_wuser_4_wuser_f;
wire [31:0]	desc_5_wuser_5_wuser_f;
wire [31:0]	desc_5_wuser_6_wuser_f;
wire [31:0]	desc_5_wuser_7_wuser_f;
wire [31:0]	desc_5_wuser_8_wuser_f;
wire [31:0]	desc_5_wuser_9_wuser_f;
wire [31:0]	desc_5_wuser_10_wuser_f;
wire [31:0]	desc_5_wuser_11_wuser_f;
wire [31:0]	desc_5_wuser_12_wuser_f;
wire [31:0]	desc_5_wuser_13_wuser_f;
wire [31:0]	desc_5_wuser_14_wuser_f;
wire [31:0]	desc_5_wuser_15_wuser_f;
wire [31:0]	desc_5_data_host_addr_0_addr_f;
wire [31:0]	desc_5_data_host_addr_1_addr_f;
wire [31:0]	desc_5_data_host_addr_2_addr_f;
wire [31:0]	desc_5_data_host_addr_3_addr_f;
wire [31:0]	desc_5_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_5_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_5_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_5_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_5_xuser_0_xuser_f;
wire [31:0]	desc_5_xuser_1_xuser_f;
wire [31:0]	desc_5_xuser_2_xuser_f;
wire [31:0]	desc_5_xuser_3_xuser_f;
wire [31:0]	desc_5_xuser_4_xuser_f;
wire [31:0]	desc_5_xuser_5_xuser_f;
wire [31:0]	desc_5_xuser_6_xuser_f;
wire [31:0]	desc_5_xuser_7_xuser_f;
wire [31:0]	desc_5_xuser_8_xuser_f;
wire [31:0]	desc_5_xuser_9_xuser_f;
wire [31:0]	desc_5_xuser_10_xuser_f;
wire [31:0]	desc_5_xuser_11_xuser_f;
wire [31:0]	desc_5_xuser_12_xuser_f;
wire [31:0]	desc_5_xuser_13_xuser_f;
wire [31:0]	desc_5_xuser_14_xuser_f;
wire [31:0]	desc_5_xuser_15_xuser_f;
wire [0:0]	desc_6_txn_type_wr_strb_f;
wire [0:0]	desc_6_txn_type_wr_rd_f;
wire [3:0]	desc_6_attr_axregion_f;
wire [3:0]	desc_6_attr_axqos_f;
wire [2:0]	desc_6_attr_axprot_f;
wire [3:0]	desc_6_attr_axcache_f;
wire [1:0]	desc_6_attr_axlock_f;
wire [1:0]	desc_6_attr_axburst_f;
wire [31:0]	desc_6_axid_0_axid_f;
wire [31:0]	desc_6_axid_1_axid_f;
wire [31:0]	desc_6_axid_2_axid_f;
wire [31:0]	desc_6_axid_3_axid_f;
wire [31:0]	desc_6_axuser_0_axuser_f;
wire [31:0]	desc_6_axuser_1_axuser_f;
wire [31:0]	desc_6_axuser_2_axuser_f;
wire [31:0]	desc_6_axuser_3_axuser_f;
wire [31:0]	desc_6_axuser_4_axuser_f;
wire [31:0]	desc_6_axuser_5_axuser_f;
wire [31:0]	desc_6_axuser_6_axuser_f;
wire [31:0]	desc_6_axuser_7_axuser_f;
wire [31:0]	desc_6_axuser_8_axuser_f;
wire [31:0]	desc_6_axuser_9_axuser_f;
wire [31:0]	desc_6_axuser_10_axuser_f;
wire [31:0]	desc_6_axuser_11_axuser_f;
wire [31:0]	desc_6_axuser_12_axuser_f;
wire [31:0]	desc_6_axuser_13_axuser_f;
wire [31:0]	desc_6_axuser_14_axuser_f;
wire [31:0]	desc_6_axuser_15_axuser_f;
wire [15:0]	desc_6_size_txn_size_f;
wire [2:0]	desc_6_axsize_axsize_f;
wire [31:0]	desc_6_axaddr_0_addr_f;
wire [31:0]	desc_6_axaddr_1_addr_f;
wire [31:0]	desc_6_axaddr_2_addr_f;
wire [31:0]	desc_6_axaddr_3_addr_f;
wire [31:0]	desc_6_data_offset_addr_f;
wire [31:0]	desc_6_wuser_0_wuser_f;
wire [31:0]	desc_6_wuser_1_wuser_f;
wire [31:0]	desc_6_wuser_2_wuser_f;
wire [31:0]	desc_6_wuser_3_wuser_f;
wire [31:0]	desc_6_wuser_4_wuser_f;
wire [31:0]	desc_6_wuser_5_wuser_f;
wire [31:0]	desc_6_wuser_6_wuser_f;
wire [31:0]	desc_6_wuser_7_wuser_f;
wire [31:0]	desc_6_wuser_8_wuser_f;
wire [31:0]	desc_6_wuser_9_wuser_f;
wire [31:0]	desc_6_wuser_10_wuser_f;
wire [31:0]	desc_6_wuser_11_wuser_f;
wire [31:0]	desc_6_wuser_12_wuser_f;
wire [31:0]	desc_6_wuser_13_wuser_f;
wire [31:0]	desc_6_wuser_14_wuser_f;
wire [31:0]	desc_6_wuser_15_wuser_f;
wire [31:0]	desc_6_data_host_addr_0_addr_f;
wire [31:0]	desc_6_data_host_addr_1_addr_f;
wire [31:0]	desc_6_data_host_addr_2_addr_f;
wire [31:0]	desc_6_data_host_addr_3_addr_f;
wire [31:0]	desc_6_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_6_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_6_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_6_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_6_xuser_0_xuser_f;
wire [31:0]	desc_6_xuser_1_xuser_f;
wire [31:0]	desc_6_xuser_2_xuser_f;
wire [31:0]	desc_6_xuser_3_xuser_f;
wire [31:0]	desc_6_xuser_4_xuser_f;
wire [31:0]	desc_6_xuser_5_xuser_f;
wire [31:0]	desc_6_xuser_6_xuser_f;
wire [31:0]	desc_6_xuser_7_xuser_f;
wire [31:0]	desc_6_xuser_8_xuser_f;
wire [31:0]	desc_6_xuser_9_xuser_f;
wire [31:0]	desc_6_xuser_10_xuser_f;
wire [31:0]	desc_6_xuser_11_xuser_f;
wire [31:0]	desc_6_xuser_12_xuser_f;
wire [31:0]	desc_6_xuser_13_xuser_f;
wire [31:0]	desc_6_xuser_14_xuser_f;
wire [31:0]	desc_6_xuser_15_xuser_f;
wire [0:0]	desc_7_txn_type_wr_strb_f;
wire [0:0]	desc_7_txn_type_wr_rd_f;
wire [3:0]	desc_7_attr_axregion_f;
wire [3:0]	desc_7_attr_axqos_f;
wire [2:0]	desc_7_attr_axprot_f;
wire [3:0]	desc_7_attr_axcache_f;
wire [1:0]	desc_7_attr_axlock_f;
wire [1:0]	desc_7_attr_axburst_f;
wire [31:0]	desc_7_axid_0_axid_f;
wire [31:0]	desc_7_axid_1_axid_f;
wire [31:0]	desc_7_axid_2_axid_f;
wire [31:0]	desc_7_axid_3_axid_f;
wire [31:0]	desc_7_axuser_0_axuser_f;
wire [31:0]	desc_7_axuser_1_axuser_f;
wire [31:0]	desc_7_axuser_2_axuser_f;
wire [31:0]	desc_7_axuser_3_axuser_f;
wire [31:0]	desc_7_axuser_4_axuser_f;
wire [31:0]	desc_7_axuser_5_axuser_f;
wire [31:0]	desc_7_axuser_6_axuser_f;
wire [31:0]	desc_7_axuser_7_axuser_f;
wire [31:0]	desc_7_axuser_8_axuser_f;
wire [31:0]	desc_7_axuser_9_axuser_f;
wire [31:0]	desc_7_axuser_10_axuser_f;
wire [31:0]	desc_7_axuser_11_axuser_f;
wire [31:0]	desc_7_axuser_12_axuser_f;
wire [31:0]	desc_7_axuser_13_axuser_f;
wire [31:0]	desc_7_axuser_14_axuser_f;
wire [31:0]	desc_7_axuser_15_axuser_f;
wire [15:0]	desc_7_size_txn_size_f;
wire [2:0]	desc_7_axsize_axsize_f;
wire [31:0]	desc_7_axaddr_0_addr_f;
wire [31:0]	desc_7_axaddr_1_addr_f;
wire [31:0]	desc_7_axaddr_2_addr_f;
wire [31:0]	desc_7_axaddr_3_addr_f;
wire [31:0]	desc_7_data_offset_addr_f;
wire [31:0]	desc_7_wuser_0_wuser_f;
wire [31:0]	desc_7_wuser_1_wuser_f;
wire [31:0]	desc_7_wuser_2_wuser_f;
wire [31:0]	desc_7_wuser_3_wuser_f;
wire [31:0]	desc_7_wuser_4_wuser_f;
wire [31:0]	desc_7_wuser_5_wuser_f;
wire [31:0]	desc_7_wuser_6_wuser_f;
wire [31:0]	desc_7_wuser_7_wuser_f;
wire [31:0]	desc_7_wuser_8_wuser_f;
wire [31:0]	desc_7_wuser_9_wuser_f;
wire [31:0]	desc_7_wuser_10_wuser_f;
wire [31:0]	desc_7_wuser_11_wuser_f;
wire [31:0]	desc_7_wuser_12_wuser_f;
wire [31:0]	desc_7_wuser_13_wuser_f;
wire [31:0]	desc_7_wuser_14_wuser_f;
wire [31:0]	desc_7_wuser_15_wuser_f;
wire [31:0]	desc_7_data_host_addr_0_addr_f;
wire [31:0]	desc_7_data_host_addr_1_addr_f;
wire [31:0]	desc_7_data_host_addr_2_addr_f;
wire [31:0]	desc_7_data_host_addr_3_addr_f;
wire [31:0]	desc_7_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_7_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_7_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_7_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_7_xuser_0_xuser_f;
wire [31:0]	desc_7_xuser_1_xuser_f;
wire [31:0]	desc_7_xuser_2_xuser_f;
wire [31:0]	desc_7_xuser_3_xuser_f;
wire [31:0]	desc_7_xuser_4_xuser_f;
wire [31:0]	desc_7_xuser_5_xuser_f;
wire [31:0]	desc_7_xuser_6_xuser_f;
wire [31:0]	desc_7_xuser_7_xuser_f;
wire [31:0]	desc_7_xuser_8_xuser_f;
wire [31:0]	desc_7_xuser_9_xuser_f;
wire [31:0]	desc_7_xuser_10_xuser_f;
wire [31:0]	desc_7_xuser_11_xuser_f;
wire [31:0]	desc_7_xuser_12_xuser_f;
wire [31:0]	desc_7_xuser_13_xuser_f;
wire [31:0]	desc_7_xuser_14_xuser_f;
wire [31:0]	desc_7_xuser_15_xuser_f;
wire [0:0]	desc_8_txn_type_wr_strb_f;
wire [0:0]	desc_8_txn_type_wr_rd_f;
wire [3:0]	desc_8_attr_axregion_f;
wire [3:0]	desc_8_attr_axqos_f;
wire [2:0]	desc_8_attr_axprot_f;
wire [3:0]	desc_8_attr_axcache_f;
wire [1:0]	desc_8_attr_axlock_f;
wire [1:0]	desc_8_attr_axburst_f;
wire [31:0]	desc_8_axid_0_axid_f;
wire [31:0]	desc_8_axid_1_axid_f;
wire [31:0]	desc_8_axid_2_axid_f;
wire [31:0]	desc_8_axid_3_axid_f;
wire [31:0]	desc_8_axuser_0_axuser_f;
wire [31:0]	desc_8_axuser_1_axuser_f;
wire [31:0]	desc_8_axuser_2_axuser_f;
wire [31:0]	desc_8_axuser_3_axuser_f;
wire [31:0]	desc_8_axuser_4_axuser_f;
wire [31:0]	desc_8_axuser_5_axuser_f;
wire [31:0]	desc_8_axuser_6_axuser_f;
wire [31:0]	desc_8_axuser_7_axuser_f;
wire [31:0]	desc_8_axuser_8_axuser_f;
wire [31:0]	desc_8_axuser_9_axuser_f;
wire [31:0]	desc_8_axuser_10_axuser_f;
wire [31:0]	desc_8_axuser_11_axuser_f;
wire [31:0]	desc_8_axuser_12_axuser_f;
wire [31:0]	desc_8_axuser_13_axuser_f;
wire [31:0]	desc_8_axuser_14_axuser_f;
wire [31:0]	desc_8_axuser_15_axuser_f;
wire [15:0]	desc_8_size_txn_size_f;
wire [2:0]	desc_8_axsize_axsize_f;
wire [31:0]	desc_8_axaddr_0_addr_f;
wire [31:0]	desc_8_axaddr_1_addr_f;
wire [31:0]	desc_8_axaddr_2_addr_f;
wire [31:0]	desc_8_axaddr_3_addr_f;
wire [31:0]	desc_8_data_offset_addr_f;
wire [31:0]	desc_8_wuser_0_wuser_f;
wire [31:0]	desc_8_wuser_1_wuser_f;
wire [31:0]	desc_8_wuser_2_wuser_f;
wire [31:0]	desc_8_wuser_3_wuser_f;
wire [31:0]	desc_8_wuser_4_wuser_f;
wire [31:0]	desc_8_wuser_5_wuser_f;
wire [31:0]	desc_8_wuser_6_wuser_f;
wire [31:0]	desc_8_wuser_7_wuser_f;
wire [31:0]	desc_8_wuser_8_wuser_f;
wire [31:0]	desc_8_wuser_9_wuser_f;
wire [31:0]	desc_8_wuser_10_wuser_f;
wire [31:0]	desc_8_wuser_11_wuser_f;
wire [31:0]	desc_8_wuser_12_wuser_f;
wire [31:0]	desc_8_wuser_13_wuser_f;
wire [31:0]	desc_8_wuser_14_wuser_f;
wire [31:0]	desc_8_wuser_15_wuser_f;
wire [31:0]	desc_8_data_host_addr_0_addr_f;
wire [31:0]	desc_8_data_host_addr_1_addr_f;
wire [31:0]	desc_8_data_host_addr_2_addr_f;
wire [31:0]	desc_8_data_host_addr_3_addr_f;
wire [31:0]	desc_8_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_8_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_8_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_8_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_8_xuser_0_xuser_f;
wire [31:0]	desc_8_xuser_1_xuser_f;
wire [31:0]	desc_8_xuser_2_xuser_f;
wire [31:0]	desc_8_xuser_3_xuser_f;
wire [31:0]	desc_8_xuser_4_xuser_f;
wire [31:0]	desc_8_xuser_5_xuser_f;
wire [31:0]	desc_8_xuser_6_xuser_f;
wire [31:0]	desc_8_xuser_7_xuser_f;
wire [31:0]	desc_8_xuser_8_xuser_f;
wire [31:0]	desc_8_xuser_9_xuser_f;
wire [31:0]	desc_8_xuser_10_xuser_f;
wire [31:0]	desc_8_xuser_11_xuser_f;
wire [31:0]	desc_8_xuser_12_xuser_f;
wire [31:0]	desc_8_xuser_13_xuser_f;
wire [31:0]	desc_8_xuser_14_xuser_f;
wire [31:0]	desc_8_xuser_15_xuser_f;
wire [0:0]	desc_9_txn_type_wr_strb_f;
wire [0:0]	desc_9_txn_type_wr_rd_f;
wire [3:0]	desc_9_attr_axregion_f;
wire [3:0]	desc_9_attr_axqos_f;
wire [2:0]	desc_9_attr_axprot_f;
wire [3:0]	desc_9_attr_axcache_f;
wire [1:0]	desc_9_attr_axlock_f;
wire [1:0]	desc_9_attr_axburst_f;
wire [31:0]	desc_9_axid_0_axid_f;
wire [31:0]	desc_9_axid_1_axid_f;
wire [31:0]	desc_9_axid_2_axid_f;
wire [31:0]	desc_9_axid_3_axid_f;
wire [31:0]	desc_9_axuser_0_axuser_f;
wire [31:0]	desc_9_axuser_1_axuser_f;
wire [31:0]	desc_9_axuser_2_axuser_f;
wire [31:0]	desc_9_axuser_3_axuser_f;
wire [31:0]	desc_9_axuser_4_axuser_f;
wire [31:0]	desc_9_axuser_5_axuser_f;
wire [31:0]	desc_9_axuser_6_axuser_f;
wire [31:0]	desc_9_axuser_7_axuser_f;
wire [31:0]	desc_9_axuser_8_axuser_f;
wire [31:0]	desc_9_axuser_9_axuser_f;
wire [31:0]	desc_9_axuser_10_axuser_f;
wire [31:0]	desc_9_axuser_11_axuser_f;
wire [31:0]	desc_9_axuser_12_axuser_f;
wire [31:0]	desc_9_axuser_13_axuser_f;
wire [31:0]	desc_9_axuser_14_axuser_f;
wire [31:0]	desc_9_axuser_15_axuser_f;
wire [15:0]	desc_9_size_txn_size_f;
wire [2:0]	desc_9_axsize_axsize_f;
wire [31:0]	desc_9_axaddr_0_addr_f;
wire [31:0]	desc_9_axaddr_1_addr_f;
wire [31:0]	desc_9_axaddr_2_addr_f;
wire [31:0]	desc_9_axaddr_3_addr_f;
wire [31:0]	desc_9_data_offset_addr_f;
wire [31:0]	desc_9_wuser_0_wuser_f;
wire [31:0]	desc_9_wuser_1_wuser_f;
wire [31:0]	desc_9_wuser_2_wuser_f;
wire [31:0]	desc_9_wuser_3_wuser_f;
wire [31:0]	desc_9_wuser_4_wuser_f;
wire [31:0]	desc_9_wuser_5_wuser_f;
wire [31:0]	desc_9_wuser_6_wuser_f;
wire [31:0]	desc_9_wuser_7_wuser_f;
wire [31:0]	desc_9_wuser_8_wuser_f;
wire [31:0]	desc_9_wuser_9_wuser_f;
wire [31:0]	desc_9_wuser_10_wuser_f;
wire [31:0]	desc_9_wuser_11_wuser_f;
wire [31:0]	desc_9_wuser_12_wuser_f;
wire [31:0]	desc_9_wuser_13_wuser_f;
wire [31:0]	desc_9_wuser_14_wuser_f;
wire [31:0]	desc_9_wuser_15_wuser_f;
wire [31:0]	desc_9_data_host_addr_0_addr_f;
wire [31:0]	desc_9_data_host_addr_1_addr_f;
wire [31:0]	desc_9_data_host_addr_2_addr_f;
wire [31:0]	desc_9_data_host_addr_3_addr_f;
wire [31:0]	desc_9_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_9_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_9_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_9_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_9_xuser_0_xuser_f;
wire [31:0]	desc_9_xuser_1_xuser_f;
wire [31:0]	desc_9_xuser_2_xuser_f;
wire [31:0]	desc_9_xuser_3_xuser_f;
wire [31:0]	desc_9_xuser_4_xuser_f;
wire [31:0]	desc_9_xuser_5_xuser_f;
wire [31:0]	desc_9_xuser_6_xuser_f;
wire [31:0]	desc_9_xuser_7_xuser_f;
wire [31:0]	desc_9_xuser_8_xuser_f;
wire [31:0]	desc_9_xuser_9_xuser_f;
wire [31:0]	desc_9_xuser_10_xuser_f;
wire [31:0]	desc_9_xuser_11_xuser_f;
wire [31:0]	desc_9_xuser_12_xuser_f;
wire [31:0]	desc_9_xuser_13_xuser_f;
wire [31:0]	desc_9_xuser_14_xuser_f;
wire [31:0]	desc_9_xuser_15_xuser_f;
wire [0:0]	desc_10_txn_type_wr_strb_f;
wire [0:0]	desc_10_txn_type_wr_rd_f;
wire [3:0]	desc_10_attr_axregion_f;
wire [3:0]	desc_10_attr_axqos_f;
wire [2:0]	desc_10_attr_axprot_f;
wire [3:0]	desc_10_attr_axcache_f;
wire [1:0]	desc_10_attr_axlock_f;
wire [1:0]	desc_10_attr_axburst_f;
wire [31:0]	desc_10_axid_0_axid_f;
wire [31:0]	desc_10_axid_1_axid_f;
wire [31:0]	desc_10_axid_2_axid_f;
wire [31:0]	desc_10_axid_3_axid_f;
wire [31:0]	desc_10_axuser_0_axuser_f;
wire [31:0]	desc_10_axuser_1_axuser_f;
wire [31:0]	desc_10_axuser_2_axuser_f;
wire [31:0]	desc_10_axuser_3_axuser_f;
wire [31:0]	desc_10_axuser_4_axuser_f;
wire [31:0]	desc_10_axuser_5_axuser_f;
wire [31:0]	desc_10_axuser_6_axuser_f;
wire [31:0]	desc_10_axuser_7_axuser_f;
wire [31:0]	desc_10_axuser_8_axuser_f;
wire [31:0]	desc_10_axuser_9_axuser_f;
wire [31:0]	desc_10_axuser_10_axuser_f;
wire [31:0]	desc_10_axuser_11_axuser_f;
wire [31:0]	desc_10_axuser_12_axuser_f;
wire [31:0]	desc_10_axuser_13_axuser_f;
wire [31:0]	desc_10_axuser_14_axuser_f;
wire [31:0]	desc_10_axuser_15_axuser_f;
wire [15:0]	desc_10_size_txn_size_f;
wire [2:0]	desc_10_axsize_axsize_f;
wire [31:0]	desc_10_axaddr_0_addr_f;
wire [31:0]	desc_10_axaddr_1_addr_f;
wire [31:0]	desc_10_axaddr_2_addr_f;
wire [31:0]	desc_10_axaddr_3_addr_f;
wire [31:0]	desc_10_data_offset_addr_f;
wire [31:0]	desc_10_wuser_0_wuser_f;
wire [31:0]	desc_10_wuser_1_wuser_f;
wire [31:0]	desc_10_wuser_2_wuser_f;
wire [31:0]	desc_10_wuser_3_wuser_f;
wire [31:0]	desc_10_wuser_4_wuser_f;
wire [31:0]	desc_10_wuser_5_wuser_f;
wire [31:0]	desc_10_wuser_6_wuser_f;
wire [31:0]	desc_10_wuser_7_wuser_f;
wire [31:0]	desc_10_wuser_8_wuser_f;
wire [31:0]	desc_10_wuser_9_wuser_f;
wire [31:0]	desc_10_wuser_10_wuser_f;
wire [31:0]	desc_10_wuser_11_wuser_f;
wire [31:0]	desc_10_wuser_12_wuser_f;
wire [31:0]	desc_10_wuser_13_wuser_f;
wire [31:0]	desc_10_wuser_14_wuser_f;
wire [31:0]	desc_10_wuser_15_wuser_f;
wire [31:0]	desc_10_data_host_addr_0_addr_f;
wire [31:0]	desc_10_data_host_addr_1_addr_f;
wire [31:0]	desc_10_data_host_addr_2_addr_f;
wire [31:0]	desc_10_data_host_addr_3_addr_f;
wire [31:0]	desc_10_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_10_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_10_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_10_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_10_xuser_0_xuser_f;
wire [31:0]	desc_10_xuser_1_xuser_f;
wire [31:0]	desc_10_xuser_2_xuser_f;
wire [31:0]	desc_10_xuser_3_xuser_f;
wire [31:0]	desc_10_xuser_4_xuser_f;
wire [31:0]	desc_10_xuser_5_xuser_f;
wire [31:0]	desc_10_xuser_6_xuser_f;
wire [31:0]	desc_10_xuser_7_xuser_f;
wire [31:0]	desc_10_xuser_8_xuser_f;
wire [31:0]	desc_10_xuser_9_xuser_f;
wire [31:0]	desc_10_xuser_10_xuser_f;
wire [31:0]	desc_10_xuser_11_xuser_f;
wire [31:0]	desc_10_xuser_12_xuser_f;
wire [31:0]	desc_10_xuser_13_xuser_f;
wire [31:0]	desc_10_xuser_14_xuser_f;
wire [31:0]	desc_10_xuser_15_xuser_f;
wire [0:0]	desc_11_txn_type_wr_strb_f;
wire [0:0]	desc_11_txn_type_wr_rd_f;
wire [3:0]	desc_11_attr_axregion_f;
wire [3:0]	desc_11_attr_axqos_f;
wire [2:0]	desc_11_attr_axprot_f;
wire [3:0]	desc_11_attr_axcache_f;
wire [1:0]	desc_11_attr_axlock_f;
wire [1:0]	desc_11_attr_axburst_f;
wire [31:0]	desc_11_axid_0_axid_f;
wire [31:0]	desc_11_axid_1_axid_f;
wire [31:0]	desc_11_axid_2_axid_f;
wire [31:0]	desc_11_axid_3_axid_f;
wire [31:0]	desc_11_axuser_0_axuser_f;
wire [31:0]	desc_11_axuser_1_axuser_f;
wire [31:0]	desc_11_axuser_2_axuser_f;
wire [31:0]	desc_11_axuser_3_axuser_f;
wire [31:0]	desc_11_axuser_4_axuser_f;
wire [31:0]	desc_11_axuser_5_axuser_f;
wire [31:0]	desc_11_axuser_6_axuser_f;
wire [31:0]	desc_11_axuser_7_axuser_f;
wire [31:0]	desc_11_axuser_8_axuser_f;
wire [31:0]	desc_11_axuser_9_axuser_f;
wire [31:0]	desc_11_axuser_10_axuser_f;
wire [31:0]	desc_11_axuser_11_axuser_f;
wire [31:0]	desc_11_axuser_12_axuser_f;
wire [31:0]	desc_11_axuser_13_axuser_f;
wire [31:0]	desc_11_axuser_14_axuser_f;
wire [31:0]	desc_11_axuser_15_axuser_f;
wire [15:0]	desc_11_size_txn_size_f;
wire [2:0]	desc_11_axsize_axsize_f;
wire [31:0]	desc_11_axaddr_0_addr_f;
wire [31:0]	desc_11_axaddr_1_addr_f;
wire [31:0]	desc_11_axaddr_2_addr_f;
wire [31:0]	desc_11_axaddr_3_addr_f;
wire [31:0]	desc_11_data_offset_addr_f;
wire [31:0]	desc_11_wuser_0_wuser_f;
wire [31:0]	desc_11_wuser_1_wuser_f;
wire [31:0]	desc_11_wuser_2_wuser_f;
wire [31:0]	desc_11_wuser_3_wuser_f;
wire [31:0]	desc_11_wuser_4_wuser_f;
wire [31:0]	desc_11_wuser_5_wuser_f;
wire [31:0]	desc_11_wuser_6_wuser_f;
wire [31:0]	desc_11_wuser_7_wuser_f;
wire [31:0]	desc_11_wuser_8_wuser_f;
wire [31:0]	desc_11_wuser_9_wuser_f;
wire [31:0]	desc_11_wuser_10_wuser_f;
wire [31:0]	desc_11_wuser_11_wuser_f;
wire [31:0]	desc_11_wuser_12_wuser_f;
wire [31:0]	desc_11_wuser_13_wuser_f;
wire [31:0]	desc_11_wuser_14_wuser_f;
wire [31:0]	desc_11_wuser_15_wuser_f;
wire [31:0]	desc_11_data_host_addr_0_addr_f;
wire [31:0]	desc_11_data_host_addr_1_addr_f;
wire [31:0]	desc_11_data_host_addr_2_addr_f;
wire [31:0]	desc_11_data_host_addr_3_addr_f;
wire [31:0]	desc_11_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_11_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_11_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_11_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_11_xuser_0_xuser_f;
wire [31:0]	desc_11_xuser_1_xuser_f;
wire [31:0]	desc_11_xuser_2_xuser_f;
wire [31:0]	desc_11_xuser_3_xuser_f;
wire [31:0]	desc_11_xuser_4_xuser_f;
wire [31:0]	desc_11_xuser_5_xuser_f;
wire [31:0]	desc_11_xuser_6_xuser_f;
wire [31:0]	desc_11_xuser_7_xuser_f;
wire [31:0]	desc_11_xuser_8_xuser_f;
wire [31:0]	desc_11_xuser_9_xuser_f;
wire [31:0]	desc_11_xuser_10_xuser_f;
wire [31:0]	desc_11_xuser_11_xuser_f;
wire [31:0]	desc_11_xuser_12_xuser_f;
wire [31:0]	desc_11_xuser_13_xuser_f;
wire [31:0]	desc_11_xuser_14_xuser_f;
wire [31:0]	desc_11_xuser_15_xuser_f;
wire [0:0]	desc_12_txn_type_wr_strb_f;
wire [0:0]	desc_12_txn_type_wr_rd_f;
wire [3:0]	desc_12_attr_axregion_f;
wire [3:0]	desc_12_attr_axqos_f;
wire [2:0]	desc_12_attr_axprot_f;
wire [3:0]	desc_12_attr_axcache_f;
wire [1:0]	desc_12_attr_axlock_f;
wire [1:0]	desc_12_attr_axburst_f;
wire [31:0]	desc_12_axid_0_axid_f;
wire [31:0]	desc_12_axid_1_axid_f;
wire [31:0]	desc_12_axid_2_axid_f;
wire [31:0]	desc_12_axid_3_axid_f;
wire [31:0]	desc_12_axuser_0_axuser_f;
wire [31:0]	desc_12_axuser_1_axuser_f;
wire [31:0]	desc_12_axuser_2_axuser_f;
wire [31:0]	desc_12_axuser_3_axuser_f;
wire [31:0]	desc_12_axuser_4_axuser_f;
wire [31:0]	desc_12_axuser_5_axuser_f;
wire [31:0]	desc_12_axuser_6_axuser_f;
wire [31:0]	desc_12_axuser_7_axuser_f;
wire [31:0]	desc_12_axuser_8_axuser_f;
wire [31:0]	desc_12_axuser_9_axuser_f;
wire [31:0]	desc_12_axuser_10_axuser_f;
wire [31:0]	desc_12_axuser_11_axuser_f;
wire [31:0]	desc_12_axuser_12_axuser_f;
wire [31:0]	desc_12_axuser_13_axuser_f;
wire [31:0]	desc_12_axuser_14_axuser_f;
wire [31:0]	desc_12_axuser_15_axuser_f;
wire [15:0]	desc_12_size_txn_size_f;
wire [2:0]	desc_12_axsize_axsize_f;
wire [31:0]	desc_12_axaddr_0_addr_f;
wire [31:0]	desc_12_axaddr_1_addr_f;
wire [31:0]	desc_12_axaddr_2_addr_f;
wire [31:0]	desc_12_axaddr_3_addr_f;
wire [31:0]	desc_12_data_offset_addr_f;
wire [31:0]	desc_12_wuser_0_wuser_f;
wire [31:0]	desc_12_wuser_1_wuser_f;
wire [31:0]	desc_12_wuser_2_wuser_f;
wire [31:0]	desc_12_wuser_3_wuser_f;
wire [31:0]	desc_12_wuser_4_wuser_f;
wire [31:0]	desc_12_wuser_5_wuser_f;
wire [31:0]	desc_12_wuser_6_wuser_f;
wire [31:0]	desc_12_wuser_7_wuser_f;
wire [31:0]	desc_12_wuser_8_wuser_f;
wire [31:0]	desc_12_wuser_9_wuser_f;
wire [31:0]	desc_12_wuser_10_wuser_f;
wire [31:0]	desc_12_wuser_11_wuser_f;
wire [31:0]	desc_12_wuser_12_wuser_f;
wire [31:0]	desc_12_wuser_13_wuser_f;
wire [31:0]	desc_12_wuser_14_wuser_f;
wire [31:0]	desc_12_wuser_15_wuser_f;
wire [31:0]	desc_12_data_host_addr_0_addr_f;
wire [31:0]	desc_12_data_host_addr_1_addr_f;
wire [31:0]	desc_12_data_host_addr_2_addr_f;
wire [31:0]	desc_12_data_host_addr_3_addr_f;
wire [31:0]	desc_12_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_12_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_12_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_12_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_12_xuser_0_xuser_f;
wire [31:0]	desc_12_xuser_1_xuser_f;
wire [31:0]	desc_12_xuser_2_xuser_f;
wire [31:0]	desc_12_xuser_3_xuser_f;
wire [31:0]	desc_12_xuser_4_xuser_f;
wire [31:0]	desc_12_xuser_5_xuser_f;
wire [31:0]	desc_12_xuser_6_xuser_f;
wire [31:0]	desc_12_xuser_7_xuser_f;
wire [31:0]	desc_12_xuser_8_xuser_f;
wire [31:0]	desc_12_xuser_9_xuser_f;
wire [31:0]	desc_12_xuser_10_xuser_f;
wire [31:0]	desc_12_xuser_11_xuser_f;
wire [31:0]	desc_12_xuser_12_xuser_f;
wire [31:0]	desc_12_xuser_13_xuser_f;
wire [31:0]	desc_12_xuser_14_xuser_f;
wire [31:0]	desc_12_xuser_15_xuser_f;
wire [0:0]	desc_13_txn_type_wr_strb_f;
wire [0:0]	desc_13_txn_type_wr_rd_f;
wire [3:0]	desc_13_attr_axregion_f;
wire [3:0]	desc_13_attr_axqos_f;
wire [2:0]	desc_13_attr_axprot_f;
wire [3:0]	desc_13_attr_axcache_f;
wire [1:0]	desc_13_attr_axlock_f;
wire [1:0]	desc_13_attr_axburst_f;
wire [31:0]	desc_13_axid_0_axid_f;
wire [31:0]	desc_13_axid_1_axid_f;
wire [31:0]	desc_13_axid_2_axid_f;
wire [31:0]	desc_13_axid_3_axid_f;
wire [31:0]	desc_13_axuser_0_axuser_f;
wire [31:0]	desc_13_axuser_1_axuser_f;
wire [31:0]	desc_13_axuser_2_axuser_f;
wire [31:0]	desc_13_axuser_3_axuser_f;
wire [31:0]	desc_13_axuser_4_axuser_f;
wire [31:0]	desc_13_axuser_5_axuser_f;
wire [31:0]	desc_13_axuser_6_axuser_f;
wire [31:0]	desc_13_axuser_7_axuser_f;
wire [31:0]	desc_13_axuser_8_axuser_f;
wire [31:0]	desc_13_axuser_9_axuser_f;
wire [31:0]	desc_13_axuser_10_axuser_f;
wire [31:0]	desc_13_axuser_11_axuser_f;
wire [31:0]	desc_13_axuser_12_axuser_f;
wire [31:0]	desc_13_axuser_13_axuser_f;
wire [31:0]	desc_13_axuser_14_axuser_f;
wire [31:0]	desc_13_axuser_15_axuser_f;
wire [15:0]	desc_13_size_txn_size_f;
wire [2:0]	desc_13_axsize_axsize_f;
wire [31:0]	desc_13_axaddr_0_addr_f;
wire [31:0]	desc_13_axaddr_1_addr_f;
wire [31:0]	desc_13_axaddr_2_addr_f;
wire [31:0]	desc_13_axaddr_3_addr_f;
wire [31:0]	desc_13_data_offset_addr_f;
wire [31:0]	desc_13_wuser_0_wuser_f;
wire [31:0]	desc_13_wuser_1_wuser_f;
wire [31:0]	desc_13_wuser_2_wuser_f;
wire [31:0]	desc_13_wuser_3_wuser_f;
wire [31:0]	desc_13_wuser_4_wuser_f;
wire [31:0]	desc_13_wuser_5_wuser_f;
wire [31:0]	desc_13_wuser_6_wuser_f;
wire [31:0]	desc_13_wuser_7_wuser_f;
wire [31:0]	desc_13_wuser_8_wuser_f;
wire [31:0]	desc_13_wuser_9_wuser_f;
wire [31:0]	desc_13_wuser_10_wuser_f;
wire [31:0]	desc_13_wuser_11_wuser_f;
wire [31:0]	desc_13_wuser_12_wuser_f;
wire [31:0]	desc_13_wuser_13_wuser_f;
wire [31:0]	desc_13_wuser_14_wuser_f;
wire [31:0]	desc_13_wuser_15_wuser_f;
wire [31:0]	desc_13_data_host_addr_0_addr_f;
wire [31:0]	desc_13_data_host_addr_1_addr_f;
wire [31:0]	desc_13_data_host_addr_2_addr_f;
wire [31:0]	desc_13_data_host_addr_3_addr_f;
wire [31:0]	desc_13_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_13_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_13_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_13_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_13_xuser_0_xuser_f;
wire [31:0]	desc_13_xuser_1_xuser_f;
wire [31:0]	desc_13_xuser_2_xuser_f;
wire [31:0]	desc_13_xuser_3_xuser_f;
wire [31:0]	desc_13_xuser_4_xuser_f;
wire [31:0]	desc_13_xuser_5_xuser_f;
wire [31:0]	desc_13_xuser_6_xuser_f;
wire [31:0]	desc_13_xuser_7_xuser_f;
wire [31:0]	desc_13_xuser_8_xuser_f;
wire [31:0]	desc_13_xuser_9_xuser_f;
wire [31:0]	desc_13_xuser_10_xuser_f;
wire [31:0]	desc_13_xuser_11_xuser_f;
wire [31:0]	desc_13_xuser_12_xuser_f;
wire [31:0]	desc_13_xuser_13_xuser_f;
wire [31:0]	desc_13_xuser_14_xuser_f;
wire [31:0]	desc_13_xuser_15_xuser_f;
wire [0:0]	desc_14_txn_type_wr_strb_f;
wire [0:0]	desc_14_txn_type_wr_rd_f;
wire [3:0]	desc_14_attr_axregion_f;
wire [3:0]	desc_14_attr_axqos_f;
wire [2:0]	desc_14_attr_axprot_f;
wire [3:0]	desc_14_attr_axcache_f;
wire [1:0]	desc_14_attr_axlock_f;
wire [1:0]	desc_14_attr_axburst_f;
wire [31:0]	desc_14_axid_0_axid_f;
wire [31:0]	desc_14_axid_1_axid_f;
wire [31:0]	desc_14_axid_2_axid_f;
wire [31:0]	desc_14_axid_3_axid_f;
wire [31:0]	desc_14_axuser_0_axuser_f;
wire [31:0]	desc_14_axuser_1_axuser_f;
wire [31:0]	desc_14_axuser_2_axuser_f;
wire [31:0]	desc_14_axuser_3_axuser_f;
wire [31:0]	desc_14_axuser_4_axuser_f;
wire [31:0]	desc_14_axuser_5_axuser_f;
wire [31:0]	desc_14_axuser_6_axuser_f;
wire [31:0]	desc_14_axuser_7_axuser_f;
wire [31:0]	desc_14_axuser_8_axuser_f;
wire [31:0]	desc_14_axuser_9_axuser_f;
wire [31:0]	desc_14_axuser_10_axuser_f;
wire [31:0]	desc_14_axuser_11_axuser_f;
wire [31:0]	desc_14_axuser_12_axuser_f;
wire [31:0]	desc_14_axuser_13_axuser_f;
wire [31:0]	desc_14_axuser_14_axuser_f;
wire [31:0]	desc_14_axuser_15_axuser_f;
wire [15:0]	desc_14_size_txn_size_f;
wire [2:0]	desc_14_axsize_axsize_f;
wire [31:0]	desc_14_axaddr_0_addr_f;
wire [31:0]	desc_14_axaddr_1_addr_f;
wire [31:0]	desc_14_axaddr_2_addr_f;
wire [31:0]	desc_14_axaddr_3_addr_f;
wire [31:0]	desc_14_data_offset_addr_f;
wire [31:0]	desc_14_wuser_0_wuser_f;
wire [31:0]	desc_14_wuser_1_wuser_f;
wire [31:0]	desc_14_wuser_2_wuser_f;
wire [31:0]	desc_14_wuser_3_wuser_f;
wire [31:0]	desc_14_wuser_4_wuser_f;
wire [31:0]	desc_14_wuser_5_wuser_f;
wire [31:0]	desc_14_wuser_6_wuser_f;
wire [31:0]	desc_14_wuser_7_wuser_f;
wire [31:0]	desc_14_wuser_8_wuser_f;
wire [31:0]	desc_14_wuser_9_wuser_f;
wire [31:0]	desc_14_wuser_10_wuser_f;
wire [31:0]	desc_14_wuser_11_wuser_f;
wire [31:0]	desc_14_wuser_12_wuser_f;
wire [31:0]	desc_14_wuser_13_wuser_f;
wire [31:0]	desc_14_wuser_14_wuser_f;
wire [31:0]	desc_14_wuser_15_wuser_f;
wire [31:0]	desc_14_data_host_addr_0_addr_f;
wire [31:0]	desc_14_data_host_addr_1_addr_f;
wire [31:0]	desc_14_data_host_addr_2_addr_f;
wire [31:0]	desc_14_data_host_addr_3_addr_f;
wire [31:0]	desc_14_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_14_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_14_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_14_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_14_xuser_0_xuser_f;
wire [31:0]	desc_14_xuser_1_xuser_f;
wire [31:0]	desc_14_xuser_2_xuser_f;
wire [31:0]	desc_14_xuser_3_xuser_f;
wire [31:0]	desc_14_xuser_4_xuser_f;
wire [31:0]	desc_14_xuser_5_xuser_f;
wire [31:0]	desc_14_xuser_6_xuser_f;
wire [31:0]	desc_14_xuser_7_xuser_f;
wire [31:0]	desc_14_xuser_8_xuser_f;
wire [31:0]	desc_14_xuser_9_xuser_f;
wire [31:0]	desc_14_xuser_10_xuser_f;
wire [31:0]	desc_14_xuser_11_xuser_f;
wire [31:0]	desc_14_xuser_12_xuser_f;
wire [31:0]	desc_14_xuser_13_xuser_f;
wire [31:0]	desc_14_xuser_14_xuser_f;
wire [31:0]	desc_14_xuser_15_xuser_f;
wire [0:0]	desc_15_txn_type_wr_strb_f;
wire [0:0]	desc_15_txn_type_wr_rd_f;
wire [3:0]	desc_15_attr_axregion_f;
wire [3:0]	desc_15_attr_axqos_f;
wire [2:0]	desc_15_attr_axprot_f;
wire [3:0]	desc_15_attr_axcache_f;
wire [1:0]	desc_15_attr_axlock_f;
wire [1:0]	desc_15_attr_axburst_f;
wire [31:0]	desc_15_axid_0_axid_f;
wire [31:0]	desc_15_axid_1_axid_f;
wire [31:0]	desc_15_axid_2_axid_f;
wire [31:0]	desc_15_axid_3_axid_f;
wire [31:0]	desc_15_axuser_0_axuser_f;
wire [31:0]	desc_15_axuser_1_axuser_f;
wire [31:0]	desc_15_axuser_2_axuser_f;
wire [31:0]	desc_15_axuser_3_axuser_f;
wire [31:0]	desc_15_axuser_4_axuser_f;
wire [31:0]	desc_15_axuser_5_axuser_f;
wire [31:0]	desc_15_axuser_6_axuser_f;
wire [31:0]	desc_15_axuser_7_axuser_f;
wire [31:0]	desc_15_axuser_8_axuser_f;
wire [31:0]	desc_15_axuser_9_axuser_f;
wire [31:0]	desc_15_axuser_10_axuser_f;
wire [31:0]	desc_15_axuser_11_axuser_f;
wire [31:0]	desc_15_axuser_12_axuser_f;
wire [31:0]	desc_15_axuser_13_axuser_f;
wire [31:0]	desc_15_axuser_14_axuser_f;
wire [31:0]	desc_15_axuser_15_axuser_f;
wire [15:0]	desc_15_size_txn_size_f;
wire [2:0]	desc_15_axsize_axsize_f;
wire [31:0]	desc_15_axaddr_0_addr_f;
wire [31:0]	desc_15_axaddr_1_addr_f;
wire [31:0]	desc_15_axaddr_2_addr_f;
wire [31:0]	desc_15_axaddr_3_addr_f;
wire [31:0]	desc_15_data_offset_addr_f;
wire [31:0]	desc_15_wuser_0_wuser_f;
wire [31:0]	desc_15_wuser_1_wuser_f;
wire [31:0]	desc_15_wuser_2_wuser_f;
wire [31:0]	desc_15_wuser_3_wuser_f;
wire [31:0]	desc_15_wuser_4_wuser_f;
wire [31:0]	desc_15_wuser_5_wuser_f;
wire [31:0]	desc_15_wuser_6_wuser_f;
wire [31:0]	desc_15_wuser_7_wuser_f;
wire [31:0]	desc_15_wuser_8_wuser_f;
wire [31:0]	desc_15_wuser_9_wuser_f;
wire [31:0]	desc_15_wuser_10_wuser_f;
wire [31:0]	desc_15_wuser_11_wuser_f;
wire [31:0]	desc_15_wuser_12_wuser_f;
wire [31:0]	desc_15_wuser_13_wuser_f;
wire [31:0]	desc_15_wuser_14_wuser_f;
wire [31:0]	desc_15_wuser_15_wuser_f;
wire [31:0]	desc_15_data_host_addr_0_addr_f;
wire [31:0]	desc_15_data_host_addr_1_addr_f;
wire [31:0]	desc_15_data_host_addr_2_addr_f;
wire [31:0]	desc_15_data_host_addr_3_addr_f;
wire [31:0]	desc_15_wstrb_host_addr_0_addr_f;
wire [31:0]	desc_15_wstrb_host_addr_1_addr_f;
wire [31:0]	desc_15_wstrb_host_addr_2_addr_f;
wire [31:0]	desc_15_wstrb_host_addr_3_addr_f;
wire [31:0]	desc_15_xuser_0_xuser_f;
wire [31:0]	desc_15_xuser_1_xuser_f;
wire [31:0]	desc_15_xuser_2_xuser_f;
wire [31:0]	desc_15_xuser_3_xuser_f;
wire [31:0]	desc_15_xuser_4_xuser_f;
wire [31:0]	desc_15_xuser_5_xuser_f;
wire [31:0]	desc_15_xuser_6_xuser_f;
wire [31:0]	desc_15_xuser_7_xuser_f;
wire [31:0]	desc_15_xuser_8_xuser_f;
wire [31:0]	desc_15_xuser_9_xuser_f;
wire [31:0]	desc_15_xuser_10_xuser_f;
wire [31:0]	desc_15_xuser_11_xuser_f;
wire [31:0]	desc_15_xuser_12_xuser_f;
wire [31:0]	desc_15_xuser_13_xuser_f;
wire [31:0]	desc_15_xuser_14_xuser_f;
wire [31:0]	desc_15_xuser_15_xuser_f;

//Fields to use in entire slave RTL ( int_<reg>_<field> )
wire	[7:0]				int_version_major_ver;
wire	[7:0]				int_version_minor_ver;
wire	[7:0]				int_bridge_type_type;
wire	[7:0]				int_axi_bridge_config_user_width;
wire	[7:0]				int_axi_bridge_config_id_width;
wire	[2:0]				int_axi_bridge_config_data_width;
wire	     				int_reset_dut_srst_3;
wire	     				int_reset_dut_srst_2;
wire	     				int_reset_dut_srst_1;
wire	     				int_reset_dut_srst_0;
wire	     				int_reset_srst;
wire	     				int_mode_select_imm_bresp;
wire	     				int_mode_select_mode_2;
wire	     				int_mode_select_mode_0_1;
wire	[MAX_DESC-1:0]			int_ownership_own;
wire	[MAX_DESC-1:0]			int_ownership_flip_flip;
wire	[MAX_DESC-1:0]			int_status_resp_comp_resp_comp;
wire	[31:0]				int_status_resp_resp;
wire	[MAX_DESC-1:0]			int_status_busy_busy;
wire	[DESC_IDX_WIDTH:0]		int_resp_fifo_free_level_level;
wire	     				int_intr_status_comp;
wire	     				int_intr_status_c2h;
wire	     				int_intr_status_error;
wire	     				int_intr_status_txn_avail;
wire	[MAX_DESC-1:0]			int_intr_txn_avail_status_avail;
wire	[MAX_DESC-1:0]			int_intr_txn_avail_clear_clr_avail;
wire	[MAX_DESC-1:0]			int_intr_txn_avail_enable_en_avail;
wire	[MAX_DESC-1:0]			int_intr_comp_status_comp;
wire	[MAX_DESC-1:0]			int_intr_comp_clear_clr_comp;
wire	[MAX_DESC-1:0]			int_intr_comp_enable_en_comp;
wire	     				int_intr_error_status_err_2;
wire	     				int_intr_error_status_err_1;
wire	     				int_intr_error_status_err_0;
wire	     				int_intr_error_clear_clr_err_2;
wire	     				int_intr_error_clear_clr_err_1;
wire	     				int_intr_error_clear_clr_err_0;
wire	     				int_intr_error_enable_en_err_2;
wire	     				int_intr_error_enable_en_err_1;
wire	     				int_intr_error_enable_en_err_0;
wire	[31:0]				int_intr_h2c_0_h2c;
wire	[31:0]				int_intr_h2c_1_h2c;
wire	[31:0]				int_intr_c2h_0_status_c2h;
wire	[31:0]				int_intr_c2h_1_status_c2h;
wire	[31:0]				int_c2h_gpio_0_status_gpio;
wire	[31:0]				int_c2h_gpio_1_status_gpio;
wire	[31:0]				int_c2h_gpio_2_status_gpio;
wire	[31:0]				int_c2h_gpio_3_status_gpio;
wire	[31:0]				int_c2h_gpio_4_status_gpio;
wire	[31:0]				int_c2h_gpio_5_status_gpio;
wire	[31:0]				int_c2h_gpio_6_status_gpio;
wire	[31:0]				int_c2h_gpio_7_status_gpio;
wire	[31:0]				int_c2h_gpio_8_status_gpio;
wire	[31:0]				int_c2h_gpio_9_status_gpio;
wire	[31:0]				int_c2h_gpio_10_status_gpio;
wire	[31:0]				int_c2h_gpio_11_status_gpio;
wire	[31:0]				int_c2h_gpio_12_status_gpio;
wire	[31:0]				int_c2h_gpio_13_status_gpio;
wire	[31:0]				int_c2h_gpio_14_status_gpio;
wire	[31:0]				int_c2h_gpio_15_status_gpio;
wire	[31:0]				int_addr_in_0_addr;
wire	[31:0]				int_addr_in_1_addr;
wire	[31:0]				int_addr_in_2_addr;
wire	[31:0]				int_addr_in_3_addr;
wire	[31:0]				int_trans_mask_0_addr;
wire	[31:0]				int_trans_mask_1_addr;
wire	[31:0]				int_trans_mask_2_addr;
wire	[31:0]				int_trans_mask_3_addr;
wire	[31:0]				int_trans_addr_0_addr;
wire	[31:0]				int_trans_addr_1_addr;
wire	[31:0]				int_trans_addr_2_addr;
wire	[31:0]				int_trans_addr_3_addr;
wire    [31:0]                          int_resp_order_field;

wire [0:0]	int_desc_0_txn_type_wr_strb;
wire [0:0]	int_desc_0_txn_type_wr_rd;
wire [3:0]	int_desc_0_attr_axregion;
wire [3:0]	int_desc_0_attr_axqos;
wire [2:0]	int_desc_0_attr_axprot;
wire [3:0]	int_desc_0_attr_axcache;
wire [1:0]	int_desc_0_attr_axlock;
wire [1:0]	int_desc_0_attr_axburst;
wire [31:0]	int_desc_0_axid_0_axid;
wire [31:0]	int_desc_0_axid_1_axid;
wire [31:0]	int_desc_0_axid_2_axid;
wire [31:0]	int_desc_0_axid_3_axid;
wire [31:0]	int_desc_0_axuser_0_axuser;
wire [31:0]	int_desc_0_axuser_1_axuser;
wire [31:0]	int_desc_0_axuser_2_axuser;
wire [31:0]	int_desc_0_axuser_3_axuser;
wire [31:0]	int_desc_0_axuser_4_axuser;
wire [31:0]	int_desc_0_axuser_5_axuser;
wire [31:0]	int_desc_0_axuser_6_axuser;
wire [31:0]	int_desc_0_axuser_7_axuser;
wire [31:0]	int_desc_0_axuser_8_axuser;
wire [31:0]	int_desc_0_axuser_9_axuser;
wire [31:0]	int_desc_0_axuser_10_axuser;
wire [31:0]	int_desc_0_axuser_11_axuser;
wire [31:0]	int_desc_0_axuser_12_axuser;
wire [31:0]	int_desc_0_axuser_13_axuser;
wire [31:0]	int_desc_0_axuser_14_axuser;
wire [31:0]	int_desc_0_axuser_15_axuser;
wire [15:0]	int_desc_0_size_txn_size;
wire [2:0]	int_desc_0_axsize_axsize;
wire [31:0]	int_desc_0_axaddr_0_addr;
wire [31:0]	int_desc_0_axaddr_1_addr;
wire [31:0]	int_desc_0_axaddr_2_addr;
wire [31:0]	int_desc_0_axaddr_3_addr;
wire [31:0]	int_desc_0_data_offset_addr;
wire [31:0]	int_desc_0_wuser_0_wuser;
wire [31:0]	int_desc_0_wuser_1_wuser;
wire [31:0]	int_desc_0_wuser_2_wuser;
wire [31:0]	int_desc_0_wuser_3_wuser;
wire [31:0]	int_desc_0_wuser_4_wuser;
wire [31:0]	int_desc_0_wuser_5_wuser;
wire [31:0]	int_desc_0_wuser_6_wuser;
wire [31:0]	int_desc_0_wuser_7_wuser;
wire [31:0]	int_desc_0_wuser_8_wuser;
wire [31:0]	int_desc_0_wuser_9_wuser;
wire [31:0]	int_desc_0_wuser_10_wuser;
wire [31:0]	int_desc_0_wuser_11_wuser;
wire [31:0]	int_desc_0_wuser_12_wuser;
wire [31:0]	int_desc_0_wuser_13_wuser;
wire [31:0]	int_desc_0_wuser_14_wuser;
wire [31:0]	int_desc_0_wuser_15_wuser;
wire [31:0]	int_desc_0_data_host_addr_0_addr;
wire [31:0]	int_desc_0_data_host_addr_1_addr;
wire [31:0]	int_desc_0_data_host_addr_2_addr;
wire [31:0]	int_desc_0_data_host_addr_3_addr;
wire [31:0]	int_desc_0_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_0_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_0_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_0_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_0_xuser_0_xuser;
wire [31:0]	int_desc_0_xuser_1_xuser;
wire [31:0]	int_desc_0_xuser_2_xuser;
wire [31:0]	int_desc_0_xuser_3_xuser;
wire [31:0]	int_desc_0_xuser_4_xuser;
wire [31:0]	int_desc_0_xuser_5_xuser;
wire [31:0]	int_desc_0_xuser_6_xuser;
wire [31:0]	int_desc_0_xuser_7_xuser;
wire [31:0]	int_desc_0_xuser_8_xuser;
wire [31:0]	int_desc_0_xuser_9_xuser;
wire [31:0]	int_desc_0_xuser_10_xuser;
wire [31:0]	int_desc_0_xuser_11_xuser;
wire [31:0]	int_desc_0_xuser_12_xuser;
wire [31:0]	int_desc_0_xuser_13_xuser;
wire [31:0]	int_desc_0_xuser_14_xuser;
wire [31:0]	int_desc_0_xuser_15_xuser;
wire [0:0]	int_desc_1_txn_type_wr_strb;
wire [0:0]	int_desc_1_txn_type_wr_rd;
wire [3:0]	int_desc_1_attr_axregion;
wire [3:0]	int_desc_1_attr_axqos;
wire [2:0]	int_desc_1_attr_axprot;
wire [3:0]	int_desc_1_attr_axcache;
wire [1:0]	int_desc_1_attr_axlock;
wire [1:0]	int_desc_1_attr_axburst;
wire [31:0]	int_desc_1_axid_0_axid;
wire [31:0]	int_desc_1_axid_1_axid;
wire [31:0]	int_desc_1_axid_2_axid;
wire [31:0]	int_desc_1_axid_3_axid;
wire [31:0]	int_desc_1_axuser_0_axuser;
wire [31:0]	int_desc_1_axuser_1_axuser;
wire [31:0]	int_desc_1_axuser_2_axuser;
wire [31:0]	int_desc_1_axuser_3_axuser;
wire [31:0]	int_desc_1_axuser_4_axuser;
wire [31:0]	int_desc_1_axuser_5_axuser;
wire [31:0]	int_desc_1_axuser_6_axuser;
wire [31:0]	int_desc_1_axuser_7_axuser;
wire [31:0]	int_desc_1_axuser_8_axuser;
wire [31:0]	int_desc_1_axuser_9_axuser;
wire [31:0]	int_desc_1_axuser_10_axuser;
wire [31:0]	int_desc_1_axuser_11_axuser;
wire [31:0]	int_desc_1_axuser_12_axuser;
wire [31:0]	int_desc_1_axuser_13_axuser;
wire [31:0]	int_desc_1_axuser_14_axuser;
wire [31:0]	int_desc_1_axuser_15_axuser;
wire [15:0]	int_desc_1_size_txn_size;
wire [2:0]	int_desc_1_axsize_axsize;
wire [31:0]	int_desc_1_axaddr_0_addr;
wire [31:0]	int_desc_1_axaddr_1_addr;
wire [31:0]	int_desc_1_axaddr_2_addr;
wire [31:0]	int_desc_1_axaddr_3_addr;
wire [31:0]	int_desc_1_data_offset_addr;
wire [31:0]	int_desc_1_wuser_0_wuser;
wire [31:0]	int_desc_1_wuser_1_wuser;
wire [31:0]	int_desc_1_wuser_2_wuser;
wire [31:0]	int_desc_1_wuser_3_wuser;
wire [31:0]	int_desc_1_wuser_4_wuser;
wire [31:0]	int_desc_1_wuser_5_wuser;
wire [31:0]	int_desc_1_wuser_6_wuser;
wire [31:0]	int_desc_1_wuser_7_wuser;
wire [31:0]	int_desc_1_wuser_8_wuser;
wire [31:0]	int_desc_1_wuser_9_wuser;
wire [31:0]	int_desc_1_wuser_10_wuser;
wire [31:0]	int_desc_1_wuser_11_wuser;
wire [31:0]	int_desc_1_wuser_12_wuser;
wire [31:0]	int_desc_1_wuser_13_wuser;
wire [31:0]	int_desc_1_wuser_14_wuser;
wire [31:0]	int_desc_1_wuser_15_wuser;
wire [31:0]	int_desc_1_data_host_addr_0_addr;
wire [31:0]	int_desc_1_data_host_addr_1_addr;
wire [31:0]	int_desc_1_data_host_addr_2_addr;
wire [31:0]	int_desc_1_data_host_addr_3_addr;
wire [31:0]	int_desc_1_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_1_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_1_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_1_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_1_xuser_0_xuser;
wire [31:0]	int_desc_1_xuser_1_xuser;
wire [31:0]	int_desc_1_xuser_2_xuser;
wire [31:0]	int_desc_1_xuser_3_xuser;
wire [31:0]	int_desc_1_xuser_4_xuser;
wire [31:0]	int_desc_1_xuser_5_xuser;
wire [31:0]	int_desc_1_xuser_6_xuser;
wire [31:0]	int_desc_1_xuser_7_xuser;
wire [31:0]	int_desc_1_xuser_8_xuser;
wire [31:0]	int_desc_1_xuser_9_xuser;
wire [31:0]	int_desc_1_xuser_10_xuser;
wire [31:0]	int_desc_1_xuser_11_xuser;
wire [31:0]	int_desc_1_xuser_12_xuser;
wire [31:0]	int_desc_1_xuser_13_xuser;
wire [31:0]	int_desc_1_xuser_14_xuser;
wire [31:0]	int_desc_1_xuser_15_xuser;
wire [0:0]	int_desc_2_txn_type_wr_strb;
wire [0:0]	int_desc_2_txn_type_wr_rd;
wire [3:0]	int_desc_2_attr_axregion;
wire [3:0]	int_desc_2_attr_axqos;
wire [2:0]	int_desc_2_attr_axprot;
wire [3:0]	int_desc_2_attr_axcache;
wire [1:0]	int_desc_2_attr_axlock;
wire [1:0]	int_desc_2_attr_axburst;
wire [31:0]	int_desc_2_axid_0_axid;
wire [31:0]	int_desc_2_axid_1_axid;
wire [31:0]	int_desc_2_axid_2_axid;
wire [31:0]	int_desc_2_axid_3_axid;
wire [31:0]	int_desc_2_axuser_0_axuser;
wire [31:0]	int_desc_2_axuser_1_axuser;
wire [31:0]	int_desc_2_axuser_2_axuser;
wire [31:0]	int_desc_2_axuser_3_axuser;
wire [31:0]	int_desc_2_axuser_4_axuser;
wire [31:0]	int_desc_2_axuser_5_axuser;
wire [31:0]	int_desc_2_axuser_6_axuser;
wire [31:0]	int_desc_2_axuser_7_axuser;
wire [31:0]	int_desc_2_axuser_8_axuser;
wire [31:0]	int_desc_2_axuser_9_axuser;
wire [31:0]	int_desc_2_axuser_10_axuser;
wire [31:0]	int_desc_2_axuser_11_axuser;
wire [31:0]	int_desc_2_axuser_12_axuser;
wire [31:0]	int_desc_2_axuser_13_axuser;
wire [31:0]	int_desc_2_axuser_14_axuser;
wire [31:0]	int_desc_2_axuser_15_axuser;
wire [15:0]	int_desc_2_size_txn_size;
wire [2:0]	int_desc_2_axsize_axsize;
wire [31:0]	int_desc_2_axaddr_0_addr;
wire [31:0]	int_desc_2_axaddr_1_addr;
wire [31:0]	int_desc_2_axaddr_2_addr;
wire [31:0]	int_desc_2_axaddr_3_addr;
wire [31:0]	int_desc_2_data_offset_addr;
wire [31:0]	int_desc_2_wuser_0_wuser;
wire [31:0]	int_desc_2_wuser_1_wuser;
wire [31:0]	int_desc_2_wuser_2_wuser;
wire [31:0]	int_desc_2_wuser_3_wuser;
wire [31:0]	int_desc_2_wuser_4_wuser;
wire [31:0]	int_desc_2_wuser_5_wuser;
wire [31:0]	int_desc_2_wuser_6_wuser;
wire [31:0]	int_desc_2_wuser_7_wuser;
wire [31:0]	int_desc_2_wuser_8_wuser;
wire [31:0]	int_desc_2_wuser_9_wuser;
wire [31:0]	int_desc_2_wuser_10_wuser;
wire [31:0]	int_desc_2_wuser_11_wuser;
wire [31:0]	int_desc_2_wuser_12_wuser;
wire [31:0]	int_desc_2_wuser_13_wuser;
wire [31:0]	int_desc_2_wuser_14_wuser;
wire [31:0]	int_desc_2_wuser_15_wuser;
wire [31:0]	int_desc_2_data_host_addr_0_addr;
wire [31:0]	int_desc_2_data_host_addr_1_addr;
wire [31:0]	int_desc_2_data_host_addr_2_addr;
wire [31:0]	int_desc_2_data_host_addr_3_addr;
wire [31:0]	int_desc_2_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_2_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_2_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_2_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_2_xuser_0_xuser;
wire [31:0]	int_desc_2_xuser_1_xuser;
wire [31:0]	int_desc_2_xuser_2_xuser;
wire [31:0]	int_desc_2_xuser_3_xuser;
wire [31:0]	int_desc_2_xuser_4_xuser;
wire [31:0]	int_desc_2_xuser_5_xuser;
wire [31:0]	int_desc_2_xuser_6_xuser;
wire [31:0]	int_desc_2_xuser_7_xuser;
wire [31:0]	int_desc_2_xuser_8_xuser;
wire [31:0]	int_desc_2_xuser_9_xuser;
wire [31:0]	int_desc_2_xuser_10_xuser;
wire [31:0]	int_desc_2_xuser_11_xuser;
wire [31:0]	int_desc_2_xuser_12_xuser;
wire [31:0]	int_desc_2_xuser_13_xuser;
wire [31:0]	int_desc_2_xuser_14_xuser;
wire [31:0]	int_desc_2_xuser_15_xuser;
wire [0:0]	int_desc_3_txn_type_wr_strb;
wire [0:0]	int_desc_3_txn_type_wr_rd;
wire [3:0]	int_desc_3_attr_axregion;
wire [3:0]	int_desc_3_attr_axqos;
wire [2:0]	int_desc_3_attr_axprot;
wire [3:0]	int_desc_3_attr_axcache;
wire [1:0]	int_desc_3_attr_axlock;
wire [1:0]	int_desc_3_attr_axburst;
wire [31:0]	int_desc_3_axid_0_axid;
wire [31:0]	int_desc_3_axid_1_axid;
wire [31:0]	int_desc_3_axid_2_axid;
wire [31:0]	int_desc_3_axid_3_axid;
wire [31:0]	int_desc_3_axuser_0_axuser;
wire [31:0]	int_desc_3_axuser_1_axuser;
wire [31:0]	int_desc_3_axuser_2_axuser;
wire [31:0]	int_desc_3_axuser_3_axuser;
wire [31:0]	int_desc_3_axuser_4_axuser;
wire [31:0]	int_desc_3_axuser_5_axuser;
wire [31:0]	int_desc_3_axuser_6_axuser;
wire [31:0]	int_desc_3_axuser_7_axuser;
wire [31:0]	int_desc_3_axuser_8_axuser;
wire [31:0]	int_desc_3_axuser_9_axuser;
wire [31:0]	int_desc_3_axuser_10_axuser;
wire [31:0]	int_desc_3_axuser_11_axuser;
wire [31:0]	int_desc_3_axuser_12_axuser;
wire [31:0]	int_desc_3_axuser_13_axuser;
wire [31:0]	int_desc_3_axuser_14_axuser;
wire [31:0]	int_desc_3_axuser_15_axuser;
wire [15:0]	int_desc_3_size_txn_size;
wire [2:0]	int_desc_3_axsize_axsize;
wire [31:0]	int_desc_3_axaddr_0_addr;
wire [31:0]	int_desc_3_axaddr_1_addr;
wire [31:0]	int_desc_3_axaddr_2_addr;
wire [31:0]	int_desc_3_axaddr_3_addr;
wire [31:0]	int_desc_3_data_offset_addr;
wire [31:0]	int_desc_3_wuser_0_wuser;
wire [31:0]	int_desc_3_wuser_1_wuser;
wire [31:0]	int_desc_3_wuser_2_wuser;
wire [31:0]	int_desc_3_wuser_3_wuser;
wire [31:0]	int_desc_3_wuser_4_wuser;
wire [31:0]	int_desc_3_wuser_5_wuser;
wire [31:0]	int_desc_3_wuser_6_wuser;
wire [31:0]	int_desc_3_wuser_7_wuser;
wire [31:0]	int_desc_3_wuser_8_wuser;
wire [31:0]	int_desc_3_wuser_9_wuser;
wire [31:0]	int_desc_3_wuser_10_wuser;
wire [31:0]	int_desc_3_wuser_11_wuser;
wire [31:0]	int_desc_3_wuser_12_wuser;
wire [31:0]	int_desc_3_wuser_13_wuser;
wire [31:0]	int_desc_3_wuser_14_wuser;
wire [31:0]	int_desc_3_wuser_15_wuser;
wire [31:0]	int_desc_3_data_host_addr_0_addr;
wire [31:0]	int_desc_3_data_host_addr_1_addr;
wire [31:0]	int_desc_3_data_host_addr_2_addr;
wire [31:0]	int_desc_3_data_host_addr_3_addr;
wire [31:0]	int_desc_3_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_3_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_3_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_3_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_3_xuser_0_xuser;
wire [31:0]	int_desc_3_xuser_1_xuser;
wire [31:0]	int_desc_3_xuser_2_xuser;
wire [31:0]	int_desc_3_xuser_3_xuser;
wire [31:0]	int_desc_3_xuser_4_xuser;
wire [31:0]	int_desc_3_xuser_5_xuser;
wire [31:0]	int_desc_3_xuser_6_xuser;
wire [31:0]	int_desc_3_xuser_7_xuser;
wire [31:0]	int_desc_3_xuser_8_xuser;
wire [31:0]	int_desc_3_xuser_9_xuser;
wire [31:0]	int_desc_3_xuser_10_xuser;
wire [31:0]	int_desc_3_xuser_11_xuser;
wire [31:0]	int_desc_3_xuser_12_xuser;
wire [31:0]	int_desc_3_xuser_13_xuser;
wire [31:0]	int_desc_3_xuser_14_xuser;
wire [31:0]	int_desc_3_xuser_15_xuser;
wire [0:0]	int_desc_4_txn_type_wr_strb;
wire [0:0]	int_desc_4_txn_type_wr_rd;
wire [3:0]	int_desc_4_attr_axregion;
wire [3:0]	int_desc_4_attr_axqos;
wire [2:0]	int_desc_4_attr_axprot;
wire [3:0]	int_desc_4_attr_axcache;
wire [1:0]	int_desc_4_attr_axlock;
wire [1:0]	int_desc_4_attr_axburst;
wire [31:0]	int_desc_4_axid_0_axid;
wire [31:0]	int_desc_4_axid_1_axid;
wire [31:0]	int_desc_4_axid_2_axid;
wire [31:0]	int_desc_4_axid_3_axid;
wire [31:0]	int_desc_4_axuser_0_axuser;
wire [31:0]	int_desc_4_axuser_1_axuser;
wire [31:0]	int_desc_4_axuser_2_axuser;
wire [31:0]	int_desc_4_axuser_3_axuser;
wire [31:0]	int_desc_4_axuser_4_axuser;
wire [31:0]	int_desc_4_axuser_5_axuser;
wire [31:0]	int_desc_4_axuser_6_axuser;
wire [31:0]	int_desc_4_axuser_7_axuser;
wire [31:0]	int_desc_4_axuser_8_axuser;
wire [31:0]	int_desc_4_axuser_9_axuser;
wire [31:0]	int_desc_4_axuser_10_axuser;
wire [31:0]	int_desc_4_axuser_11_axuser;
wire [31:0]	int_desc_4_axuser_12_axuser;
wire [31:0]	int_desc_4_axuser_13_axuser;
wire [31:0]	int_desc_4_axuser_14_axuser;
wire [31:0]	int_desc_4_axuser_15_axuser;
wire [15:0]	int_desc_4_size_txn_size;
wire [2:0]	int_desc_4_axsize_axsize;
wire [31:0]	int_desc_4_axaddr_0_addr;
wire [31:0]	int_desc_4_axaddr_1_addr;
wire [31:0]	int_desc_4_axaddr_2_addr;
wire [31:0]	int_desc_4_axaddr_3_addr;
wire [31:0]	int_desc_4_data_offset_addr;
wire [31:0]	int_desc_4_wuser_0_wuser;
wire [31:0]	int_desc_4_wuser_1_wuser;
wire [31:0]	int_desc_4_wuser_2_wuser;
wire [31:0]	int_desc_4_wuser_3_wuser;
wire [31:0]	int_desc_4_wuser_4_wuser;
wire [31:0]	int_desc_4_wuser_5_wuser;
wire [31:0]	int_desc_4_wuser_6_wuser;
wire [31:0]	int_desc_4_wuser_7_wuser;
wire [31:0]	int_desc_4_wuser_8_wuser;
wire [31:0]	int_desc_4_wuser_9_wuser;
wire [31:0]	int_desc_4_wuser_10_wuser;
wire [31:0]	int_desc_4_wuser_11_wuser;
wire [31:0]	int_desc_4_wuser_12_wuser;
wire [31:0]	int_desc_4_wuser_13_wuser;
wire [31:0]	int_desc_4_wuser_14_wuser;
wire [31:0]	int_desc_4_wuser_15_wuser;
wire [31:0]	int_desc_4_data_host_addr_0_addr;
wire [31:0]	int_desc_4_data_host_addr_1_addr;
wire [31:0]	int_desc_4_data_host_addr_2_addr;
wire [31:0]	int_desc_4_data_host_addr_3_addr;
wire [31:0]	int_desc_4_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_4_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_4_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_4_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_4_xuser_0_xuser;
wire [31:0]	int_desc_4_xuser_1_xuser;
wire [31:0]	int_desc_4_xuser_2_xuser;
wire [31:0]	int_desc_4_xuser_3_xuser;
wire [31:0]	int_desc_4_xuser_4_xuser;
wire [31:0]	int_desc_4_xuser_5_xuser;
wire [31:0]	int_desc_4_xuser_6_xuser;
wire [31:0]	int_desc_4_xuser_7_xuser;
wire [31:0]	int_desc_4_xuser_8_xuser;
wire [31:0]	int_desc_4_xuser_9_xuser;
wire [31:0]	int_desc_4_xuser_10_xuser;
wire [31:0]	int_desc_4_xuser_11_xuser;
wire [31:0]	int_desc_4_xuser_12_xuser;
wire [31:0]	int_desc_4_xuser_13_xuser;
wire [31:0]	int_desc_4_xuser_14_xuser;
wire [31:0]	int_desc_4_xuser_15_xuser;
wire [0:0]	int_desc_5_txn_type_wr_strb;
wire [0:0]	int_desc_5_txn_type_wr_rd;
wire [3:0]	int_desc_5_attr_axregion;
wire [3:0]	int_desc_5_attr_axqos;
wire [2:0]	int_desc_5_attr_axprot;
wire [3:0]	int_desc_5_attr_axcache;
wire [1:0]	int_desc_5_attr_axlock;
wire [1:0]	int_desc_5_attr_axburst;
wire [31:0]	int_desc_5_axid_0_axid;
wire [31:0]	int_desc_5_axid_1_axid;
wire [31:0]	int_desc_5_axid_2_axid;
wire [31:0]	int_desc_5_axid_3_axid;
wire [31:0]	int_desc_5_axuser_0_axuser;
wire [31:0]	int_desc_5_axuser_1_axuser;
wire [31:0]	int_desc_5_axuser_2_axuser;
wire [31:0]	int_desc_5_axuser_3_axuser;
wire [31:0]	int_desc_5_axuser_4_axuser;
wire [31:0]	int_desc_5_axuser_5_axuser;
wire [31:0]	int_desc_5_axuser_6_axuser;
wire [31:0]	int_desc_5_axuser_7_axuser;
wire [31:0]	int_desc_5_axuser_8_axuser;
wire [31:0]	int_desc_5_axuser_9_axuser;
wire [31:0]	int_desc_5_axuser_10_axuser;
wire [31:0]	int_desc_5_axuser_11_axuser;
wire [31:0]	int_desc_5_axuser_12_axuser;
wire [31:0]	int_desc_5_axuser_13_axuser;
wire [31:0]	int_desc_5_axuser_14_axuser;
wire [31:0]	int_desc_5_axuser_15_axuser;
wire [15:0]	int_desc_5_size_txn_size;
wire [2:0]	int_desc_5_axsize_axsize;
wire [31:0]	int_desc_5_axaddr_0_addr;
wire [31:0]	int_desc_5_axaddr_1_addr;
wire [31:0]	int_desc_5_axaddr_2_addr;
wire [31:0]	int_desc_5_axaddr_3_addr;
wire [31:0]	int_desc_5_data_offset_addr;
wire [31:0]	int_desc_5_wuser_0_wuser;
wire [31:0]	int_desc_5_wuser_1_wuser;
wire [31:0]	int_desc_5_wuser_2_wuser;
wire [31:0]	int_desc_5_wuser_3_wuser;
wire [31:0]	int_desc_5_wuser_4_wuser;
wire [31:0]	int_desc_5_wuser_5_wuser;
wire [31:0]	int_desc_5_wuser_6_wuser;
wire [31:0]	int_desc_5_wuser_7_wuser;
wire [31:0]	int_desc_5_wuser_8_wuser;
wire [31:0]	int_desc_5_wuser_9_wuser;
wire [31:0]	int_desc_5_wuser_10_wuser;
wire [31:0]	int_desc_5_wuser_11_wuser;
wire [31:0]	int_desc_5_wuser_12_wuser;
wire [31:0]	int_desc_5_wuser_13_wuser;
wire [31:0]	int_desc_5_wuser_14_wuser;
wire [31:0]	int_desc_5_wuser_15_wuser;
wire [31:0]	int_desc_5_data_host_addr_0_addr;
wire [31:0]	int_desc_5_data_host_addr_1_addr;
wire [31:0]	int_desc_5_data_host_addr_2_addr;
wire [31:0]	int_desc_5_data_host_addr_3_addr;
wire [31:0]	int_desc_5_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_5_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_5_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_5_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_5_xuser_0_xuser;
wire [31:0]	int_desc_5_xuser_1_xuser;
wire [31:0]	int_desc_5_xuser_2_xuser;
wire [31:0]	int_desc_5_xuser_3_xuser;
wire [31:0]	int_desc_5_xuser_4_xuser;
wire [31:0]	int_desc_5_xuser_5_xuser;
wire [31:0]	int_desc_5_xuser_6_xuser;
wire [31:0]	int_desc_5_xuser_7_xuser;
wire [31:0]	int_desc_5_xuser_8_xuser;
wire [31:0]	int_desc_5_xuser_9_xuser;
wire [31:0]	int_desc_5_xuser_10_xuser;
wire [31:0]	int_desc_5_xuser_11_xuser;
wire [31:0]	int_desc_5_xuser_12_xuser;
wire [31:0]	int_desc_5_xuser_13_xuser;
wire [31:0]	int_desc_5_xuser_14_xuser;
wire [31:0]	int_desc_5_xuser_15_xuser;
wire [0:0]	int_desc_6_txn_type_wr_strb;
wire [0:0]	int_desc_6_txn_type_wr_rd;
wire [3:0]	int_desc_6_attr_axregion;
wire [3:0]	int_desc_6_attr_axqos;
wire [2:0]	int_desc_6_attr_axprot;
wire [3:0]	int_desc_6_attr_axcache;
wire [1:0]	int_desc_6_attr_axlock;
wire [1:0]	int_desc_6_attr_axburst;
wire [31:0]	int_desc_6_axid_0_axid;
wire [31:0]	int_desc_6_axid_1_axid;
wire [31:0]	int_desc_6_axid_2_axid;
wire [31:0]	int_desc_6_axid_3_axid;
wire [31:0]	int_desc_6_axuser_0_axuser;
wire [31:0]	int_desc_6_axuser_1_axuser;
wire [31:0]	int_desc_6_axuser_2_axuser;
wire [31:0]	int_desc_6_axuser_3_axuser;
wire [31:0]	int_desc_6_axuser_4_axuser;
wire [31:0]	int_desc_6_axuser_5_axuser;
wire [31:0]	int_desc_6_axuser_6_axuser;
wire [31:0]	int_desc_6_axuser_7_axuser;
wire [31:0]	int_desc_6_axuser_8_axuser;
wire [31:0]	int_desc_6_axuser_9_axuser;
wire [31:0]	int_desc_6_axuser_10_axuser;
wire [31:0]	int_desc_6_axuser_11_axuser;
wire [31:0]	int_desc_6_axuser_12_axuser;
wire [31:0]	int_desc_6_axuser_13_axuser;
wire [31:0]	int_desc_6_axuser_14_axuser;
wire [31:0]	int_desc_6_axuser_15_axuser;
wire [15:0]	int_desc_6_size_txn_size;
wire [2:0]	int_desc_6_axsize_axsize;
wire [31:0]	int_desc_6_axaddr_0_addr;
wire [31:0]	int_desc_6_axaddr_1_addr;
wire [31:0]	int_desc_6_axaddr_2_addr;
wire [31:0]	int_desc_6_axaddr_3_addr;
wire [31:0]	int_desc_6_data_offset_addr;
wire [31:0]	int_desc_6_wuser_0_wuser;
wire [31:0]	int_desc_6_wuser_1_wuser;
wire [31:0]	int_desc_6_wuser_2_wuser;
wire [31:0]	int_desc_6_wuser_3_wuser;
wire [31:0]	int_desc_6_wuser_4_wuser;
wire [31:0]	int_desc_6_wuser_5_wuser;
wire [31:0]	int_desc_6_wuser_6_wuser;
wire [31:0]	int_desc_6_wuser_7_wuser;
wire [31:0]	int_desc_6_wuser_8_wuser;
wire [31:0]	int_desc_6_wuser_9_wuser;
wire [31:0]	int_desc_6_wuser_10_wuser;
wire [31:0]	int_desc_6_wuser_11_wuser;
wire [31:0]	int_desc_6_wuser_12_wuser;
wire [31:0]	int_desc_6_wuser_13_wuser;
wire [31:0]	int_desc_6_wuser_14_wuser;
wire [31:0]	int_desc_6_wuser_15_wuser;
wire [31:0]	int_desc_6_data_host_addr_0_addr;
wire [31:0]	int_desc_6_data_host_addr_1_addr;
wire [31:0]	int_desc_6_data_host_addr_2_addr;
wire [31:0]	int_desc_6_data_host_addr_3_addr;
wire [31:0]	int_desc_6_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_6_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_6_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_6_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_6_xuser_0_xuser;
wire [31:0]	int_desc_6_xuser_1_xuser;
wire [31:0]	int_desc_6_xuser_2_xuser;
wire [31:0]	int_desc_6_xuser_3_xuser;
wire [31:0]	int_desc_6_xuser_4_xuser;
wire [31:0]	int_desc_6_xuser_5_xuser;
wire [31:0]	int_desc_6_xuser_6_xuser;
wire [31:0]	int_desc_6_xuser_7_xuser;
wire [31:0]	int_desc_6_xuser_8_xuser;
wire [31:0]	int_desc_6_xuser_9_xuser;
wire [31:0]	int_desc_6_xuser_10_xuser;
wire [31:0]	int_desc_6_xuser_11_xuser;
wire [31:0]	int_desc_6_xuser_12_xuser;
wire [31:0]	int_desc_6_xuser_13_xuser;
wire [31:0]	int_desc_6_xuser_14_xuser;
wire [31:0]	int_desc_6_xuser_15_xuser;
wire [0:0]	int_desc_7_txn_type_wr_strb;
wire [0:0]	int_desc_7_txn_type_wr_rd;
wire [3:0]	int_desc_7_attr_axregion;
wire [3:0]	int_desc_7_attr_axqos;
wire [2:0]	int_desc_7_attr_axprot;
wire [3:0]	int_desc_7_attr_axcache;
wire [1:0]	int_desc_7_attr_axlock;
wire [1:0]	int_desc_7_attr_axburst;
wire [31:0]	int_desc_7_axid_0_axid;
wire [31:0]	int_desc_7_axid_1_axid;
wire [31:0]	int_desc_7_axid_2_axid;
wire [31:0]	int_desc_7_axid_3_axid;
wire [31:0]	int_desc_7_axuser_0_axuser;
wire [31:0]	int_desc_7_axuser_1_axuser;
wire [31:0]	int_desc_7_axuser_2_axuser;
wire [31:0]	int_desc_7_axuser_3_axuser;
wire [31:0]	int_desc_7_axuser_4_axuser;
wire [31:0]	int_desc_7_axuser_5_axuser;
wire [31:0]	int_desc_7_axuser_6_axuser;
wire [31:0]	int_desc_7_axuser_7_axuser;
wire [31:0]	int_desc_7_axuser_8_axuser;
wire [31:0]	int_desc_7_axuser_9_axuser;
wire [31:0]	int_desc_7_axuser_10_axuser;
wire [31:0]	int_desc_7_axuser_11_axuser;
wire [31:0]	int_desc_7_axuser_12_axuser;
wire [31:0]	int_desc_7_axuser_13_axuser;
wire [31:0]	int_desc_7_axuser_14_axuser;
wire [31:0]	int_desc_7_axuser_15_axuser;
wire [15:0]	int_desc_7_size_txn_size;
wire [2:0]	int_desc_7_axsize_axsize;
wire [31:0]	int_desc_7_axaddr_0_addr;
wire [31:0]	int_desc_7_axaddr_1_addr;
wire [31:0]	int_desc_7_axaddr_2_addr;
wire [31:0]	int_desc_7_axaddr_3_addr;
wire [31:0]	int_desc_7_data_offset_addr;
wire [31:0]	int_desc_7_wuser_0_wuser;
wire [31:0]	int_desc_7_wuser_1_wuser;
wire [31:0]	int_desc_7_wuser_2_wuser;
wire [31:0]	int_desc_7_wuser_3_wuser;
wire [31:0]	int_desc_7_wuser_4_wuser;
wire [31:0]	int_desc_7_wuser_5_wuser;
wire [31:0]	int_desc_7_wuser_6_wuser;
wire [31:0]	int_desc_7_wuser_7_wuser;
wire [31:0]	int_desc_7_wuser_8_wuser;
wire [31:0]	int_desc_7_wuser_9_wuser;
wire [31:0]	int_desc_7_wuser_10_wuser;
wire [31:0]	int_desc_7_wuser_11_wuser;
wire [31:0]	int_desc_7_wuser_12_wuser;
wire [31:0]	int_desc_7_wuser_13_wuser;
wire [31:0]	int_desc_7_wuser_14_wuser;
wire [31:0]	int_desc_7_wuser_15_wuser;
wire [31:0]	int_desc_7_data_host_addr_0_addr;
wire [31:0]	int_desc_7_data_host_addr_1_addr;
wire [31:0]	int_desc_7_data_host_addr_2_addr;
wire [31:0]	int_desc_7_data_host_addr_3_addr;
wire [31:0]	int_desc_7_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_7_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_7_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_7_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_7_xuser_0_xuser;
wire [31:0]	int_desc_7_xuser_1_xuser;
wire [31:0]	int_desc_7_xuser_2_xuser;
wire [31:0]	int_desc_7_xuser_3_xuser;
wire [31:0]	int_desc_7_xuser_4_xuser;
wire [31:0]	int_desc_7_xuser_5_xuser;
wire [31:0]	int_desc_7_xuser_6_xuser;
wire [31:0]	int_desc_7_xuser_7_xuser;
wire [31:0]	int_desc_7_xuser_8_xuser;
wire [31:0]	int_desc_7_xuser_9_xuser;
wire [31:0]	int_desc_7_xuser_10_xuser;
wire [31:0]	int_desc_7_xuser_11_xuser;
wire [31:0]	int_desc_7_xuser_12_xuser;
wire [31:0]	int_desc_7_xuser_13_xuser;
wire [31:0]	int_desc_7_xuser_14_xuser;
wire [31:0]	int_desc_7_xuser_15_xuser;
wire [0:0]	int_desc_8_txn_type_wr_strb;
wire [0:0]	int_desc_8_txn_type_wr_rd;
wire [3:0]	int_desc_8_attr_axregion;
wire [3:0]	int_desc_8_attr_axqos;
wire [2:0]	int_desc_8_attr_axprot;
wire [3:0]	int_desc_8_attr_axcache;
wire [1:0]	int_desc_8_attr_axlock;
wire [1:0]	int_desc_8_attr_axburst;
wire [31:0]	int_desc_8_axid_0_axid;
wire [31:0]	int_desc_8_axid_1_axid;
wire [31:0]	int_desc_8_axid_2_axid;
wire [31:0]	int_desc_8_axid_3_axid;
wire [31:0]	int_desc_8_axuser_0_axuser;
wire [31:0]	int_desc_8_axuser_1_axuser;
wire [31:0]	int_desc_8_axuser_2_axuser;
wire [31:0]	int_desc_8_axuser_3_axuser;
wire [31:0]	int_desc_8_axuser_4_axuser;
wire [31:0]	int_desc_8_axuser_5_axuser;
wire [31:0]	int_desc_8_axuser_6_axuser;
wire [31:0]	int_desc_8_axuser_7_axuser;
wire [31:0]	int_desc_8_axuser_8_axuser;
wire [31:0]	int_desc_8_axuser_9_axuser;
wire [31:0]	int_desc_8_axuser_10_axuser;
wire [31:0]	int_desc_8_axuser_11_axuser;
wire [31:0]	int_desc_8_axuser_12_axuser;
wire [31:0]	int_desc_8_axuser_13_axuser;
wire [31:0]	int_desc_8_axuser_14_axuser;
wire [31:0]	int_desc_8_axuser_15_axuser;
wire [15:0]	int_desc_8_size_txn_size;
wire [2:0]	int_desc_8_axsize_axsize;
wire [31:0]	int_desc_8_axaddr_0_addr;
wire [31:0]	int_desc_8_axaddr_1_addr;
wire [31:0]	int_desc_8_axaddr_2_addr;
wire [31:0]	int_desc_8_axaddr_3_addr;
wire [31:0]	int_desc_8_data_offset_addr;
wire [31:0]	int_desc_8_wuser_0_wuser;
wire [31:0]	int_desc_8_wuser_1_wuser;
wire [31:0]	int_desc_8_wuser_2_wuser;
wire [31:0]	int_desc_8_wuser_3_wuser;
wire [31:0]	int_desc_8_wuser_4_wuser;
wire [31:0]	int_desc_8_wuser_5_wuser;
wire [31:0]	int_desc_8_wuser_6_wuser;
wire [31:0]	int_desc_8_wuser_7_wuser;
wire [31:0]	int_desc_8_wuser_8_wuser;
wire [31:0]	int_desc_8_wuser_9_wuser;
wire [31:0]	int_desc_8_wuser_10_wuser;
wire [31:0]	int_desc_8_wuser_11_wuser;
wire [31:0]	int_desc_8_wuser_12_wuser;
wire [31:0]	int_desc_8_wuser_13_wuser;
wire [31:0]	int_desc_8_wuser_14_wuser;
wire [31:0]	int_desc_8_wuser_15_wuser;
wire [31:0]	int_desc_8_data_host_addr_0_addr;
wire [31:0]	int_desc_8_data_host_addr_1_addr;
wire [31:0]	int_desc_8_data_host_addr_2_addr;
wire [31:0]	int_desc_8_data_host_addr_3_addr;
wire [31:0]	int_desc_8_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_8_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_8_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_8_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_8_xuser_0_xuser;
wire [31:0]	int_desc_8_xuser_1_xuser;
wire [31:0]	int_desc_8_xuser_2_xuser;
wire [31:0]	int_desc_8_xuser_3_xuser;
wire [31:0]	int_desc_8_xuser_4_xuser;
wire [31:0]	int_desc_8_xuser_5_xuser;
wire [31:0]	int_desc_8_xuser_6_xuser;
wire [31:0]	int_desc_8_xuser_7_xuser;
wire [31:0]	int_desc_8_xuser_8_xuser;
wire [31:0]	int_desc_8_xuser_9_xuser;
wire [31:0]	int_desc_8_xuser_10_xuser;
wire [31:0]	int_desc_8_xuser_11_xuser;
wire [31:0]	int_desc_8_xuser_12_xuser;
wire [31:0]	int_desc_8_xuser_13_xuser;
wire [31:0]	int_desc_8_xuser_14_xuser;
wire [31:0]	int_desc_8_xuser_15_xuser;
wire [0:0]	int_desc_9_txn_type_wr_strb;
wire [0:0]	int_desc_9_txn_type_wr_rd;
wire [3:0]	int_desc_9_attr_axregion;
wire [3:0]	int_desc_9_attr_axqos;
wire [2:0]	int_desc_9_attr_axprot;
wire [3:0]	int_desc_9_attr_axcache;
wire [1:0]	int_desc_9_attr_axlock;
wire [1:0]	int_desc_9_attr_axburst;
wire [31:0]	int_desc_9_axid_0_axid;
wire [31:0]	int_desc_9_axid_1_axid;
wire [31:0]	int_desc_9_axid_2_axid;
wire [31:0]	int_desc_9_axid_3_axid;
wire [31:0]	int_desc_9_axuser_0_axuser;
wire [31:0]	int_desc_9_axuser_1_axuser;
wire [31:0]	int_desc_9_axuser_2_axuser;
wire [31:0]	int_desc_9_axuser_3_axuser;
wire [31:0]	int_desc_9_axuser_4_axuser;
wire [31:0]	int_desc_9_axuser_5_axuser;
wire [31:0]	int_desc_9_axuser_6_axuser;
wire [31:0]	int_desc_9_axuser_7_axuser;
wire [31:0]	int_desc_9_axuser_8_axuser;
wire [31:0]	int_desc_9_axuser_9_axuser;
wire [31:0]	int_desc_9_axuser_10_axuser;
wire [31:0]	int_desc_9_axuser_11_axuser;
wire [31:0]	int_desc_9_axuser_12_axuser;
wire [31:0]	int_desc_9_axuser_13_axuser;
wire [31:0]	int_desc_9_axuser_14_axuser;
wire [31:0]	int_desc_9_axuser_15_axuser;
wire [15:0]	int_desc_9_size_txn_size;
wire [2:0]	int_desc_9_axsize_axsize;
wire [31:0]	int_desc_9_axaddr_0_addr;
wire [31:0]	int_desc_9_axaddr_1_addr;
wire [31:0]	int_desc_9_axaddr_2_addr;
wire [31:0]	int_desc_9_axaddr_3_addr;
wire [31:0]	int_desc_9_data_offset_addr;
wire [31:0]	int_desc_9_wuser_0_wuser;
wire [31:0]	int_desc_9_wuser_1_wuser;
wire [31:0]	int_desc_9_wuser_2_wuser;
wire [31:0]	int_desc_9_wuser_3_wuser;
wire [31:0]	int_desc_9_wuser_4_wuser;
wire [31:0]	int_desc_9_wuser_5_wuser;
wire [31:0]	int_desc_9_wuser_6_wuser;
wire [31:0]	int_desc_9_wuser_7_wuser;
wire [31:0]	int_desc_9_wuser_8_wuser;
wire [31:0]	int_desc_9_wuser_9_wuser;
wire [31:0]	int_desc_9_wuser_10_wuser;
wire [31:0]	int_desc_9_wuser_11_wuser;
wire [31:0]	int_desc_9_wuser_12_wuser;
wire [31:0]	int_desc_9_wuser_13_wuser;
wire [31:0]	int_desc_9_wuser_14_wuser;
wire [31:0]	int_desc_9_wuser_15_wuser;
wire [31:0]	int_desc_9_data_host_addr_0_addr;
wire [31:0]	int_desc_9_data_host_addr_1_addr;
wire [31:0]	int_desc_9_data_host_addr_2_addr;
wire [31:0]	int_desc_9_data_host_addr_3_addr;
wire [31:0]	int_desc_9_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_9_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_9_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_9_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_9_xuser_0_xuser;
wire [31:0]	int_desc_9_xuser_1_xuser;
wire [31:0]	int_desc_9_xuser_2_xuser;
wire [31:0]	int_desc_9_xuser_3_xuser;
wire [31:0]	int_desc_9_xuser_4_xuser;
wire [31:0]	int_desc_9_xuser_5_xuser;
wire [31:0]	int_desc_9_xuser_6_xuser;
wire [31:0]	int_desc_9_xuser_7_xuser;
wire [31:0]	int_desc_9_xuser_8_xuser;
wire [31:0]	int_desc_9_xuser_9_xuser;
wire [31:0]	int_desc_9_xuser_10_xuser;
wire [31:0]	int_desc_9_xuser_11_xuser;
wire [31:0]	int_desc_9_xuser_12_xuser;
wire [31:0]	int_desc_9_xuser_13_xuser;
wire [31:0]	int_desc_9_xuser_14_xuser;
wire [31:0]	int_desc_9_xuser_15_xuser;
wire [0:0]	int_desc_10_txn_type_wr_strb;
wire [0:0]	int_desc_10_txn_type_wr_rd;
wire [3:0]	int_desc_10_attr_axregion;
wire [3:0]	int_desc_10_attr_axqos;
wire [2:0]	int_desc_10_attr_axprot;
wire [3:0]	int_desc_10_attr_axcache;
wire [1:0]	int_desc_10_attr_axlock;
wire [1:0]	int_desc_10_attr_axburst;
wire [31:0]	int_desc_10_axid_0_axid;
wire [31:0]	int_desc_10_axid_1_axid;
wire [31:0]	int_desc_10_axid_2_axid;
wire [31:0]	int_desc_10_axid_3_axid;
wire [31:0]	int_desc_10_axuser_0_axuser;
wire [31:0]	int_desc_10_axuser_1_axuser;
wire [31:0]	int_desc_10_axuser_2_axuser;
wire [31:0]	int_desc_10_axuser_3_axuser;
wire [31:0]	int_desc_10_axuser_4_axuser;
wire [31:0]	int_desc_10_axuser_5_axuser;
wire [31:0]	int_desc_10_axuser_6_axuser;
wire [31:0]	int_desc_10_axuser_7_axuser;
wire [31:0]	int_desc_10_axuser_8_axuser;
wire [31:0]	int_desc_10_axuser_9_axuser;
wire [31:0]	int_desc_10_axuser_10_axuser;
wire [31:0]	int_desc_10_axuser_11_axuser;
wire [31:0]	int_desc_10_axuser_12_axuser;
wire [31:0]	int_desc_10_axuser_13_axuser;
wire [31:0]	int_desc_10_axuser_14_axuser;
wire [31:0]	int_desc_10_axuser_15_axuser;
wire [15:0]	int_desc_10_size_txn_size;
wire [2:0]	int_desc_10_axsize_axsize;
wire [31:0]	int_desc_10_axaddr_0_addr;
wire [31:0]	int_desc_10_axaddr_1_addr;
wire [31:0]	int_desc_10_axaddr_2_addr;
wire [31:0]	int_desc_10_axaddr_3_addr;
wire [31:0]	int_desc_10_data_offset_addr;
wire [31:0]	int_desc_10_wuser_0_wuser;
wire [31:0]	int_desc_10_wuser_1_wuser;
wire [31:0]	int_desc_10_wuser_2_wuser;
wire [31:0]	int_desc_10_wuser_3_wuser;
wire [31:0]	int_desc_10_wuser_4_wuser;
wire [31:0]	int_desc_10_wuser_5_wuser;
wire [31:0]	int_desc_10_wuser_6_wuser;
wire [31:0]	int_desc_10_wuser_7_wuser;
wire [31:0]	int_desc_10_wuser_8_wuser;
wire [31:0]	int_desc_10_wuser_9_wuser;
wire [31:0]	int_desc_10_wuser_10_wuser;
wire [31:0]	int_desc_10_wuser_11_wuser;
wire [31:0]	int_desc_10_wuser_12_wuser;
wire [31:0]	int_desc_10_wuser_13_wuser;
wire [31:0]	int_desc_10_wuser_14_wuser;
wire [31:0]	int_desc_10_wuser_15_wuser;
wire [31:0]	int_desc_10_data_host_addr_0_addr;
wire [31:0]	int_desc_10_data_host_addr_1_addr;
wire [31:0]	int_desc_10_data_host_addr_2_addr;
wire [31:0]	int_desc_10_data_host_addr_3_addr;
wire [31:0]	int_desc_10_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_10_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_10_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_10_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_10_xuser_0_xuser;
wire [31:0]	int_desc_10_xuser_1_xuser;
wire [31:0]	int_desc_10_xuser_2_xuser;
wire [31:0]	int_desc_10_xuser_3_xuser;
wire [31:0]	int_desc_10_xuser_4_xuser;
wire [31:0]	int_desc_10_xuser_5_xuser;
wire [31:0]	int_desc_10_xuser_6_xuser;
wire [31:0]	int_desc_10_xuser_7_xuser;
wire [31:0]	int_desc_10_xuser_8_xuser;
wire [31:0]	int_desc_10_xuser_9_xuser;
wire [31:0]	int_desc_10_xuser_10_xuser;
wire [31:0]	int_desc_10_xuser_11_xuser;
wire [31:0]	int_desc_10_xuser_12_xuser;
wire [31:0]	int_desc_10_xuser_13_xuser;
wire [31:0]	int_desc_10_xuser_14_xuser;
wire [31:0]	int_desc_10_xuser_15_xuser;
wire [0:0]	int_desc_11_txn_type_wr_strb;
wire [0:0]	int_desc_11_txn_type_wr_rd;
wire [3:0]	int_desc_11_attr_axregion;
wire [3:0]	int_desc_11_attr_axqos;
wire [2:0]	int_desc_11_attr_axprot;
wire [3:0]	int_desc_11_attr_axcache;
wire [1:0]	int_desc_11_attr_axlock;
wire [1:0]	int_desc_11_attr_axburst;
wire [31:0]	int_desc_11_axid_0_axid;
wire [31:0]	int_desc_11_axid_1_axid;
wire [31:0]	int_desc_11_axid_2_axid;
wire [31:0]	int_desc_11_axid_3_axid;
wire [31:0]	int_desc_11_axuser_0_axuser;
wire [31:0]	int_desc_11_axuser_1_axuser;
wire [31:0]	int_desc_11_axuser_2_axuser;
wire [31:0]	int_desc_11_axuser_3_axuser;
wire [31:0]	int_desc_11_axuser_4_axuser;
wire [31:0]	int_desc_11_axuser_5_axuser;
wire [31:0]	int_desc_11_axuser_6_axuser;
wire [31:0]	int_desc_11_axuser_7_axuser;
wire [31:0]	int_desc_11_axuser_8_axuser;
wire [31:0]	int_desc_11_axuser_9_axuser;
wire [31:0]	int_desc_11_axuser_10_axuser;
wire [31:0]	int_desc_11_axuser_11_axuser;
wire [31:0]	int_desc_11_axuser_12_axuser;
wire [31:0]	int_desc_11_axuser_13_axuser;
wire [31:0]	int_desc_11_axuser_14_axuser;
wire [31:0]	int_desc_11_axuser_15_axuser;
wire [15:0]	int_desc_11_size_txn_size;
wire [2:0]	int_desc_11_axsize_axsize;
wire [31:0]	int_desc_11_axaddr_0_addr;
wire [31:0]	int_desc_11_axaddr_1_addr;
wire [31:0]	int_desc_11_axaddr_2_addr;
wire [31:0]	int_desc_11_axaddr_3_addr;
wire [31:0]	int_desc_11_data_offset_addr;
wire [31:0]	int_desc_11_wuser_0_wuser;
wire [31:0]	int_desc_11_wuser_1_wuser;
wire [31:0]	int_desc_11_wuser_2_wuser;
wire [31:0]	int_desc_11_wuser_3_wuser;
wire [31:0]	int_desc_11_wuser_4_wuser;
wire [31:0]	int_desc_11_wuser_5_wuser;
wire [31:0]	int_desc_11_wuser_6_wuser;
wire [31:0]	int_desc_11_wuser_7_wuser;
wire [31:0]	int_desc_11_wuser_8_wuser;
wire [31:0]	int_desc_11_wuser_9_wuser;
wire [31:0]	int_desc_11_wuser_10_wuser;
wire [31:0]	int_desc_11_wuser_11_wuser;
wire [31:0]	int_desc_11_wuser_12_wuser;
wire [31:0]	int_desc_11_wuser_13_wuser;
wire [31:0]	int_desc_11_wuser_14_wuser;
wire [31:0]	int_desc_11_wuser_15_wuser;
wire [31:0]	int_desc_11_data_host_addr_0_addr;
wire [31:0]	int_desc_11_data_host_addr_1_addr;
wire [31:0]	int_desc_11_data_host_addr_2_addr;
wire [31:0]	int_desc_11_data_host_addr_3_addr;
wire [31:0]	int_desc_11_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_11_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_11_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_11_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_11_xuser_0_xuser;
wire [31:0]	int_desc_11_xuser_1_xuser;
wire [31:0]	int_desc_11_xuser_2_xuser;
wire [31:0]	int_desc_11_xuser_3_xuser;
wire [31:0]	int_desc_11_xuser_4_xuser;
wire [31:0]	int_desc_11_xuser_5_xuser;
wire [31:0]	int_desc_11_xuser_6_xuser;
wire [31:0]	int_desc_11_xuser_7_xuser;
wire [31:0]	int_desc_11_xuser_8_xuser;
wire [31:0]	int_desc_11_xuser_9_xuser;
wire [31:0]	int_desc_11_xuser_10_xuser;
wire [31:0]	int_desc_11_xuser_11_xuser;
wire [31:0]	int_desc_11_xuser_12_xuser;
wire [31:0]	int_desc_11_xuser_13_xuser;
wire [31:0]	int_desc_11_xuser_14_xuser;
wire [31:0]	int_desc_11_xuser_15_xuser;
wire [0:0]	int_desc_12_txn_type_wr_strb;
wire [0:0]	int_desc_12_txn_type_wr_rd;
wire [3:0]	int_desc_12_attr_axregion;
wire [3:0]	int_desc_12_attr_axqos;
wire [2:0]	int_desc_12_attr_axprot;
wire [3:0]	int_desc_12_attr_axcache;
wire [1:0]	int_desc_12_attr_axlock;
wire [1:0]	int_desc_12_attr_axburst;
wire [31:0]	int_desc_12_axid_0_axid;
wire [31:0]	int_desc_12_axid_1_axid;
wire [31:0]	int_desc_12_axid_2_axid;
wire [31:0]	int_desc_12_axid_3_axid;
wire [31:0]	int_desc_12_axuser_0_axuser;
wire [31:0]	int_desc_12_axuser_1_axuser;
wire [31:0]	int_desc_12_axuser_2_axuser;
wire [31:0]	int_desc_12_axuser_3_axuser;
wire [31:0]	int_desc_12_axuser_4_axuser;
wire [31:0]	int_desc_12_axuser_5_axuser;
wire [31:0]	int_desc_12_axuser_6_axuser;
wire [31:0]	int_desc_12_axuser_7_axuser;
wire [31:0]	int_desc_12_axuser_8_axuser;
wire [31:0]	int_desc_12_axuser_9_axuser;
wire [31:0]	int_desc_12_axuser_10_axuser;
wire [31:0]	int_desc_12_axuser_11_axuser;
wire [31:0]	int_desc_12_axuser_12_axuser;
wire [31:0]	int_desc_12_axuser_13_axuser;
wire [31:0]	int_desc_12_axuser_14_axuser;
wire [31:0]	int_desc_12_axuser_15_axuser;
wire [15:0]	int_desc_12_size_txn_size;
wire [2:0]	int_desc_12_axsize_axsize;
wire [31:0]	int_desc_12_axaddr_0_addr;
wire [31:0]	int_desc_12_axaddr_1_addr;
wire [31:0]	int_desc_12_axaddr_2_addr;
wire [31:0]	int_desc_12_axaddr_3_addr;
wire [31:0]	int_desc_12_data_offset_addr;
wire [31:0]	int_desc_12_wuser_0_wuser;
wire [31:0]	int_desc_12_wuser_1_wuser;
wire [31:0]	int_desc_12_wuser_2_wuser;
wire [31:0]	int_desc_12_wuser_3_wuser;
wire [31:0]	int_desc_12_wuser_4_wuser;
wire [31:0]	int_desc_12_wuser_5_wuser;
wire [31:0]	int_desc_12_wuser_6_wuser;
wire [31:0]	int_desc_12_wuser_7_wuser;
wire [31:0]	int_desc_12_wuser_8_wuser;
wire [31:0]	int_desc_12_wuser_9_wuser;
wire [31:0]	int_desc_12_wuser_10_wuser;
wire [31:0]	int_desc_12_wuser_11_wuser;
wire [31:0]	int_desc_12_wuser_12_wuser;
wire [31:0]	int_desc_12_wuser_13_wuser;
wire [31:0]	int_desc_12_wuser_14_wuser;
wire [31:0]	int_desc_12_wuser_15_wuser;
wire [31:0]	int_desc_12_data_host_addr_0_addr;
wire [31:0]	int_desc_12_data_host_addr_1_addr;
wire [31:0]	int_desc_12_data_host_addr_2_addr;
wire [31:0]	int_desc_12_data_host_addr_3_addr;
wire [31:0]	int_desc_12_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_12_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_12_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_12_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_12_xuser_0_xuser;
wire [31:0]	int_desc_12_xuser_1_xuser;
wire [31:0]	int_desc_12_xuser_2_xuser;
wire [31:0]	int_desc_12_xuser_3_xuser;
wire [31:0]	int_desc_12_xuser_4_xuser;
wire [31:0]	int_desc_12_xuser_5_xuser;
wire [31:0]	int_desc_12_xuser_6_xuser;
wire [31:0]	int_desc_12_xuser_7_xuser;
wire [31:0]	int_desc_12_xuser_8_xuser;
wire [31:0]	int_desc_12_xuser_9_xuser;
wire [31:0]	int_desc_12_xuser_10_xuser;
wire [31:0]	int_desc_12_xuser_11_xuser;
wire [31:0]	int_desc_12_xuser_12_xuser;
wire [31:0]	int_desc_12_xuser_13_xuser;
wire [31:0]	int_desc_12_xuser_14_xuser;
wire [31:0]	int_desc_12_xuser_15_xuser;
wire [0:0]	int_desc_13_txn_type_wr_strb;
wire [0:0]	int_desc_13_txn_type_wr_rd;
wire [3:0]	int_desc_13_attr_axregion;
wire [3:0]	int_desc_13_attr_axqos;
wire [2:0]	int_desc_13_attr_axprot;
wire [3:0]	int_desc_13_attr_axcache;
wire [1:0]	int_desc_13_attr_axlock;
wire [1:0]	int_desc_13_attr_axburst;
wire [31:0]	int_desc_13_axid_0_axid;
wire [31:0]	int_desc_13_axid_1_axid;
wire [31:0]	int_desc_13_axid_2_axid;
wire [31:0]	int_desc_13_axid_3_axid;
wire [31:0]	int_desc_13_axuser_0_axuser;
wire [31:0]	int_desc_13_axuser_1_axuser;
wire [31:0]	int_desc_13_axuser_2_axuser;
wire [31:0]	int_desc_13_axuser_3_axuser;
wire [31:0]	int_desc_13_axuser_4_axuser;
wire [31:0]	int_desc_13_axuser_5_axuser;
wire [31:0]	int_desc_13_axuser_6_axuser;
wire [31:0]	int_desc_13_axuser_7_axuser;
wire [31:0]	int_desc_13_axuser_8_axuser;
wire [31:0]	int_desc_13_axuser_9_axuser;
wire [31:0]	int_desc_13_axuser_10_axuser;
wire [31:0]	int_desc_13_axuser_11_axuser;
wire [31:0]	int_desc_13_axuser_12_axuser;
wire [31:0]	int_desc_13_axuser_13_axuser;
wire [31:0]	int_desc_13_axuser_14_axuser;
wire [31:0]	int_desc_13_axuser_15_axuser;
wire [15:0]	int_desc_13_size_txn_size;
wire [2:0]	int_desc_13_axsize_axsize;
wire [31:0]	int_desc_13_axaddr_0_addr;
wire [31:0]	int_desc_13_axaddr_1_addr;
wire [31:0]	int_desc_13_axaddr_2_addr;
wire [31:0]	int_desc_13_axaddr_3_addr;
wire [31:0]	int_desc_13_data_offset_addr;
wire [31:0]	int_desc_13_wuser_0_wuser;
wire [31:0]	int_desc_13_wuser_1_wuser;
wire [31:0]	int_desc_13_wuser_2_wuser;
wire [31:0]	int_desc_13_wuser_3_wuser;
wire [31:0]	int_desc_13_wuser_4_wuser;
wire [31:0]	int_desc_13_wuser_5_wuser;
wire [31:0]	int_desc_13_wuser_6_wuser;
wire [31:0]	int_desc_13_wuser_7_wuser;
wire [31:0]	int_desc_13_wuser_8_wuser;
wire [31:0]	int_desc_13_wuser_9_wuser;
wire [31:0]	int_desc_13_wuser_10_wuser;
wire [31:0]	int_desc_13_wuser_11_wuser;
wire [31:0]	int_desc_13_wuser_12_wuser;
wire [31:0]	int_desc_13_wuser_13_wuser;
wire [31:0]	int_desc_13_wuser_14_wuser;
wire [31:0]	int_desc_13_wuser_15_wuser;
wire [31:0]	int_desc_13_data_host_addr_0_addr;
wire [31:0]	int_desc_13_data_host_addr_1_addr;
wire [31:0]	int_desc_13_data_host_addr_2_addr;
wire [31:0]	int_desc_13_data_host_addr_3_addr;
wire [31:0]	int_desc_13_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_13_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_13_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_13_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_13_xuser_0_xuser;
wire [31:0]	int_desc_13_xuser_1_xuser;
wire [31:0]	int_desc_13_xuser_2_xuser;
wire [31:0]	int_desc_13_xuser_3_xuser;
wire [31:0]	int_desc_13_xuser_4_xuser;
wire [31:0]	int_desc_13_xuser_5_xuser;
wire [31:0]	int_desc_13_xuser_6_xuser;
wire [31:0]	int_desc_13_xuser_7_xuser;
wire [31:0]	int_desc_13_xuser_8_xuser;
wire [31:0]	int_desc_13_xuser_9_xuser;
wire [31:0]	int_desc_13_xuser_10_xuser;
wire [31:0]	int_desc_13_xuser_11_xuser;
wire [31:0]	int_desc_13_xuser_12_xuser;
wire [31:0]	int_desc_13_xuser_13_xuser;
wire [31:0]	int_desc_13_xuser_14_xuser;
wire [31:0]	int_desc_13_xuser_15_xuser;
wire [0:0]	int_desc_14_txn_type_wr_strb;
wire [0:0]	int_desc_14_txn_type_wr_rd;
wire [3:0]	int_desc_14_attr_axregion;
wire [3:0]	int_desc_14_attr_axqos;
wire [2:0]	int_desc_14_attr_axprot;
wire [3:0]	int_desc_14_attr_axcache;
wire [1:0]	int_desc_14_attr_axlock;
wire [1:0]	int_desc_14_attr_axburst;
wire [31:0]	int_desc_14_axid_0_axid;
wire [31:0]	int_desc_14_axid_1_axid;
wire [31:0]	int_desc_14_axid_2_axid;
wire [31:0]	int_desc_14_axid_3_axid;
wire [31:0]	int_desc_14_axuser_0_axuser;
wire [31:0]	int_desc_14_axuser_1_axuser;
wire [31:0]	int_desc_14_axuser_2_axuser;
wire [31:0]	int_desc_14_axuser_3_axuser;
wire [31:0]	int_desc_14_axuser_4_axuser;
wire [31:0]	int_desc_14_axuser_5_axuser;
wire [31:0]	int_desc_14_axuser_6_axuser;
wire [31:0]	int_desc_14_axuser_7_axuser;
wire [31:0]	int_desc_14_axuser_8_axuser;
wire [31:0]	int_desc_14_axuser_9_axuser;
wire [31:0]	int_desc_14_axuser_10_axuser;
wire [31:0]	int_desc_14_axuser_11_axuser;
wire [31:0]	int_desc_14_axuser_12_axuser;
wire [31:0]	int_desc_14_axuser_13_axuser;
wire [31:0]	int_desc_14_axuser_14_axuser;
wire [31:0]	int_desc_14_axuser_15_axuser;
wire [15:0]	int_desc_14_size_txn_size;
wire [2:0]	int_desc_14_axsize_axsize;
wire [31:0]	int_desc_14_axaddr_0_addr;
wire [31:0]	int_desc_14_axaddr_1_addr;
wire [31:0]	int_desc_14_axaddr_2_addr;
wire [31:0]	int_desc_14_axaddr_3_addr;
wire [31:0]	int_desc_14_data_offset_addr;
wire [31:0]	int_desc_14_wuser_0_wuser;
wire [31:0]	int_desc_14_wuser_1_wuser;
wire [31:0]	int_desc_14_wuser_2_wuser;
wire [31:0]	int_desc_14_wuser_3_wuser;
wire [31:0]	int_desc_14_wuser_4_wuser;
wire [31:0]	int_desc_14_wuser_5_wuser;
wire [31:0]	int_desc_14_wuser_6_wuser;
wire [31:0]	int_desc_14_wuser_7_wuser;
wire [31:0]	int_desc_14_wuser_8_wuser;
wire [31:0]	int_desc_14_wuser_9_wuser;
wire [31:0]	int_desc_14_wuser_10_wuser;
wire [31:0]	int_desc_14_wuser_11_wuser;
wire [31:0]	int_desc_14_wuser_12_wuser;
wire [31:0]	int_desc_14_wuser_13_wuser;
wire [31:0]	int_desc_14_wuser_14_wuser;
wire [31:0]	int_desc_14_wuser_15_wuser;
wire [31:0]	int_desc_14_data_host_addr_0_addr;
wire [31:0]	int_desc_14_data_host_addr_1_addr;
wire [31:0]	int_desc_14_data_host_addr_2_addr;
wire [31:0]	int_desc_14_data_host_addr_3_addr;
wire [31:0]	int_desc_14_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_14_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_14_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_14_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_14_xuser_0_xuser;
wire [31:0]	int_desc_14_xuser_1_xuser;
wire [31:0]	int_desc_14_xuser_2_xuser;
wire [31:0]	int_desc_14_xuser_3_xuser;
wire [31:0]	int_desc_14_xuser_4_xuser;
wire [31:0]	int_desc_14_xuser_5_xuser;
wire [31:0]	int_desc_14_xuser_6_xuser;
wire [31:0]	int_desc_14_xuser_7_xuser;
wire [31:0]	int_desc_14_xuser_8_xuser;
wire [31:0]	int_desc_14_xuser_9_xuser;
wire [31:0]	int_desc_14_xuser_10_xuser;
wire [31:0]	int_desc_14_xuser_11_xuser;
wire [31:0]	int_desc_14_xuser_12_xuser;
wire [31:0]	int_desc_14_xuser_13_xuser;
wire [31:0]	int_desc_14_xuser_14_xuser;
wire [31:0]	int_desc_14_xuser_15_xuser;
wire [0:0]	int_desc_15_txn_type_wr_strb;
wire [0:0]	int_desc_15_txn_type_wr_rd;
wire [3:0]	int_desc_15_attr_axregion;
wire [3:0]	int_desc_15_attr_axqos;
wire [2:0]	int_desc_15_attr_axprot;
wire [3:0]	int_desc_15_attr_axcache;
wire [1:0]	int_desc_15_attr_axlock;
wire [1:0]	int_desc_15_attr_axburst;
wire [31:0]	int_desc_15_axid_0_axid;
wire [31:0]	int_desc_15_axid_1_axid;
wire [31:0]	int_desc_15_axid_2_axid;
wire [31:0]	int_desc_15_axid_3_axid;
wire [31:0]	int_desc_15_axuser_0_axuser;
wire [31:0]	int_desc_15_axuser_1_axuser;
wire [31:0]	int_desc_15_axuser_2_axuser;
wire [31:0]	int_desc_15_axuser_3_axuser;
wire [31:0]	int_desc_15_axuser_4_axuser;
wire [31:0]	int_desc_15_axuser_5_axuser;
wire [31:0]	int_desc_15_axuser_6_axuser;
wire [31:0]	int_desc_15_axuser_7_axuser;
wire [31:0]	int_desc_15_axuser_8_axuser;
wire [31:0]	int_desc_15_axuser_9_axuser;
wire [31:0]	int_desc_15_axuser_10_axuser;
wire [31:0]	int_desc_15_axuser_11_axuser;
wire [31:0]	int_desc_15_axuser_12_axuser;
wire [31:0]	int_desc_15_axuser_13_axuser;
wire [31:0]	int_desc_15_axuser_14_axuser;
wire [31:0]	int_desc_15_axuser_15_axuser;
wire [15:0]	int_desc_15_size_txn_size;
wire [2:0]	int_desc_15_axsize_axsize;
wire [31:0]	int_desc_15_axaddr_0_addr;
wire [31:0]	int_desc_15_axaddr_1_addr;
wire [31:0]	int_desc_15_axaddr_2_addr;
wire [31:0]	int_desc_15_axaddr_3_addr;
wire [31:0]	int_desc_15_data_offset_addr;
wire [31:0]	int_desc_15_wuser_0_wuser;
wire [31:0]	int_desc_15_wuser_1_wuser;
wire [31:0]	int_desc_15_wuser_2_wuser;
wire [31:0]	int_desc_15_wuser_3_wuser;
wire [31:0]	int_desc_15_wuser_4_wuser;
wire [31:0]	int_desc_15_wuser_5_wuser;
wire [31:0]	int_desc_15_wuser_6_wuser;
wire [31:0]	int_desc_15_wuser_7_wuser;
wire [31:0]	int_desc_15_wuser_8_wuser;
wire [31:0]	int_desc_15_wuser_9_wuser;
wire [31:0]	int_desc_15_wuser_10_wuser;
wire [31:0]	int_desc_15_wuser_11_wuser;
wire [31:0]	int_desc_15_wuser_12_wuser;
wire [31:0]	int_desc_15_wuser_13_wuser;
wire [31:0]	int_desc_15_wuser_14_wuser;
wire [31:0]	int_desc_15_wuser_15_wuser;
wire [31:0]	int_desc_15_data_host_addr_0_addr;
wire [31:0]	int_desc_15_data_host_addr_1_addr;
wire [31:0]	int_desc_15_data_host_addr_2_addr;
wire [31:0]	int_desc_15_data_host_addr_3_addr;
wire [31:0]	int_desc_15_wstrb_host_addr_0_addr;
wire [31:0]	int_desc_15_wstrb_host_addr_1_addr;
wire [31:0]	int_desc_15_wstrb_host_addr_2_addr;
wire [31:0]	int_desc_15_wstrb_host_addr_3_addr;
wire [31:0]	int_desc_15_xuser_0_xuser;
wire [31:0]	int_desc_15_xuser_1_xuser;
wire [31:0]	int_desc_15_xuser_2_xuser;
wire [31:0]	int_desc_15_xuser_3_xuser;
wire [31:0]	int_desc_15_xuser_4_xuser;
wire [31:0]	int_desc_15_xuser_5_xuser;
wire [31:0]	int_desc_15_xuser_6_xuser;
wire [31:0]	int_desc_15_xuser_7_xuser;
wire [31:0]	int_desc_15_xuser_8_xuser;
wire [31:0]	int_desc_15_xuser_9_xuser;
wire [31:0]	int_desc_15_xuser_10_xuser;
wire [31:0]	int_desc_15_xuser_11_xuser;
wire [31:0]	int_desc_15_xuser_12_xuser;
wire [31:0]	int_desc_15_xuser_13_xuser;
wire [31:0]	int_desc_15_xuser_14_xuser;
wire [31:0]	int_desc_15_xuser_15_xuser;

//////////////////////
//Derive fields from registers of RB
//////////////////////

assign version_major_ver_f = version_reg[15:8];
assign version_minor_ver_f = version_reg[7:0];
assign bridge_type_type_f = bridge_type_reg[7:0];
assign axi_bridge_config_user_width_f = axi_bridge_config_reg[23:16];
assign axi_bridge_config_id_width_f = axi_bridge_config_reg[11:4];
assign axi_bridge_config_data_width_f = axi_bridge_config_reg[2:0];
assign reset_dut_srst_3_f = reset_reg[4];
assign reset_dut_srst_2_f = reset_reg[3];
assign reset_dut_srst_1_f = reset_reg[2];
assign reset_dut_srst_0_f = reset_reg[1];
assign reset_srst_f = reset_reg[0];
assign mode_select_imm_bresp_f = mode_select_reg[2];
assign mode_select_mode_2_f = mode_select_reg[1];
assign mode_select_mode_0_1_f = mode_select_reg[0];
assign ownership_own_f = ownership_reg[MAX_DESC-1:0];
assign ownership_flip_flip_f = ownership_flip_reg[MAX_DESC-1:0];
assign status_resp_comp_resp_comp_f = status_resp_comp_reg[MAX_DESC-1:0];
assign status_resp_resp_f = status_resp_reg[31:0];
assign status_busy_busy_f = status_busy_reg[MAX_DESC-1:0];
assign resp_fifo_free_level_level_f = resp_fifo_free_level_reg[DESC_IDX_WIDTH:0];
assign intr_status_comp_f = intr_status_reg[3];
assign intr_status_c2h_f = intr_status_reg[2];
assign intr_status_error_f = intr_status_reg[1];
assign intr_status_txn_avail_f = intr_status_reg[0];
assign intr_txn_avail_status_avail_f = intr_txn_avail_status_reg[MAX_DESC-1:0];
assign intr_txn_avail_clear_clr_avail_f = intr_txn_avail_clear_reg[MAX_DESC-1:0];
assign intr_txn_avail_enable_en_avail_f = intr_txn_avail_enable_reg[MAX_DESC-1:0];
assign intr_comp_status_comp_f = intr_comp_status_reg[MAX_DESC-1:0];
assign intr_comp_clear_clr_comp_f = intr_comp_clear_reg[MAX_DESC-1:0];
assign intr_comp_enable_en_comp_f = intr_comp_enable_reg[MAX_DESC-1:0];
assign intr_error_status_err_2_f = intr_error_status_reg[2];
assign intr_error_status_err_1_f = intr_error_status_reg[1];
assign intr_error_status_err_0_f = intr_error_status_reg[0];
assign intr_error_clear_clr_err_2_f = intr_error_clear_reg[2];
assign intr_error_clear_clr_err_1_f = intr_error_clear_reg[1];
assign intr_error_clear_clr_err_0_f = intr_error_clear_reg[0];
assign intr_error_enable_en_err_2_f = intr_error_enable_reg[2];
assign intr_error_enable_en_err_1_f = intr_error_enable_reg[1];
assign intr_error_enable_en_err_0_f = intr_error_enable_reg[0];
assign intr_h2c_0_h2c_f = intr_h2c_0_reg[31:0];
assign intr_h2c_1_h2c_f = intr_h2c_1_reg[31:0];
assign intr_c2h_0_status_c2h_f = intr_c2h_0_status_reg[31:0];
assign intr_c2h_1_status_c2h_f = intr_c2h_1_status_reg[31:0];
assign c2h_gpio_0_status_gpio_f = c2h_gpio_0_status_reg[31:0];
assign c2h_gpio_1_status_gpio_f = c2h_gpio_1_status_reg[31:0];
assign c2h_gpio_2_status_gpio_f = c2h_gpio_2_status_reg[31:0];
assign c2h_gpio_3_status_gpio_f = c2h_gpio_3_status_reg[31:0];
assign c2h_gpio_4_status_gpio_f = c2h_gpio_4_status_reg[31:0];
assign c2h_gpio_5_status_gpio_f = c2h_gpio_5_status_reg[31:0];
assign c2h_gpio_6_status_gpio_f = c2h_gpio_6_status_reg[31:0];
assign c2h_gpio_7_status_gpio_f = c2h_gpio_7_status_reg[31:0];
assign c2h_gpio_8_status_gpio_f = c2h_gpio_8_status_reg[31:0];
assign c2h_gpio_9_status_gpio_f = c2h_gpio_9_status_reg[31:0];
assign c2h_gpio_10_status_gpio_f = c2h_gpio_10_status_reg[31:0];
assign c2h_gpio_11_status_gpio_f = c2h_gpio_11_status_reg[31:0];
assign c2h_gpio_12_status_gpio_f = c2h_gpio_12_status_reg[31:0];
assign c2h_gpio_13_status_gpio_f = c2h_gpio_13_status_reg[31:0];
assign c2h_gpio_14_status_gpio_f = c2h_gpio_14_status_reg[31:0];
assign c2h_gpio_15_status_gpio_f = c2h_gpio_15_status_reg[31:0];
assign addr_in_0_addr_f = addr_in_0_reg[31:0];
assign addr_in_1_addr_f = addr_in_1_reg[31:0];
assign addr_in_2_addr_f = addr_in_2_reg[31:0];
assign addr_in_3_addr_f = addr_in_3_reg[31:0];
assign trans_mask_0_addr_f = trans_mask_0_reg[31:0];
assign trans_mask_1_addr_f = trans_mask_1_reg[31:0];
assign trans_mask_2_addr_f = trans_mask_2_reg[31:0];
assign trans_mask_3_addr_f = trans_mask_3_reg[31:0];
assign trans_addr_0_addr_f = trans_addr_0_reg[31:0];
assign trans_addr_1_addr_f = trans_addr_1_reg[31:0];
assign trans_addr_2_addr_f = trans_addr_2_reg[31:0];
assign trans_addr_3_addr_f = trans_addr_3_reg[31:0];
assign resp_order_field_f = resp_order_reg[31:0];

assign desc_0_txn_type_wr_strb_f = desc_0_txn_type_reg[1];
assign desc_0_txn_type_wr_rd_f = desc_0_txn_type_reg[0];
assign desc_0_attr_axregion_f = desc_0_attr_reg[18:15];
assign desc_0_attr_axqos_f = desc_0_attr_reg[14:11];
assign desc_0_attr_axprot_f = desc_0_attr_reg[10:8];
assign desc_0_attr_axcache_f = desc_0_attr_reg[7:4];
assign desc_0_attr_axlock_f = desc_0_attr_reg[3:2];
assign desc_0_attr_axburst_f = desc_0_attr_reg[1:0];
assign desc_0_axid_0_axid_f = desc_0_axid_0_reg[31:0];
assign desc_0_axid_1_axid_f = desc_0_axid_1_reg[31:0];
assign desc_0_axid_2_axid_f = desc_0_axid_2_reg[31:0];
assign desc_0_axid_3_axid_f = desc_0_axid_3_reg[31:0];
assign desc_0_axuser_0_axuser_f = desc_0_axuser_0_reg[31:0];
assign desc_0_axuser_1_axuser_f = desc_0_axuser_1_reg[31:0];
assign desc_0_axuser_2_axuser_f = desc_0_axuser_2_reg[31:0];
assign desc_0_axuser_3_axuser_f = desc_0_axuser_3_reg[31:0];
assign desc_0_axuser_4_axuser_f = desc_0_axuser_4_reg[31:0];
assign desc_0_axuser_5_axuser_f = desc_0_axuser_5_reg[31:0];
assign desc_0_axuser_6_axuser_f = desc_0_axuser_6_reg[31:0];
assign desc_0_axuser_7_axuser_f = desc_0_axuser_7_reg[31:0];
assign desc_0_axuser_8_axuser_f = desc_0_axuser_8_reg[31:0];
assign desc_0_axuser_9_axuser_f = desc_0_axuser_9_reg[31:0];
assign desc_0_axuser_10_axuser_f = desc_0_axuser_10_reg[31:0];
assign desc_0_axuser_11_axuser_f = desc_0_axuser_11_reg[31:0];
assign desc_0_axuser_12_axuser_f = desc_0_axuser_12_reg[31:0];
assign desc_0_axuser_13_axuser_f = desc_0_axuser_13_reg[31:0];
assign desc_0_axuser_14_axuser_f = desc_0_axuser_14_reg[31:0];
assign desc_0_axuser_15_axuser_f = desc_0_axuser_15_reg[31:0];
assign desc_0_size_txn_size_f = desc_0_size_reg[15:0];
assign desc_0_axsize_axsize_f = desc_0_axsize_reg[2:0];
assign desc_0_axaddr_0_addr_f = desc_0_axaddr_0_reg[31:0];
assign desc_0_axaddr_1_addr_f = desc_0_axaddr_1_reg[31:0];
assign desc_0_axaddr_2_addr_f = desc_0_axaddr_2_reg[31:0];
assign desc_0_axaddr_3_addr_f = desc_0_axaddr_3_reg[31:0];
assign desc_0_data_offset_addr_f = desc_0_data_offset_reg[31:0];
assign desc_0_wuser_0_wuser_f = desc_0_wuser_0_reg[31:0];
assign desc_0_wuser_1_wuser_f = desc_0_wuser_1_reg[31:0];
assign desc_0_wuser_2_wuser_f = desc_0_wuser_2_reg[31:0];
assign desc_0_wuser_3_wuser_f = desc_0_wuser_3_reg[31:0];
assign desc_0_wuser_4_wuser_f = desc_0_wuser_4_reg[31:0];
assign desc_0_wuser_5_wuser_f = desc_0_wuser_5_reg[31:0];
assign desc_0_wuser_6_wuser_f = desc_0_wuser_6_reg[31:0];
assign desc_0_wuser_7_wuser_f = desc_0_wuser_7_reg[31:0];
assign desc_0_wuser_8_wuser_f = desc_0_wuser_8_reg[31:0];
assign desc_0_wuser_9_wuser_f = desc_0_wuser_9_reg[31:0];
assign desc_0_wuser_10_wuser_f = desc_0_wuser_10_reg[31:0];
assign desc_0_wuser_11_wuser_f = desc_0_wuser_11_reg[31:0];
assign desc_0_wuser_12_wuser_f = desc_0_wuser_12_reg[31:0];
assign desc_0_wuser_13_wuser_f = desc_0_wuser_13_reg[31:0];
assign desc_0_wuser_14_wuser_f = desc_0_wuser_14_reg[31:0];
assign desc_0_wuser_15_wuser_f = desc_0_wuser_15_reg[31:0];
assign desc_0_data_host_addr_0_addr_f = desc_0_data_host_addr_0_reg[31:0];
assign desc_0_data_host_addr_1_addr_f = desc_0_data_host_addr_1_reg[31:0];
assign desc_0_data_host_addr_2_addr_f = desc_0_data_host_addr_2_reg[31:0];
assign desc_0_data_host_addr_3_addr_f = desc_0_data_host_addr_3_reg[31:0];
assign desc_0_wstrb_host_addr_0_addr_f = desc_0_wstrb_host_addr_0_reg[31:0];
assign desc_0_wstrb_host_addr_1_addr_f = desc_0_wstrb_host_addr_1_reg[31:0];
assign desc_0_wstrb_host_addr_2_addr_f = desc_0_wstrb_host_addr_2_reg[31:0];
assign desc_0_wstrb_host_addr_3_addr_f = desc_0_wstrb_host_addr_3_reg[31:0];
assign desc_0_xuser_0_xuser_f = desc_0_xuser_0_reg[31:0];
assign desc_0_xuser_1_xuser_f = desc_0_xuser_1_reg[31:0];
assign desc_0_xuser_2_xuser_f = desc_0_xuser_2_reg[31:0];
assign desc_0_xuser_3_xuser_f = desc_0_xuser_3_reg[31:0];
assign desc_0_xuser_4_xuser_f = desc_0_xuser_4_reg[31:0];
assign desc_0_xuser_5_xuser_f = desc_0_xuser_5_reg[31:0];
assign desc_0_xuser_6_xuser_f = desc_0_xuser_6_reg[31:0];
assign desc_0_xuser_7_xuser_f = desc_0_xuser_7_reg[31:0];
assign desc_0_xuser_8_xuser_f = desc_0_xuser_8_reg[31:0];
assign desc_0_xuser_9_xuser_f = desc_0_xuser_9_reg[31:0];
assign desc_0_xuser_10_xuser_f = desc_0_xuser_10_reg[31:0];
assign desc_0_xuser_11_xuser_f = desc_0_xuser_11_reg[31:0];
assign desc_0_xuser_12_xuser_f = desc_0_xuser_12_reg[31:0];
assign desc_0_xuser_13_xuser_f = desc_0_xuser_13_reg[31:0];
assign desc_0_xuser_14_xuser_f = desc_0_xuser_14_reg[31:0];
assign desc_0_xuser_15_xuser_f = desc_0_xuser_15_reg[31:0];
assign desc_1_txn_type_wr_strb_f = desc_1_txn_type_reg[1];
assign desc_1_txn_type_wr_rd_f = desc_1_txn_type_reg[0];
assign desc_1_attr_axregion_f = desc_1_attr_reg[18:15];
assign desc_1_attr_axqos_f = desc_1_attr_reg[14:11];
assign desc_1_attr_axprot_f = desc_1_attr_reg[10:8];
assign desc_1_attr_axcache_f = desc_1_attr_reg[7:4];
assign desc_1_attr_axlock_f = desc_1_attr_reg[3:2];
assign desc_1_attr_axburst_f = desc_1_attr_reg[1:0];
assign desc_1_axid_0_axid_f = desc_1_axid_0_reg[31:0];
assign desc_1_axid_1_axid_f = desc_1_axid_1_reg[31:0];
assign desc_1_axid_2_axid_f = desc_1_axid_2_reg[31:0];
assign desc_1_axid_3_axid_f = desc_1_axid_3_reg[31:0];
assign desc_1_axuser_0_axuser_f = desc_1_axuser_0_reg[31:0];
assign desc_1_axuser_1_axuser_f = desc_1_axuser_1_reg[31:0];
assign desc_1_axuser_2_axuser_f = desc_1_axuser_2_reg[31:0];
assign desc_1_axuser_3_axuser_f = desc_1_axuser_3_reg[31:0];
assign desc_1_axuser_4_axuser_f = desc_1_axuser_4_reg[31:0];
assign desc_1_axuser_5_axuser_f = desc_1_axuser_5_reg[31:0];
assign desc_1_axuser_6_axuser_f = desc_1_axuser_6_reg[31:0];
assign desc_1_axuser_7_axuser_f = desc_1_axuser_7_reg[31:0];
assign desc_1_axuser_8_axuser_f = desc_1_axuser_8_reg[31:0];
assign desc_1_axuser_9_axuser_f = desc_1_axuser_9_reg[31:0];
assign desc_1_axuser_10_axuser_f = desc_1_axuser_10_reg[31:0];
assign desc_1_axuser_11_axuser_f = desc_1_axuser_11_reg[31:0];
assign desc_1_axuser_12_axuser_f = desc_1_axuser_12_reg[31:0];
assign desc_1_axuser_13_axuser_f = desc_1_axuser_13_reg[31:0];
assign desc_1_axuser_14_axuser_f = desc_1_axuser_14_reg[31:0];
assign desc_1_axuser_15_axuser_f = desc_1_axuser_15_reg[31:0];
assign desc_1_size_txn_size_f = desc_1_size_reg[15:0];
assign desc_1_axsize_axsize_f = desc_1_axsize_reg[2:0];
assign desc_1_axaddr_0_addr_f = desc_1_axaddr_0_reg[31:0];
assign desc_1_axaddr_1_addr_f = desc_1_axaddr_1_reg[31:0];
assign desc_1_axaddr_2_addr_f = desc_1_axaddr_2_reg[31:0];
assign desc_1_axaddr_3_addr_f = desc_1_axaddr_3_reg[31:0];
assign desc_1_data_offset_addr_f = desc_1_data_offset_reg[31:0];
assign desc_1_wuser_0_wuser_f = desc_1_wuser_0_reg[31:0];
assign desc_1_wuser_1_wuser_f = desc_1_wuser_1_reg[31:0];
assign desc_1_wuser_2_wuser_f = desc_1_wuser_2_reg[31:0];
assign desc_1_wuser_3_wuser_f = desc_1_wuser_3_reg[31:0];
assign desc_1_wuser_4_wuser_f = desc_1_wuser_4_reg[31:0];
assign desc_1_wuser_5_wuser_f = desc_1_wuser_5_reg[31:0];
assign desc_1_wuser_6_wuser_f = desc_1_wuser_6_reg[31:0];
assign desc_1_wuser_7_wuser_f = desc_1_wuser_7_reg[31:0];
assign desc_1_wuser_8_wuser_f = desc_1_wuser_8_reg[31:0];
assign desc_1_wuser_9_wuser_f = desc_1_wuser_9_reg[31:0];
assign desc_1_wuser_10_wuser_f = desc_1_wuser_10_reg[31:0];
assign desc_1_wuser_11_wuser_f = desc_1_wuser_11_reg[31:0];
assign desc_1_wuser_12_wuser_f = desc_1_wuser_12_reg[31:0];
assign desc_1_wuser_13_wuser_f = desc_1_wuser_13_reg[31:0];
assign desc_1_wuser_14_wuser_f = desc_1_wuser_14_reg[31:0];
assign desc_1_wuser_15_wuser_f = desc_1_wuser_15_reg[31:0];
assign desc_1_data_host_addr_0_addr_f = desc_1_data_host_addr_0_reg[31:0];
assign desc_1_data_host_addr_1_addr_f = desc_1_data_host_addr_1_reg[31:0];
assign desc_1_data_host_addr_2_addr_f = desc_1_data_host_addr_2_reg[31:0];
assign desc_1_data_host_addr_3_addr_f = desc_1_data_host_addr_3_reg[31:0];
assign desc_1_wstrb_host_addr_0_addr_f = desc_1_wstrb_host_addr_0_reg[31:0];
assign desc_1_wstrb_host_addr_1_addr_f = desc_1_wstrb_host_addr_1_reg[31:0];
assign desc_1_wstrb_host_addr_2_addr_f = desc_1_wstrb_host_addr_2_reg[31:0];
assign desc_1_wstrb_host_addr_3_addr_f = desc_1_wstrb_host_addr_3_reg[31:0];
assign desc_1_xuser_0_xuser_f = desc_1_xuser_0_reg[31:0];
assign desc_1_xuser_1_xuser_f = desc_1_xuser_1_reg[31:0];
assign desc_1_xuser_2_xuser_f = desc_1_xuser_2_reg[31:0];
assign desc_1_xuser_3_xuser_f = desc_1_xuser_3_reg[31:0];
assign desc_1_xuser_4_xuser_f = desc_1_xuser_4_reg[31:0];
assign desc_1_xuser_5_xuser_f = desc_1_xuser_5_reg[31:0];
assign desc_1_xuser_6_xuser_f = desc_1_xuser_6_reg[31:0];
assign desc_1_xuser_7_xuser_f = desc_1_xuser_7_reg[31:0];
assign desc_1_xuser_8_xuser_f = desc_1_xuser_8_reg[31:0];
assign desc_1_xuser_9_xuser_f = desc_1_xuser_9_reg[31:0];
assign desc_1_xuser_10_xuser_f = desc_1_xuser_10_reg[31:0];
assign desc_1_xuser_11_xuser_f = desc_1_xuser_11_reg[31:0];
assign desc_1_xuser_12_xuser_f = desc_1_xuser_12_reg[31:0];
assign desc_1_xuser_13_xuser_f = desc_1_xuser_13_reg[31:0];
assign desc_1_xuser_14_xuser_f = desc_1_xuser_14_reg[31:0];
assign desc_1_xuser_15_xuser_f = desc_1_xuser_15_reg[31:0];
assign desc_2_txn_type_wr_strb_f = desc_2_txn_type_reg[1];
assign desc_2_txn_type_wr_rd_f = desc_2_txn_type_reg[0];
assign desc_2_attr_axregion_f = desc_2_attr_reg[18:15];
assign desc_2_attr_axqos_f = desc_2_attr_reg[14:11];
assign desc_2_attr_axprot_f = desc_2_attr_reg[10:8];
assign desc_2_attr_axcache_f = desc_2_attr_reg[7:4];
assign desc_2_attr_axlock_f = desc_2_attr_reg[3:2];
assign desc_2_attr_axburst_f = desc_2_attr_reg[1:0];
assign desc_2_axid_0_axid_f = desc_2_axid_0_reg[31:0];
assign desc_2_axid_1_axid_f = desc_2_axid_1_reg[31:0];
assign desc_2_axid_2_axid_f = desc_2_axid_2_reg[31:0];
assign desc_2_axid_3_axid_f = desc_2_axid_3_reg[31:0];
assign desc_2_axuser_0_axuser_f = desc_2_axuser_0_reg[31:0];
assign desc_2_axuser_1_axuser_f = desc_2_axuser_1_reg[31:0];
assign desc_2_axuser_2_axuser_f = desc_2_axuser_2_reg[31:0];
assign desc_2_axuser_3_axuser_f = desc_2_axuser_3_reg[31:0];
assign desc_2_axuser_4_axuser_f = desc_2_axuser_4_reg[31:0];
assign desc_2_axuser_5_axuser_f = desc_2_axuser_5_reg[31:0];
assign desc_2_axuser_6_axuser_f = desc_2_axuser_6_reg[31:0];
assign desc_2_axuser_7_axuser_f = desc_2_axuser_7_reg[31:0];
assign desc_2_axuser_8_axuser_f = desc_2_axuser_8_reg[31:0];
assign desc_2_axuser_9_axuser_f = desc_2_axuser_9_reg[31:0];
assign desc_2_axuser_10_axuser_f = desc_2_axuser_10_reg[31:0];
assign desc_2_axuser_11_axuser_f = desc_2_axuser_11_reg[31:0];
assign desc_2_axuser_12_axuser_f = desc_2_axuser_12_reg[31:0];
assign desc_2_axuser_13_axuser_f = desc_2_axuser_13_reg[31:0];
assign desc_2_axuser_14_axuser_f = desc_2_axuser_14_reg[31:0];
assign desc_2_axuser_15_axuser_f = desc_2_axuser_15_reg[31:0];
assign desc_2_size_txn_size_f = desc_2_size_reg[15:0];
assign desc_2_axsize_axsize_f = desc_2_axsize_reg[2:0];
assign desc_2_axaddr_0_addr_f = desc_2_axaddr_0_reg[31:0];
assign desc_2_axaddr_1_addr_f = desc_2_axaddr_1_reg[31:0];
assign desc_2_axaddr_2_addr_f = desc_2_axaddr_2_reg[31:0];
assign desc_2_axaddr_3_addr_f = desc_2_axaddr_3_reg[31:0];
assign desc_2_data_offset_addr_f = desc_2_data_offset_reg[31:0];
assign desc_2_wuser_0_wuser_f = desc_2_wuser_0_reg[31:0];
assign desc_2_wuser_1_wuser_f = desc_2_wuser_1_reg[31:0];
assign desc_2_wuser_2_wuser_f = desc_2_wuser_2_reg[31:0];
assign desc_2_wuser_3_wuser_f = desc_2_wuser_3_reg[31:0];
assign desc_2_wuser_4_wuser_f = desc_2_wuser_4_reg[31:0];
assign desc_2_wuser_5_wuser_f = desc_2_wuser_5_reg[31:0];
assign desc_2_wuser_6_wuser_f = desc_2_wuser_6_reg[31:0];
assign desc_2_wuser_7_wuser_f = desc_2_wuser_7_reg[31:0];
assign desc_2_wuser_8_wuser_f = desc_2_wuser_8_reg[31:0];
assign desc_2_wuser_9_wuser_f = desc_2_wuser_9_reg[31:0];
assign desc_2_wuser_10_wuser_f = desc_2_wuser_10_reg[31:0];
assign desc_2_wuser_11_wuser_f = desc_2_wuser_11_reg[31:0];
assign desc_2_wuser_12_wuser_f = desc_2_wuser_12_reg[31:0];
assign desc_2_wuser_13_wuser_f = desc_2_wuser_13_reg[31:0];
assign desc_2_wuser_14_wuser_f = desc_2_wuser_14_reg[31:0];
assign desc_2_wuser_15_wuser_f = desc_2_wuser_15_reg[31:0];
assign desc_2_data_host_addr_0_addr_f = desc_2_data_host_addr_0_reg[31:0];
assign desc_2_data_host_addr_1_addr_f = desc_2_data_host_addr_1_reg[31:0];
assign desc_2_data_host_addr_2_addr_f = desc_2_data_host_addr_2_reg[31:0];
assign desc_2_data_host_addr_3_addr_f = desc_2_data_host_addr_3_reg[31:0];
assign desc_2_wstrb_host_addr_0_addr_f = desc_2_wstrb_host_addr_0_reg[31:0];
assign desc_2_wstrb_host_addr_1_addr_f = desc_2_wstrb_host_addr_1_reg[31:0];
assign desc_2_wstrb_host_addr_2_addr_f = desc_2_wstrb_host_addr_2_reg[31:0];
assign desc_2_wstrb_host_addr_3_addr_f = desc_2_wstrb_host_addr_3_reg[31:0];
assign desc_2_xuser_0_xuser_f = desc_2_xuser_0_reg[31:0];
assign desc_2_xuser_1_xuser_f = desc_2_xuser_1_reg[31:0];
assign desc_2_xuser_2_xuser_f = desc_2_xuser_2_reg[31:0];
assign desc_2_xuser_3_xuser_f = desc_2_xuser_3_reg[31:0];
assign desc_2_xuser_4_xuser_f = desc_2_xuser_4_reg[31:0];
assign desc_2_xuser_5_xuser_f = desc_2_xuser_5_reg[31:0];
assign desc_2_xuser_6_xuser_f = desc_2_xuser_6_reg[31:0];
assign desc_2_xuser_7_xuser_f = desc_2_xuser_7_reg[31:0];
assign desc_2_xuser_8_xuser_f = desc_2_xuser_8_reg[31:0];
assign desc_2_xuser_9_xuser_f = desc_2_xuser_9_reg[31:0];
assign desc_2_xuser_10_xuser_f = desc_2_xuser_10_reg[31:0];
assign desc_2_xuser_11_xuser_f = desc_2_xuser_11_reg[31:0];
assign desc_2_xuser_12_xuser_f = desc_2_xuser_12_reg[31:0];
assign desc_2_xuser_13_xuser_f = desc_2_xuser_13_reg[31:0];
assign desc_2_xuser_14_xuser_f = desc_2_xuser_14_reg[31:0];
assign desc_2_xuser_15_xuser_f = desc_2_xuser_15_reg[31:0];
assign desc_3_txn_type_wr_strb_f = desc_3_txn_type_reg[1];
assign desc_3_txn_type_wr_rd_f = desc_3_txn_type_reg[0];
assign desc_3_attr_axregion_f = desc_3_attr_reg[18:15];
assign desc_3_attr_axqos_f = desc_3_attr_reg[14:11];
assign desc_3_attr_axprot_f = desc_3_attr_reg[10:8];
assign desc_3_attr_axcache_f = desc_3_attr_reg[7:4];
assign desc_3_attr_axlock_f = desc_3_attr_reg[3:2];
assign desc_3_attr_axburst_f = desc_3_attr_reg[1:0];
assign desc_3_axid_0_axid_f = desc_3_axid_0_reg[31:0];
assign desc_3_axid_1_axid_f = desc_3_axid_1_reg[31:0];
assign desc_3_axid_2_axid_f = desc_3_axid_2_reg[31:0];
assign desc_3_axid_3_axid_f = desc_3_axid_3_reg[31:0];
assign desc_3_axuser_0_axuser_f = desc_3_axuser_0_reg[31:0];
assign desc_3_axuser_1_axuser_f = desc_3_axuser_1_reg[31:0];
assign desc_3_axuser_2_axuser_f = desc_3_axuser_2_reg[31:0];
assign desc_3_axuser_3_axuser_f = desc_3_axuser_3_reg[31:0];
assign desc_3_axuser_4_axuser_f = desc_3_axuser_4_reg[31:0];
assign desc_3_axuser_5_axuser_f = desc_3_axuser_5_reg[31:0];
assign desc_3_axuser_6_axuser_f = desc_3_axuser_6_reg[31:0];
assign desc_3_axuser_7_axuser_f = desc_3_axuser_7_reg[31:0];
assign desc_3_axuser_8_axuser_f = desc_3_axuser_8_reg[31:0];
assign desc_3_axuser_9_axuser_f = desc_3_axuser_9_reg[31:0];
assign desc_3_axuser_10_axuser_f = desc_3_axuser_10_reg[31:0];
assign desc_3_axuser_11_axuser_f = desc_3_axuser_11_reg[31:0];
assign desc_3_axuser_12_axuser_f = desc_3_axuser_12_reg[31:0];
assign desc_3_axuser_13_axuser_f = desc_3_axuser_13_reg[31:0];
assign desc_3_axuser_14_axuser_f = desc_3_axuser_14_reg[31:0];
assign desc_3_axuser_15_axuser_f = desc_3_axuser_15_reg[31:0];
assign desc_3_size_txn_size_f = desc_3_size_reg[15:0];
assign desc_3_axsize_axsize_f = desc_3_axsize_reg[2:0];
assign desc_3_axaddr_0_addr_f = desc_3_axaddr_0_reg[31:0];
assign desc_3_axaddr_1_addr_f = desc_3_axaddr_1_reg[31:0];
assign desc_3_axaddr_2_addr_f = desc_3_axaddr_2_reg[31:0];
assign desc_3_axaddr_3_addr_f = desc_3_axaddr_3_reg[31:0];
assign desc_3_data_offset_addr_f = desc_3_data_offset_reg[31:0];
assign desc_3_wuser_0_wuser_f = desc_3_wuser_0_reg[31:0];
assign desc_3_wuser_1_wuser_f = desc_3_wuser_1_reg[31:0];
assign desc_3_wuser_2_wuser_f = desc_3_wuser_2_reg[31:0];
assign desc_3_wuser_3_wuser_f = desc_3_wuser_3_reg[31:0];
assign desc_3_wuser_4_wuser_f = desc_3_wuser_4_reg[31:0];
assign desc_3_wuser_5_wuser_f = desc_3_wuser_5_reg[31:0];
assign desc_3_wuser_6_wuser_f = desc_3_wuser_6_reg[31:0];
assign desc_3_wuser_7_wuser_f = desc_3_wuser_7_reg[31:0];
assign desc_3_wuser_8_wuser_f = desc_3_wuser_8_reg[31:0];
assign desc_3_wuser_9_wuser_f = desc_3_wuser_9_reg[31:0];
assign desc_3_wuser_10_wuser_f = desc_3_wuser_10_reg[31:0];
assign desc_3_wuser_11_wuser_f = desc_3_wuser_11_reg[31:0];
assign desc_3_wuser_12_wuser_f = desc_3_wuser_12_reg[31:0];
assign desc_3_wuser_13_wuser_f = desc_3_wuser_13_reg[31:0];
assign desc_3_wuser_14_wuser_f = desc_3_wuser_14_reg[31:0];
assign desc_3_wuser_15_wuser_f = desc_3_wuser_15_reg[31:0];
assign desc_3_data_host_addr_0_addr_f = desc_3_data_host_addr_0_reg[31:0];
assign desc_3_data_host_addr_1_addr_f = desc_3_data_host_addr_1_reg[31:0];
assign desc_3_data_host_addr_2_addr_f = desc_3_data_host_addr_2_reg[31:0];
assign desc_3_data_host_addr_3_addr_f = desc_3_data_host_addr_3_reg[31:0];
assign desc_3_wstrb_host_addr_0_addr_f = desc_3_wstrb_host_addr_0_reg[31:0];
assign desc_3_wstrb_host_addr_1_addr_f = desc_3_wstrb_host_addr_1_reg[31:0];
assign desc_3_wstrb_host_addr_2_addr_f = desc_3_wstrb_host_addr_2_reg[31:0];
assign desc_3_wstrb_host_addr_3_addr_f = desc_3_wstrb_host_addr_3_reg[31:0];
assign desc_3_xuser_0_xuser_f = desc_3_xuser_0_reg[31:0];
assign desc_3_xuser_1_xuser_f = desc_3_xuser_1_reg[31:0];
assign desc_3_xuser_2_xuser_f = desc_3_xuser_2_reg[31:0];
assign desc_3_xuser_3_xuser_f = desc_3_xuser_3_reg[31:0];
assign desc_3_xuser_4_xuser_f = desc_3_xuser_4_reg[31:0];
assign desc_3_xuser_5_xuser_f = desc_3_xuser_5_reg[31:0];
assign desc_3_xuser_6_xuser_f = desc_3_xuser_6_reg[31:0];
assign desc_3_xuser_7_xuser_f = desc_3_xuser_7_reg[31:0];
assign desc_3_xuser_8_xuser_f = desc_3_xuser_8_reg[31:0];
assign desc_3_xuser_9_xuser_f = desc_3_xuser_9_reg[31:0];
assign desc_3_xuser_10_xuser_f = desc_3_xuser_10_reg[31:0];
assign desc_3_xuser_11_xuser_f = desc_3_xuser_11_reg[31:0];
assign desc_3_xuser_12_xuser_f = desc_3_xuser_12_reg[31:0];
assign desc_3_xuser_13_xuser_f = desc_3_xuser_13_reg[31:0];
assign desc_3_xuser_14_xuser_f = desc_3_xuser_14_reg[31:0];
assign desc_3_xuser_15_xuser_f = desc_3_xuser_15_reg[31:0];
assign desc_4_txn_type_wr_strb_f = desc_4_txn_type_reg[1];
assign desc_4_txn_type_wr_rd_f = desc_4_txn_type_reg[0];
assign desc_4_attr_axregion_f = desc_4_attr_reg[18:15];
assign desc_4_attr_axqos_f = desc_4_attr_reg[14:11];
assign desc_4_attr_axprot_f = desc_4_attr_reg[10:8];
assign desc_4_attr_axcache_f = desc_4_attr_reg[7:4];
assign desc_4_attr_axlock_f = desc_4_attr_reg[3:2];
assign desc_4_attr_axburst_f = desc_4_attr_reg[1:0];
assign desc_4_axid_0_axid_f = desc_4_axid_0_reg[31:0];
assign desc_4_axid_1_axid_f = desc_4_axid_1_reg[31:0];
assign desc_4_axid_2_axid_f = desc_4_axid_2_reg[31:0];
assign desc_4_axid_3_axid_f = desc_4_axid_3_reg[31:0];
assign desc_4_axuser_0_axuser_f = desc_4_axuser_0_reg[31:0];
assign desc_4_axuser_1_axuser_f = desc_4_axuser_1_reg[31:0];
assign desc_4_axuser_2_axuser_f = desc_4_axuser_2_reg[31:0];
assign desc_4_axuser_3_axuser_f = desc_4_axuser_3_reg[31:0];
assign desc_4_axuser_4_axuser_f = desc_4_axuser_4_reg[31:0];
assign desc_4_axuser_5_axuser_f = desc_4_axuser_5_reg[31:0];
assign desc_4_axuser_6_axuser_f = desc_4_axuser_6_reg[31:0];
assign desc_4_axuser_7_axuser_f = desc_4_axuser_7_reg[31:0];
assign desc_4_axuser_8_axuser_f = desc_4_axuser_8_reg[31:0];
assign desc_4_axuser_9_axuser_f = desc_4_axuser_9_reg[31:0];
assign desc_4_axuser_10_axuser_f = desc_4_axuser_10_reg[31:0];
assign desc_4_axuser_11_axuser_f = desc_4_axuser_11_reg[31:0];
assign desc_4_axuser_12_axuser_f = desc_4_axuser_12_reg[31:0];
assign desc_4_axuser_13_axuser_f = desc_4_axuser_13_reg[31:0];
assign desc_4_axuser_14_axuser_f = desc_4_axuser_14_reg[31:0];
assign desc_4_axuser_15_axuser_f = desc_4_axuser_15_reg[31:0];
assign desc_4_size_txn_size_f = desc_4_size_reg[15:0];
assign desc_4_axsize_axsize_f = desc_4_axsize_reg[2:0];
assign desc_4_axaddr_0_addr_f = desc_4_axaddr_0_reg[31:0];
assign desc_4_axaddr_1_addr_f = desc_4_axaddr_1_reg[31:0];
assign desc_4_axaddr_2_addr_f = desc_4_axaddr_2_reg[31:0];
assign desc_4_axaddr_3_addr_f = desc_4_axaddr_3_reg[31:0];
assign desc_4_data_offset_addr_f = desc_4_data_offset_reg[31:0];
assign desc_4_wuser_0_wuser_f = desc_4_wuser_0_reg[31:0];
assign desc_4_wuser_1_wuser_f = desc_4_wuser_1_reg[31:0];
assign desc_4_wuser_2_wuser_f = desc_4_wuser_2_reg[31:0];
assign desc_4_wuser_3_wuser_f = desc_4_wuser_3_reg[31:0];
assign desc_4_wuser_4_wuser_f = desc_4_wuser_4_reg[31:0];
assign desc_4_wuser_5_wuser_f = desc_4_wuser_5_reg[31:0];
assign desc_4_wuser_6_wuser_f = desc_4_wuser_6_reg[31:0];
assign desc_4_wuser_7_wuser_f = desc_4_wuser_7_reg[31:0];
assign desc_4_wuser_8_wuser_f = desc_4_wuser_8_reg[31:0];
assign desc_4_wuser_9_wuser_f = desc_4_wuser_9_reg[31:0];
assign desc_4_wuser_10_wuser_f = desc_4_wuser_10_reg[31:0];
assign desc_4_wuser_11_wuser_f = desc_4_wuser_11_reg[31:0];
assign desc_4_wuser_12_wuser_f = desc_4_wuser_12_reg[31:0];
assign desc_4_wuser_13_wuser_f = desc_4_wuser_13_reg[31:0];
assign desc_4_wuser_14_wuser_f = desc_4_wuser_14_reg[31:0];
assign desc_4_wuser_15_wuser_f = desc_4_wuser_15_reg[31:0];
assign desc_4_data_host_addr_0_addr_f = desc_4_data_host_addr_0_reg[31:0];
assign desc_4_data_host_addr_1_addr_f = desc_4_data_host_addr_1_reg[31:0];
assign desc_4_data_host_addr_2_addr_f = desc_4_data_host_addr_2_reg[31:0];
assign desc_4_data_host_addr_3_addr_f = desc_4_data_host_addr_3_reg[31:0];
assign desc_4_wstrb_host_addr_0_addr_f = desc_4_wstrb_host_addr_0_reg[31:0];
assign desc_4_wstrb_host_addr_1_addr_f = desc_4_wstrb_host_addr_1_reg[31:0];
assign desc_4_wstrb_host_addr_2_addr_f = desc_4_wstrb_host_addr_2_reg[31:0];
assign desc_4_wstrb_host_addr_3_addr_f = desc_4_wstrb_host_addr_3_reg[31:0];
assign desc_4_xuser_0_xuser_f = desc_4_xuser_0_reg[31:0];
assign desc_4_xuser_1_xuser_f = desc_4_xuser_1_reg[31:0];
assign desc_4_xuser_2_xuser_f = desc_4_xuser_2_reg[31:0];
assign desc_4_xuser_3_xuser_f = desc_4_xuser_3_reg[31:0];
assign desc_4_xuser_4_xuser_f = desc_4_xuser_4_reg[31:0];
assign desc_4_xuser_5_xuser_f = desc_4_xuser_5_reg[31:0];
assign desc_4_xuser_6_xuser_f = desc_4_xuser_6_reg[31:0];
assign desc_4_xuser_7_xuser_f = desc_4_xuser_7_reg[31:0];
assign desc_4_xuser_8_xuser_f = desc_4_xuser_8_reg[31:0];
assign desc_4_xuser_9_xuser_f = desc_4_xuser_9_reg[31:0];
assign desc_4_xuser_10_xuser_f = desc_4_xuser_10_reg[31:0];
assign desc_4_xuser_11_xuser_f = desc_4_xuser_11_reg[31:0];
assign desc_4_xuser_12_xuser_f = desc_4_xuser_12_reg[31:0];
assign desc_4_xuser_13_xuser_f = desc_4_xuser_13_reg[31:0];
assign desc_4_xuser_14_xuser_f = desc_4_xuser_14_reg[31:0];
assign desc_4_xuser_15_xuser_f = desc_4_xuser_15_reg[31:0];
assign desc_5_txn_type_wr_strb_f = desc_5_txn_type_reg[1];
assign desc_5_txn_type_wr_rd_f = desc_5_txn_type_reg[0];
assign desc_5_attr_axregion_f = desc_5_attr_reg[18:15];
assign desc_5_attr_axqos_f = desc_5_attr_reg[14:11];
assign desc_5_attr_axprot_f = desc_5_attr_reg[10:8];
assign desc_5_attr_axcache_f = desc_5_attr_reg[7:4];
assign desc_5_attr_axlock_f = desc_5_attr_reg[3:2];
assign desc_5_attr_axburst_f = desc_5_attr_reg[1:0];
assign desc_5_axid_0_axid_f = desc_5_axid_0_reg[31:0];
assign desc_5_axid_1_axid_f = desc_5_axid_1_reg[31:0];
assign desc_5_axid_2_axid_f = desc_5_axid_2_reg[31:0];
assign desc_5_axid_3_axid_f = desc_5_axid_3_reg[31:0];
assign desc_5_axuser_0_axuser_f = desc_5_axuser_0_reg[31:0];
assign desc_5_axuser_1_axuser_f = desc_5_axuser_1_reg[31:0];
assign desc_5_axuser_2_axuser_f = desc_5_axuser_2_reg[31:0];
assign desc_5_axuser_3_axuser_f = desc_5_axuser_3_reg[31:0];
assign desc_5_axuser_4_axuser_f = desc_5_axuser_4_reg[31:0];
assign desc_5_axuser_5_axuser_f = desc_5_axuser_5_reg[31:0];
assign desc_5_axuser_6_axuser_f = desc_5_axuser_6_reg[31:0];
assign desc_5_axuser_7_axuser_f = desc_5_axuser_7_reg[31:0];
assign desc_5_axuser_8_axuser_f = desc_5_axuser_8_reg[31:0];
assign desc_5_axuser_9_axuser_f = desc_5_axuser_9_reg[31:0];
assign desc_5_axuser_10_axuser_f = desc_5_axuser_10_reg[31:0];
assign desc_5_axuser_11_axuser_f = desc_5_axuser_11_reg[31:0];
assign desc_5_axuser_12_axuser_f = desc_5_axuser_12_reg[31:0];
assign desc_5_axuser_13_axuser_f = desc_5_axuser_13_reg[31:0];
assign desc_5_axuser_14_axuser_f = desc_5_axuser_14_reg[31:0];
assign desc_5_axuser_15_axuser_f = desc_5_axuser_15_reg[31:0];
assign desc_5_size_txn_size_f = desc_5_size_reg[15:0];
assign desc_5_axsize_axsize_f = desc_5_axsize_reg[2:0];
assign desc_5_axaddr_0_addr_f = desc_5_axaddr_0_reg[31:0];
assign desc_5_axaddr_1_addr_f = desc_5_axaddr_1_reg[31:0];
assign desc_5_axaddr_2_addr_f = desc_5_axaddr_2_reg[31:0];
assign desc_5_axaddr_3_addr_f = desc_5_axaddr_3_reg[31:0];
assign desc_5_data_offset_addr_f = desc_5_data_offset_reg[31:0];
assign desc_5_wuser_0_wuser_f = desc_5_wuser_0_reg[31:0];
assign desc_5_wuser_1_wuser_f = desc_5_wuser_1_reg[31:0];
assign desc_5_wuser_2_wuser_f = desc_5_wuser_2_reg[31:0];
assign desc_5_wuser_3_wuser_f = desc_5_wuser_3_reg[31:0];
assign desc_5_wuser_4_wuser_f = desc_5_wuser_4_reg[31:0];
assign desc_5_wuser_5_wuser_f = desc_5_wuser_5_reg[31:0];
assign desc_5_wuser_6_wuser_f = desc_5_wuser_6_reg[31:0];
assign desc_5_wuser_7_wuser_f = desc_5_wuser_7_reg[31:0];
assign desc_5_wuser_8_wuser_f = desc_5_wuser_8_reg[31:0];
assign desc_5_wuser_9_wuser_f = desc_5_wuser_9_reg[31:0];
assign desc_5_wuser_10_wuser_f = desc_5_wuser_10_reg[31:0];
assign desc_5_wuser_11_wuser_f = desc_5_wuser_11_reg[31:0];
assign desc_5_wuser_12_wuser_f = desc_5_wuser_12_reg[31:0];
assign desc_5_wuser_13_wuser_f = desc_5_wuser_13_reg[31:0];
assign desc_5_wuser_14_wuser_f = desc_5_wuser_14_reg[31:0];
assign desc_5_wuser_15_wuser_f = desc_5_wuser_15_reg[31:0];
assign desc_5_data_host_addr_0_addr_f = desc_5_data_host_addr_0_reg[31:0];
assign desc_5_data_host_addr_1_addr_f = desc_5_data_host_addr_1_reg[31:0];
assign desc_5_data_host_addr_2_addr_f = desc_5_data_host_addr_2_reg[31:0];
assign desc_5_data_host_addr_3_addr_f = desc_5_data_host_addr_3_reg[31:0];
assign desc_5_wstrb_host_addr_0_addr_f = desc_5_wstrb_host_addr_0_reg[31:0];
assign desc_5_wstrb_host_addr_1_addr_f = desc_5_wstrb_host_addr_1_reg[31:0];
assign desc_5_wstrb_host_addr_2_addr_f = desc_5_wstrb_host_addr_2_reg[31:0];
assign desc_5_wstrb_host_addr_3_addr_f = desc_5_wstrb_host_addr_3_reg[31:0];
assign desc_5_xuser_0_xuser_f = desc_5_xuser_0_reg[31:0];
assign desc_5_xuser_1_xuser_f = desc_5_xuser_1_reg[31:0];
assign desc_5_xuser_2_xuser_f = desc_5_xuser_2_reg[31:0];
assign desc_5_xuser_3_xuser_f = desc_5_xuser_3_reg[31:0];
assign desc_5_xuser_4_xuser_f = desc_5_xuser_4_reg[31:0];
assign desc_5_xuser_5_xuser_f = desc_5_xuser_5_reg[31:0];
assign desc_5_xuser_6_xuser_f = desc_5_xuser_6_reg[31:0];
assign desc_5_xuser_7_xuser_f = desc_5_xuser_7_reg[31:0];
assign desc_5_xuser_8_xuser_f = desc_5_xuser_8_reg[31:0];
assign desc_5_xuser_9_xuser_f = desc_5_xuser_9_reg[31:0];
assign desc_5_xuser_10_xuser_f = desc_5_xuser_10_reg[31:0];
assign desc_5_xuser_11_xuser_f = desc_5_xuser_11_reg[31:0];
assign desc_5_xuser_12_xuser_f = desc_5_xuser_12_reg[31:0];
assign desc_5_xuser_13_xuser_f = desc_5_xuser_13_reg[31:0];
assign desc_5_xuser_14_xuser_f = desc_5_xuser_14_reg[31:0];
assign desc_5_xuser_15_xuser_f = desc_5_xuser_15_reg[31:0];
assign desc_6_txn_type_wr_strb_f = desc_6_txn_type_reg[1];
assign desc_6_txn_type_wr_rd_f = desc_6_txn_type_reg[0];
assign desc_6_attr_axregion_f = desc_6_attr_reg[18:15];
assign desc_6_attr_axqos_f = desc_6_attr_reg[14:11];
assign desc_6_attr_axprot_f = desc_6_attr_reg[10:8];
assign desc_6_attr_axcache_f = desc_6_attr_reg[7:4];
assign desc_6_attr_axlock_f = desc_6_attr_reg[3:2];
assign desc_6_attr_axburst_f = desc_6_attr_reg[1:0];
assign desc_6_axid_0_axid_f = desc_6_axid_0_reg[31:0];
assign desc_6_axid_1_axid_f = desc_6_axid_1_reg[31:0];
assign desc_6_axid_2_axid_f = desc_6_axid_2_reg[31:0];
assign desc_6_axid_3_axid_f = desc_6_axid_3_reg[31:0];
assign desc_6_axuser_0_axuser_f = desc_6_axuser_0_reg[31:0];
assign desc_6_axuser_1_axuser_f = desc_6_axuser_1_reg[31:0];
assign desc_6_axuser_2_axuser_f = desc_6_axuser_2_reg[31:0];
assign desc_6_axuser_3_axuser_f = desc_6_axuser_3_reg[31:0];
assign desc_6_axuser_4_axuser_f = desc_6_axuser_4_reg[31:0];
assign desc_6_axuser_5_axuser_f = desc_6_axuser_5_reg[31:0];
assign desc_6_axuser_6_axuser_f = desc_6_axuser_6_reg[31:0];
assign desc_6_axuser_7_axuser_f = desc_6_axuser_7_reg[31:0];
assign desc_6_axuser_8_axuser_f = desc_6_axuser_8_reg[31:0];
assign desc_6_axuser_9_axuser_f = desc_6_axuser_9_reg[31:0];
assign desc_6_axuser_10_axuser_f = desc_6_axuser_10_reg[31:0];
assign desc_6_axuser_11_axuser_f = desc_6_axuser_11_reg[31:0];
assign desc_6_axuser_12_axuser_f = desc_6_axuser_12_reg[31:0];
assign desc_6_axuser_13_axuser_f = desc_6_axuser_13_reg[31:0];
assign desc_6_axuser_14_axuser_f = desc_6_axuser_14_reg[31:0];
assign desc_6_axuser_15_axuser_f = desc_6_axuser_15_reg[31:0];
assign desc_6_size_txn_size_f = desc_6_size_reg[15:0];
assign desc_6_axsize_axsize_f = desc_6_axsize_reg[2:0];
assign desc_6_axaddr_0_addr_f = desc_6_axaddr_0_reg[31:0];
assign desc_6_axaddr_1_addr_f = desc_6_axaddr_1_reg[31:0];
assign desc_6_axaddr_2_addr_f = desc_6_axaddr_2_reg[31:0];
assign desc_6_axaddr_3_addr_f = desc_6_axaddr_3_reg[31:0];
assign desc_6_data_offset_addr_f = desc_6_data_offset_reg[31:0];
assign desc_6_wuser_0_wuser_f = desc_6_wuser_0_reg[31:0];
assign desc_6_wuser_1_wuser_f = desc_6_wuser_1_reg[31:0];
assign desc_6_wuser_2_wuser_f = desc_6_wuser_2_reg[31:0];
assign desc_6_wuser_3_wuser_f = desc_6_wuser_3_reg[31:0];
assign desc_6_wuser_4_wuser_f = desc_6_wuser_4_reg[31:0];
assign desc_6_wuser_5_wuser_f = desc_6_wuser_5_reg[31:0];
assign desc_6_wuser_6_wuser_f = desc_6_wuser_6_reg[31:0];
assign desc_6_wuser_7_wuser_f = desc_6_wuser_7_reg[31:0];
assign desc_6_wuser_8_wuser_f = desc_6_wuser_8_reg[31:0];
assign desc_6_wuser_9_wuser_f = desc_6_wuser_9_reg[31:0];
assign desc_6_wuser_10_wuser_f = desc_6_wuser_10_reg[31:0];
assign desc_6_wuser_11_wuser_f = desc_6_wuser_11_reg[31:0];
assign desc_6_wuser_12_wuser_f = desc_6_wuser_12_reg[31:0];
assign desc_6_wuser_13_wuser_f = desc_6_wuser_13_reg[31:0];
assign desc_6_wuser_14_wuser_f = desc_6_wuser_14_reg[31:0];
assign desc_6_wuser_15_wuser_f = desc_6_wuser_15_reg[31:0];
assign desc_6_data_host_addr_0_addr_f = desc_6_data_host_addr_0_reg[31:0];
assign desc_6_data_host_addr_1_addr_f = desc_6_data_host_addr_1_reg[31:0];
assign desc_6_data_host_addr_2_addr_f = desc_6_data_host_addr_2_reg[31:0];
assign desc_6_data_host_addr_3_addr_f = desc_6_data_host_addr_3_reg[31:0];
assign desc_6_wstrb_host_addr_0_addr_f = desc_6_wstrb_host_addr_0_reg[31:0];
assign desc_6_wstrb_host_addr_1_addr_f = desc_6_wstrb_host_addr_1_reg[31:0];
assign desc_6_wstrb_host_addr_2_addr_f = desc_6_wstrb_host_addr_2_reg[31:0];
assign desc_6_wstrb_host_addr_3_addr_f = desc_6_wstrb_host_addr_3_reg[31:0];
assign desc_6_xuser_0_xuser_f = desc_6_xuser_0_reg[31:0];
assign desc_6_xuser_1_xuser_f = desc_6_xuser_1_reg[31:0];
assign desc_6_xuser_2_xuser_f = desc_6_xuser_2_reg[31:0];
assign desc_6_xuser_3_xuser_f = desc_6_xuser_3_reg[31:0];
assign desc_6_xuser_4_xuser_f = desc_6_xuser_4_reg[31:0];
assign desc_6_xuser_5_xuser_f = desc_6_xuser_5_reg[31:0];
assign desc_6_xuser_6_xuser_f = desc_6_xuser_6_reg[31:0];
assign desc_6_xuser_7_xuser_f = desc_6_xuser_7_reg[31:0];
assign desc_6_xuser_8_xuser_f = desc_6_xuser_8_reg[31:0];
assign desc_6_xuser_9_xuser_f = desc_6_xuser_9_reg[31:0];
assign desc_6_xuser_10_xuser_f = desc_6_xuser_10_reg[31:0];
assign desc_6_xuser_11_xuser_f = desc_6_xuser_11_reg[31:0];
assign desc_6_xuser_12_xuser_f = desc_6_xuser_12_reg[31:0];
assign desc_6_xuser_13_xuser_f = desc_6_xuser_13_reg[31:0];
assign desc_6_xuser_14_xuser_f = desc_6_xuser_14_reg[31:0];
assign desc_6_xuser_15_xuser_f = desc_6_xuser_15_reg[31:0];
assign desc_7_txn_type_wr_strb_f = desc_7_txn_type_reg[1];
assign desc_7_txn_type_wr_rd_f = desc_7_txn_type_reg[0];
assign desc_7_attr_axregion_f = desc_7_attr_reg[18:15];
assign desc_7_attr_axqos_f = desc_7_attr_reg[14:11];
assign desc_7_attr_axprot_f = desc_7_attr_reg[10:8];
assign desc_7_attr_axcache_f = desc_7_attr_reg[7:4];
assign desc_7_attr_axlock_f = desc_7_attr_reg[3:2];
assign desc_7_attr_axburst_f = desc_7_attr_reg[1:0];
assign desc_7_axid_0_axid_f = desc_7_axid_0_reg[31:0];
assign desc_7_axid_1_axid_f = desc_7_axid_1_reg[31:0];
assign desc_7_axid_2_axid_f = desc_7_axid_2_reg[31:0];
assign desc_7_axid_3_axid_f = desc_7_axid_3_reg[31:0];
assign desc_7_axuser_0_axuser_f = desc_7_axuser_0_reg[31:0];
assign desc_7_axuser_1_axuser_f = desc_7_axuser_1_reg[31:0];
assign desc_7_axuser_2_axuser_f = desc_7_axuser_2_reg[31:0];
assign desc_7_axuser_3_axuser_f = desc_7_axuser_3_reg[31:0];
assign desc_7_axuser_4_axuser_f = desc_7_axuser_4_reg[31:0];
assign desc_7_axuser_5_axuser_f = desc_7_axuser_5_reg[31:0];
assign desc_7_axuser_6_axuser_f = desc_7_axuser_6_reg[31:0];
assign desc_7_axuser_7_axuser_f = desc_7_axuser_7_reg[31:0];
assign desc_7_axuser_8_axuser_f = desc_7_axuser_8_reg[31:0];
assign desc_7_axuser_9_axuser_f = desc_7_axuser_9_reg[31:0];
assign desc_7_axuser_10_axuser_f = desc_7_axuser_10_reg[31:0];
assign desc_7_axuser_11_axuser_f = desc_7_axuser_11_reg[31:0];
assign desc_7_axuser_12_axuser_f = desc_7_axuser_12_reg[31:0];
assign desc_7_axuser_13_axuser_f = desc_7_axuser_13_reg[31:0];
assign desc_7_axuser_14_axuser_f = desc_7_axuser_14_reg[31:0];
assign desc_7_axuser_15_axuser_f = desc_7_axuser_15_reg[31:0];
assign desc_7_size_txn_size_f = desc_7_size_reg[15:0];
assign desc_7_axsize_axsize_f = desc_7_axsize_reg[2:0];
assign desc_7_axaddr_0_addr_f = desc_7_axaddr_0_reg[31:0];
assign desc_7_axaddr_1_addr_f = desc_7_axaddr_1_reg[31:0];
assign desc_7_axaddr_2_addr_f = desc_7_axaddr_2_reg[31:0];
assign desc_7_axaddr_3_addr_f = desc_7_axaddr_3_reg[31:0];
assign desc_7_data_offset_addr_f = desc_7_data_offset_reg[31:0];
assign desc_7_wuser_0_wuser_f = desc_7_wuser_0_reg[31:0];
assign desc_7_wuser_1_wuser_f = desc_7_wuser_1_reg[31:0];
assign desc_7_wuser_2_wuser_f = desc_7_wuser_2_reg[31:0];
assign desc_7_wuser_3_wuser_f = desc_7_wuser_3_reg[31:0];
assign desc_7_wuser_4_wuser_f = desc_7_wuser_4_reg[31:0];
assign desc_7_wuser_5_wuser_f = desc_7_wuser_5_reg[31:0];
assign desc_7_wuser_6_wuser_f = desc_7_wuser_6_reg[31:0];
assign desc_7_wuser_7_wuser_f = desc_7_wuser_7_reg[31:0];
assign desc_7_wuser_8_wuser_f = desc_7_wuser_8_reg[31:0];
assign desc_7_wuser_9_wuser_f = desc_7_wuser_9_reg[31:0];
assign desc_7_wuser_10_wuser_f = desc_7_wuser_10_reg[31:0];
assign desc_7_wuser_11_wuser_f = desc_7_wuser_11_reg[31:0];
assign desc_7_wuser_12_wuser_f = desc_7_wuser_12_reg[31:0];
assign desc_7_wuser_13_wuser_f = desc_7_wuser_13_reg[31:0];
assign desc_7_wuser_14_wuser_f = desc_7_wuser_14_reg[31:0];
assign desc_7_wuser_15_wuser_f = desc_7_wuser_15_reg[31:0];
assign desc_7_data_host_addr_0_addr_f = desc_7_data_host_addr_0_reg[31:0];
assign desc_7_data_host_addr_1_addr_f = desc_7_data_host_addr_1_reg[31:0];
assign desc_7_data_host_addr_2_addr_f = desc_7_data_host_addr_2_reg[31:0];
assign desc_7_data_host_addr_3_addr_f = desc_7_data_host_addr_3_reg[31:0];
assign desc_7_wstrb_host_addr_0_addr_f = desc_7_wstrb_host_addr_0_reg[31:0];
assign desc_7_wstrb_host_addr_1_addr_f = desc_7_wstrb_host_addr_1_reg[31:0];
assign desc_7_wstrb_host_addr_2_addr_f = desc_7_wstrb_host_addr_2_reg[31:0];
assign desc_7_wstrb_host_addr_3_addr_f = desc_7_wstrb_host_addr_3_reg[31:0];
assign desc_7_xuser_0_xuser_f = desc_7_xuser_0_reg[31:0];
assign desc_7_xuser_1_xuser_f = desc_7_xuser_1_reg[31:0];
assign desc_7_xuser_2_xuser_f = desc_7_xuser_2_reg[31:0];
assign desc_7_xuser_3_xuser_f = desc_7_xuser_3_reg[31:0];
assign desc_7_xuser_4_xuser_f = desc_7_xuser_4_reg[31:0];
assign desc_7_xuser_5_xuser_f = desc_7_xuser_5_reg[31:0];
assign desc_7_xuser_6_xuser_f = desc_7_xuser_6_reg[31:0];
assign desc_7_xuser_7_xuser_f = desc_7_xuser_7_reg[31:0];
assign desc_7_xuser_8_xuser_f = desc_7_xuser_8_reg[31:0];
assign desc_7_xuser_9_xuser_f = desc_7_xuser_9_reg[31:0];
assign desc_7_xuser_10_xuser_f = desc_7_xuser_10_reg[31:0];
assign desc_7_xuser_11_xuser_f = desc_7_xuser_11_reg[31:0];
assign desc_7_xuser_12_xuser_f = desc_7_xuser_12_reg[31:0];
assign desc_7_xuser_13_xuser_f = desc_7_xuser_13_reg[31:0];
assign desc_7_xuser_14_xuser_f = desc_7_xuser_14_reg[31:0];
assign desc_7_xuser_15_xuser_f = desc_7_xuser_15_reg[31:0];
assign desc_8_txn_type_wr_strb_f = desc_8_txn_type_reg[1];
assign desc_8_txn_type_wr_rd_f = desc_8_txn_type_reg[0];
assign desc_8_attr_axregion_f = desc_8_attr_reg[18:15];
assign desc_8_attr_axqos_f = desc_8_attr_reg[14:11];
assign desc_8_attr_axprot_f = desc_8_attr_reg[10:8];
assign desc_8_attr_axcache_f = desc_8_attr_reg[7:4];
assign desc_8_attr_axlock_f = desc_8_attr_reg[3:2];
assign desc_8_attr_axburst_f = desc_8_attr_reg[1:0];
assign desc_8_axid_0_axid_f = desc_8_axid_0_reg[31:0];
assign desc_8_axid_1_axid_f = desc_8_axid_1_reg[31:0];
assign desc_8_axid_2_axid_f = desc_8_axid_2_reg[31:0];
assign desc_8_axid_3_axid_f = desc_8_axid_3_reg[31:0];
assign desc_8_axuser_0_axuser_f = desc_8_axuser_0_reg[31:0];
assign desc_8_axuser_1_axuser_f = desc_8_axuser_1_reg[31:0];
assign desc_8_axuser_2_axuser_f = desc_8_axuser_2_reg[31:0];
assign desc_8_axuser_3_axuser_f = desc_8_axuser_3_reg[31:0];
assign desc_8_axuser_4_axuser_f = desc_8_axuser_4_reg[31:0];
assign desc_8_axuser_5_axuser_f = desc_8_axuser_5_reg[31:0];
assign desc_8_axuser_6_axuser_f = desc_8_axuser_6_reg[31:0];
assign desc_8_axuser_7_axuser_f = desc_8_axuser_7_reg[31:0];
assign desc_8_axuser_8_axuser_f = desc_8_axuser_8_reg[31:0];
assign desc_8_axuser_9_axuser_f = desc_8_axuser_9_reg[31:0];
assign desc_8_axuser_10_axuser_f = desc_8_axuser_10_reg[31:0];
assign desc_8_axuser_11_axuser_f = desc_8_axuser_11_reg[31:0];
assign desc_8_axuser_12_axuser_f = desc_8_axuser_12_reg[31:0];
assign desc_8_axuser_13_axuser_f = desc_8_axuser_13_reg[31:0];
assign desc_8_axuser_14_axuser_f = desc_8_axuser_14_reg[31:0];
assign desc_8_axuser_15_axuser_f = desc_8_axuser_15_reg[31:0];
assign desc_8_size_txn_size_f = desc_8_size_reg[15:0];
assign desc_8_axsize_axsize_f = desc_8_axsize_reg[2:0];
assign desc_8_axaddr_0_addr_f = desc_8_axaddr_0_reg[31:0];
assign desc_8_axaddr_1_addr_f = desc_8_axaddr_1_reg[31:0];
assign desc_8_axaddr_2_addr_f = desc_8_axaddr_2_reg[31:0];
assign desc_8_axaddr_3_addr_f = desc_8_axaddr_3_reg[31:0];
assign desc_8_data_offset_addr_f = desc_8_data_offset_reg[31:0];
assign desc_8_wuser_0_wuser_f = desc_8_wuser_0_reg[31:0];
assign desc_8_wuser_1_wuser_f = desc_8_wuser_1_reg[31:0];
assign desc_8_wuser_2_wuser_f = desc_8_wuser_2_reg[31:0];
assign desc_8_wuser_3_wuser_f = desc_8_wuser_3_reg[31:0];
assign desc_8_wuser_4_wuser_f = desc_8_wuser_4_reg[31:0];
assign desc_8_wuser_5_wuser_f = desc_8_wuser_5_reg[31:0];
assign desc_8_wuser_6_wuser_f = desc_8_wuser_6_reg[31:0];
assign desc_8_wuser_7_wuser_f = desc_8_wuser_7_reg[31:0];
assign desc_8_wuser_8_wuser_f = desc_8_wuser_8_reg[31:0];
assign desc_8_wuser_9_wuser_f = desc_8_wuser_9_reg[31:0];
assign desc_8_wuser_10_wuser_f = desc_8_wuser_10_reg[31:0];
assign desc_8_wuser_11_wuser_f = desc_8_wuser_11_reg[31:0];
assign desc_8_wuser_12_wuser_f = desc_8_wuser_12_reg[31:0];
assign desc_8_wuser_13_wuser_f = desc_8_wuser_13_reg[31:0];
assign desc_8_wuser_14_wuser_f = desc_8_wuser_14_reg[31:0];
assign desc_8_wuser_15_wuser_f = desc_8_wuser_15_reg[31:0];
assign desc_8_data_host_addr_0_addr_f = desc_8_data_host_addr_0_reg[31:0];
assign desc_8_data_host_addr_1_addr_f = desc_8_data_host_addr_1_reg[31:0];
assign desc_8_data_host_addr_2_addr_f = desc_8_data_host_addr_2_reg[31:0];
assign desc_8_data_host_addr_3_addr_f = desc_8_data_host_addr_3_reg[31:0];
assign desc_8_wstrb_host_addr_0_addr_f = desc_8_wstrb_host_addr_0_reg[31:0];
assign desc_8_wstrb_host_addr_1_addr_f = desc_8_wstrb_host_addr_1_reg[31:0];
assign desc_8_wstrb_host_addr_2_addr_f = desc_8_wstrb_host_addr_2_reg[31:0];
assign desc_8_wstrb_host_addr_3_addr_f = desc_8_wstrb_host_addr_3_reg[31:0];
assign desc_8_xuser_0_xuser_f = desc_8_xuser_0_reg[31:0];
assign desc_8_xuser_1_xuser_f = desc_8_xuser_1_reg[31:0];
assign desc_8_xuser_2_xuser_f = desc_8_xuser_2_reg[31:0];
assign desc_8_xuser_3_xuser_f = desc_8_xuser_3_reg[31:0];
assign desc_8_xuser_4_xuser_f = desc_8_xuser_4_reg[31:0];
assign desc_8_xuser_5_xuser_f = desc_8_xuser_5_reg[31:0];
assign desc_8_xuser_6_xuser_f = desc_8_xuser_6_reg[31:0];
assign desc_8_xuser_7_xuser_f = desc_8_xuser_7_reg[31:0];
assign desc_8_xuser_8_xuser_f = desc_8_xuser_8_reg[31:0];
assign desc_8_xuser_9_xuser_f = desc_8_xuser_9_reg[31:0];
assign desc_8_xuser_10_xuser_f = desc_8_xuser_10_reg[31:0];
assign desc_8_xuser_11_xuser_f = desc_8_xuser_11_reg[31:0];
assign desc_8_xuser_12_xuser_f = desc_8_xuser_12_reg[31:0];
assign desc_8_xuser_13_xuser_f = desc_8_xuser_13_reg[31:0];
assign desc_8_xuser_14_xuser_f = desc_8_xuser_14_reg[31:0];
assign desc_8_xuser_15_xuser_f = desc_8_xuser_15_reg[31:0];
assign desc_9_txn_type_wr_strb_f = desc_9_txn_type_reg[1];
assign desc_9_txn_type_wr_rd_f = desc_9_txn_type_reg[0];
assign desc_9_attr_axregion_f = desc_9_attr_reg[18:15];
assign desc_9_attr_axqos_f = desc_9_attr_reg[14:11];
assign desc_9_attr_axprot_f = desc_9_attr_reg[10:8];
assign desc_9_attr_axcache_f = desc_9_attr_reg[7:4];
assign desc_9_attr_axlock_f = desc_9_attr_reg[3:2];
assign desc_9_attr_axburst_f = desc_9_attr_reg[1:0];
assign desc_9_axid_0_axid_f = desc_9_axid_0_reg[31:0];
assign desc_9_axid_1_axid_f = desc_9_axid_1_reg[31:0];
assign desc_9_axid_2_axid_f = desc_9_axid_2_reg[31:0];
assign desc_9_axid_3_axid_f = desc_9_axid_3_reg[31:0];
assign desc_9_axuser_0_axuser_f = desc_9_axuser_0_reg[31:0];
assign desc_9_axuser_1_axuser_f = desc_9_axuser_1_reg[31:0];
assign desc_9_axuser_2_axuser_f = desc_9_axuser_2_reg[31:0];
assign desc_9_axuser_3_axuser_f = desc_9_axuser_3_reg[31:0];
assign desc_9_axuser_4_axuser_f = desc_9_axuser_4_reg[31:0];
assign desc_9_axuser_5_axuser_f = desc_9_axuser_5_reg[31:0];
assign desc_9_axuser_6_axuser_f = desc_9_axuser_6_reg[31:0];
assign desc_9_axuser_7_axuser_f = desc_9_axuser_7_reg[31:0];
assign desc_9_axuser_8_axuser_f = desc_9_axuser_8_reg[31:0];
assign desc_9_axuser_9_axuser_f = desc_9_axuser_9_reg[31:0];
assign desc_9_axuser_10_axuser_f = desc_9_axuser_10_reg[31:0];
assign desc_9_axuser_11_axuser_f = desc_9_axuser_11_reg[31:0];
assign desc_9_axuser_12_axuser_f = desc_9_axuser_12_reg[31:0];
assign desc_9_axuser_13_axuser_f = desc_9_axuser_13_reg[31:0];
assign desc_9_axuser_14_axuser_f = desc_9_axuser_14_reg[31:0];
assign desc_9_axuser_15_axuser_f = desc_9_axuser_15_reg[31:0];
assign desc_9_size_txn_size_f = desc_9_size_reg[15:0];
assign desc_9_axsize_axsize_f = desc_9_axsize_reg[2:0];
assign desc_9_axaddr_0_addr_f = desc_9_axaddr_0_reg[31:0];
assign desc_9_axaddr_1_addr_f = desc_9_axaddr_1_reg[31:0];
assign desc_9_axaddr_2_addr_f = desc_9_axaddr_2_reg[31:0];
assign desc_9_axaddr_3_addr_f = desc_9_axaddr_3_reg[31:0];
assign desc_9_data_offset_addr_f = desc_9_data_offset_reg[31:0];
assign desc_9_wuser_0_wuser_f = desc_9_wuser_0_reg[31:0];
assign desc_9_wuser_1_wuser_f = desc_9_wuser_1_reg[31:0];
assign desc_9_wuser_2_wuser_f = desc_9_wuser_2_reg[31:0];
assign desc_9_wuser_3_wuser_f = desc_9_wuser_3_reg[31:0];
assign desc_9_wuser_4_wuser_f = desc_9_wuser_4_reg[31:0];
assign desc_9_wuser_5_wuser_f = desc_9_wuser_5_reg[31:0];
assign desc_9_wuser_6_wuser_f = desc_9_wuser_6_reg[31:0];
assign desc_9_wuser_7_wuser_f = desc_9_wuser_7_reg[31:0];
assign desc_9_wuser_8_wuser_f = desc_9_wuser_8_reg[31:0];
assign desc_9_wuser_9_wuser_f = desc_9_wuser_9_reg[31:0];
assign desc_9_wuser_10_wuser_f = desc_9_wuser_10_reg[31:0];
assign desc_9_wuser_11_wuser_f = desc_9_wuser_11_reg[31:0];
assign desc_9_wuser_12_wuser_f = desc_9_wuser_12_reg[31:0];
assign desc_9_wuser_13_wuser_f = desc_9_wuser_13_reg[31:0];
assign desc_9_wuser_14_wuser_f = desc_9_wuser_14_reg[31:0];
assign desc_9_wuser_15_wuser_f = desc_9_wuser_15_reg[31:0];
assign desc_9_data_host_addr_0_addr_f = desc_9_data_host_addr_0_reg[31:0];
assign desc_9_data_host_addr_1_addr_f = desc_9_data_host_addr_1_reg[31:0];
assign desc_9_data_host_addr_2_addr_f = desc_9_data_host_addr_2_reg[31:0];
assign desc_9_data_host_addr_3_addr_f = desc_9_data_host_addr_3_reg[31:0];
assign desc_9_wstrb_host_addr_0_addr_f = desc_9_wstrb_host_addr_0_reg[31:0];
assign desc_9_wstrb_host_addr_1_addr_f = desc_9_wstrb_host_addr_1_reg[31:0];
assign desc_9_wstrb_host_addr_2_addr_f = desc_9_wstrb_host_addr_2_reg[31:0];
assign desc_9_wstrb_host_addr_3_addr_f = desc_9_wstrb_host_addr_3_reg[31:0];
assign desc_9_xuser_0_xuser_f = desc_9_xuser_0_reg[31:0];
assign desc_9_xuser_1_xuser_f = desc_9_xuser_1_reg[31:0];
assign desc_9_xuser_2_xuser_f = desc_9_xuser_2_reg[31:0];
assign desc_9_xuser_3_xuser_f = desc_9_xuser_3_reg[31:0];
assign desc_9_xuser_4_xuser_f = desc_9_xuser_4_reg[31:0];
assign desc_9_xuser_5_xuser_f = desc_9_xuser_5_reg[31:0];
assign desc_9_xuser_6_xuser_f = desc_9_xuser_6_reg[31:0];
assign desc_9_xuser_7_xuser_f = desc_9_xuser_7_reg[31:0];
assign desc_9_xuser_8_xuser_f = desc_9_xuser_8_reg[31:0];
assign desc_9_xuser_9_xuser_f = desc_9_xuser_9_reg[31:0];
assign desc_9_xuser_10_xuser_f = desc_9_xuser_10_reg[31:0];
assign desc_9_xuser_11_xuser_f = desc_9_xuser_11_reg[31:0];
assign desc_9_xuser_12_xuser_f = desc_9_xuser_12_reg[31:0];
assign desc_9_xuser_13_xuser_f = desc_9_xuser_13_reg[31:0];
assign desc_9_xuser_14_xuser_f = desc_9_xuser_14_reg[31:0];
assign desc_9_xuser_15_xuser_f = desc_9_xuser_15_reg[31:0];
assign desc_10_txn_type_wr_strb_f = desc_10_txn_type_reg[1];
assign desc_10_txn_type_wr_rd_f = desc_10_txn_type_reg[0];
assign desc_10_attr_axregion_f = desc_10_attr_reg[18:15];
assign desc_10_attr_axqos_f = desc_10_attr_reg[14:11];
assign desc_10_attr_axprot_f = desc_10_attr_reg[10:8];
assign desc_10_attr_axcache_f = desc_10_attr_reg[7:4];
assign desc_10_attr_axlock_f = desc_10_attr_reg[3:2];
assign desc_10_attr_axburst_f = desc_10_attr_reg[1:0];
assign desc_10_axid_0_axid_f = desc_10_axid_0_reg[31:0];
assign desc_10_axid_1_axid_f = desc_10_axid_1_reg[31:0];
assign desc_10_axid_2_axid_f = desc_10_axid_2_reg[31:0];
assign desc_10_axid_3_axid_f = desc_10_axid_3_reg[31:0];
assign desc_10_axuser_0_axuser_f = desc_10_axuser_0_reg[31:0];
assign desc_10_axuser_1_axuser_f = desc_10_axuser_1_reg[31:0];
assign desc_10_axuser_2_axuser_f = desc_10_axuser_2_reg[31:0];
assign desc_10_axuser_3_axuser_f = desc_10_axuser_3_reg[31:0];
assign desc_10_axuser_4_axuser_f = desc_10_axuser_4_reg[31:0];
assign desc_10_axuser_5_axuser_f = desc_10_axuser_5_reg[31:0];
assign desc_10_axuser_6_axuser_f = desc_10_axuser_6_reg[31:0];
assign desc_10_axuser_7_axuser_f = desc_10_axuser_7_reg[31:0];
assign desc_10_axuser_8_axuser_f = desc_10_axuser_8_reg[31:0];
assign desc_10_axuser_9_axuser_f = desc_10_axuser_9_reg[31:0];
assign desc_10_axuser_10_axuser_f = desc_10_axuser_10_reg[31:0];
assign desc_10_axuser_11_axuser_f = desc_10_axuser_11_reg[31:0];
assign desc_10_axuser_12_axuser_f = desc_10_axuser_12_reg[31:0];
assign desc_10_axuser_13_axuser_f = desc_10_axuser_13_reg[31:0];
assign desc_10_axuser_14_axuser_f = desc_10_axuser_14_reg[31:0];
assign desc_10_axuser_15_axuser_f = desc_10_axuser_15_reg[31:0];
assign desc_10_size_txn_size_f = desc_10_size_reg[15:0];
assign desc_10_axsize_axsize_f = desc_10_axsize_reg[2:0];
assign desc_10_axaddr_0_addr_f = desc_10_axaddr_0_reg[31:0];
assign desc_10_axaddr_1_addr_f = desc_10_axaddr_1_reg[31:0];
assign desc_10_axaddr_2_addr_f = desc_10_axaddr_2_reg[31:0];
assign desc_10_axaddr_3_addr_f = desc_10_axaddr_3_reg[31:0];
assign desc_10_data_offset_addr_f = desc_10_data_offset_reg[31:0];
assign desc_10_wuser_0_wuser_f = desc_10_wuser_0_reg[31:0];
assign desc_10_wuser_1_wuser_f = desc_10_wuser_1_reg[31:0];
assign desc_10_wuser_2_wuser_f = desc_10_wuser_2_reg[31:0];
assign desc_10_wuser_3_wuser_f = desc_10_wuser_3_reg[31:0];
assign desc_10_wuser_4_wuser_f = desc_10_wuser_4_reg[31:0];
assign desc_10_wuser_5_wuser_f = desc_10_wuser_5_reg[31:0];
assign desc_10_wuser_6_wuser_f = desc_10_wuser_6_reg[31:0];
assign desc_10_wuser_7_wuser_f = desc_10_wuser_7_reg[31:0];
assign desc_10_wuser_8_wuser_f = desc_10_wuser_8_reg[31:0];
assign desc_10_wuser_9_wuser_f = desc_10_wuser_9_reg[31:0];
assign desc_10_wuser_10_wuser_f = desc_10_wuser_10_reg[31:0];
assign desc_10_wuser_11_wuser_f = desc_10_wuser_11_reg[31:0];
assign desc_10_wuser_12_wuser_f = desc_10_wuser_12_reg[31:0];
assign desc_10_wuser_13_wuser_f = desc_10_wuser_13_reg[31:0];
assign desc_10_wuser_14_wuser_f = desc_10_wuser_14_reg[31:0];
assign desc_10_wuser_15_wuser_f = desc_10_wuser_15_reg[31:0];
assign desc_10_data_host_addr_0_addr_f = desc_10_data_host_addr_0_reg[31:0];
assign desc_10_data_host_addr_1_addr_f = desc_10_data_host_addr_1_reg[31:0];
assign desc_10_data_host_addr_2_addr_f = desc_10_data_host_addr_2_reg[31:0];
assign desc_10_data_host_addr_3_addr_f = desc_10_data_host_addr_3_reg[31:0];
assign desc_10_wstrb_host_addr_0_addr_f = desc_10_wstrb_host_addr_0_reg[31:0];
assign desc_10_wstrb_host_addr_1_addr_f = desc_10_wstrb_host_addr_1_reg[31:0];
assign desc_10_wstrb_host_addr_2_addr_f = desc_10_wstrb_host_addr_2_reg[31:0];
assign desc_10_wstrb_host_addr_3_addr_f = desc_10_wstrb_host_addr_3_reg[31:0];
assign desc_10_xuser_0_xuser_f = desc_10_xuser_0_reg[31:0];
assign desc_10_xuser_1_xuser_f = desc_10_xuser_1_reg[31:0];
assign desc_10_xuser_2_xuser_f = desc_10_xuser_2_reg[31:0];
assign desc_10_xuser_3_xuser_f = desc_10_xuser_3_reg[31:0];
assign desc_10_xuser_4_xuser_f = desc_10_xuser_4_reg[31:0];
assign desc_10_xuser_5_xuser_f = desc_10_xuser_5_reg[31:0];
assign desc_10_xuser_6_xuser_f = desc_10_xuser_6_reg[31:0];
assign desc_10_xuser_7_xuser_f = desc_10_xuser_7_reg[31:0];
assign desc_10_xuser_8_xuser_f = desc_10_xuser_8_reg[31:0];
assign desc_10_xuser_9_xuser_f = desc_10_xuser_9_reg[31:0];
assign desc_10_xuser_10_xuser_f = desc_10_xuser_10_reg[31:0];
assign desc_10_xuser_11_xuser_f = desc_10_xuser_11_reg[31:0];
assign desc_10_xuser_12_xuser_f = desc_10_xuser_12_reg[31:0];
assign desc_10_xuser_13_xuser_f = desc_10_xuser_13_reg[31:0];
assign desc_10_xuser_14_xuser_f = desc_10_xuser_14_reg[31:0];
assign desc_10_xuser_15_xuser_f = desc_10_xuser_15_reg[31:0];
assign desc_11_txn_type_wr_strb_f = desc_11_txn_type_reg[1];
assign desc_11_txn_type_wr_rd_f = desc_11_txn_type_reg[0];
assign desc_11_attr_axregion_f = desc_11_attr_reg[18:15];
assign desc_11_attr_axqos_f = desc_11_attr_reg[14:11];
assign desc_11_attr_axprot_f = desc_11_attr_reg[10:8];
assign desc_11_attr_axcache_f = desc_11_attr_reg[7:4];
assign desc_11_attr_axlock_f = desc_11_attr_reg[3:2];
assign desc_11_attr_axburst_f = desc_11_attr_reg[1:0];
assign desc_11_axid_0_axid_f = desc_11_axid_0_reg[31:0];
assign desc_11_axid_1_axid_f = desc_11_axid_1_reg[31:0];
assign desc_11_axid_2_axid_f = desc_11_axid_2_reg[31:0];
assign desc_11_axid_3_axid_f = desc_11_axid_3_reg[31:0];
assign desc_11_axuser_0_axuser_f = desc_11_axuser_0_reg[31:0];
assign desc_11_axuser_1_axuser_f = desc_11_axuser_1_reg[31:0];
assign desc_11_axuser_2_axuser_f = desc_11_axuser_2_reg[31:0];
assign desc_11_axuser_3_axuser_f = desc_11_axuser_3_reg[31:0];
assign desc_11_axuser_4_axuser_f = desc_11_axuser_4_reg[31:0];
assign desc_11_axuser_5_axuser_f = desc_11_axuser_5_reg[31:0];
assign desc_11_axuser_6_axuser_f = desc_11_axuser_6_reg[31:0];
assign desc_11_axuser_7_axuser_f = desc_11_axuser_7_reg[31:0];
assign desc_11_axuser_8_axuser_f = desc_11_axuser_8_reg[31:0];
assign desc_11_axuser_9_axuser_f = desc_11_axuser_9_reg[31:0];
assign desc_11_axuser_10_axuser_f = desc_11_axuser_10_reg[31:0];
assign desc_11_axuser_11_axuser_f = desc_11_axuser_11_reg[31:0];
assign desc_11_axuser_12_axuser_f = desc_11_axuser_12_reg[31:0];
assign desc_11_axuser_13_axuser_f = desc_11_axuser_13_reg[31:0];
assign desc_11_axuser_14_axuser_f = desc_11_axuser_14_reg[31:0];
assign desc_11_axuser_15_axuser_f = desc_11_axuser_15_reg[31:0];
assign desc_11_size_txn_size_f = desc_11_size_reg[15:0];
assign desc_11_axsize_axsize_f = desc_11_axsize_reg[2:0];
assign desc_11_axaddr_0_addr_f = desc_11_axaddr_0_reg[31:0];
assign desc_11_axaddr_1_addr_f = desc_11_axaddr_1_reg[31:0];
assign desc_11_axaddr_2_addr_f = desc_11_axaddr_2_reg[31:0];
assign desc_11_axaddr_3_addr_f = desc_11_axaddr_3_reg[31:0];
assign desc_11_data_offset_addr_f = desc_11_data_offset_reg[31:0];
assign desc_11_wuser_0_wuser_f = desc_11_wuser_0_reg[31:0];
assign desc_11_wuser_1_wuser_f = desc_11_wuser_1_reg[31:0];
assign desc_11_wuser_2_wuser_f = desc_11_wuser_2_reg[31:0];
assign desc_11_wuser_3_wuser_f = desc_11_wuser_3_reg[31:0];
assign desc_11_wuser_4_wuser_f = desc_11_wuser_4_reg[31:0];
assign desc_11_wuser_5_wuser_f = desc_11_wuser_5_reg[31:0];
assign desc_11_wuser_6_wuser_f = desc_11_wuser_6_reg[31:0];
assign desc_11_wuser_7_wuser_f = desc_11_wuser_7_reg[31:0];
assign desc_11_wuser_8_wuser_f = desc_11_wuser_8_reg[31:0];
assign desc_11_wuser_9_wuser_f = desc_11_wuser_9_reg[31:0];
assign desc_11_wuser_10_wuser_f = desc_11_wuser_10_reg[31:0];
assign desc_11_wuser_11_wuser_f = desc_11_wuser_11_reg[31:0];
assign desc_11_wuser_12_wuser_f = desc_11_wuser_12_reg[31:0];
assign desc_11_wuser_13_wuser_f = desc_11_wuser_13_reg[31:0];
assign desc_11_wuser_14_wuser_f = desc_11_wuser_14_reg[31:0];
assign desc_11_wuser_15_wuser_f = desc_11_wuser_15_reg[31:0];
assign desc_11_data_host_addr_0_addr_f = desc_11_data_host_addr_0_reg[31:0];
assign desc_11_data_host_addr_1_addr_f = desc_11_data_host_addr_1_reg[31:0];
assign desc_11_data_host_addr_2_addr_f = desc_11_data_host_addr_2_reg[31:0];
assign desc_11_data_host_addr_3_addr_f = desc_11_data_host_addr_3_reg[31:0];
assign desc_11_wstrb_host_addr_0_addr_f = desc_11_wstrb_host_addr_0_reg[31:0];
assign desc_11_wstrb_host_addr_1_addr_f = desc_11_wstrb_host_addr_1_reg[31:0];
assign desc_11_wstrb_host_addr_2_addr_f = desc_11_wstrb_host_addr_2_reg[31:0];
assign desc_11_wstrb_host_addr_3_addr_f = desc_11_wstrb_host_addr_3_reg[31:0];
assign desc_11_xuser_0_xuser_f = desc_11_xuser_0_reg[31:0];
assign desc_11_xuser_1_xuser_f = desc_11_xuser_1_reg[31:0];
assign desc_11_xuser_2_xuser_f = desc_11_xuser_2_reg[31:0];
assign desc_11_xuser_3_xuser_f = desc_11_xuser_3_reg[31:0];
assign desc_11_xuser_4_xuser_f = desc_11_xuser_4_reg[31:0];
assign desc_11_xuser_5_xuser_f = desc_11_xuser_5_reg[31:0];
assign desc_11_xuser_6_xuser_f = desc_11_xuser_6_reg[31:0];
assign desc_11_xuser_7_xuser_f = desc_11_xuser_7_reg[31:0];
assign desc_11_xuser_8_xuser_f = desc_11_xuser_8_reg[31:0];
assign desc_11_xuser_9_xuser_f = desc_11_xuser_9_reg[31:0];
assign desc_11_xuser_10_xuser_f = desc_11_xuser_10_reg[31:0];
assign desc_11_xuser_11_xuser_f = desc_11_xuser_11_reg[31:0];
assign desc_11_xuser_12_xuser_f = desc_11_xuser_12_reg[31:0];
assign desc_11_xuser_13_xuser_f = desc_11_xuser_13_reg[31:0];
assign desc_11_xuser_14_xuser_f = desc_11_xuser_14_reg[31:0];
assign desc_11_xuser_15_xuser_f = desc_11_xuser_15_reg[31:0];
assign desc_12_txn_type_wr_strb_f = desc_12_txn_type_reg[1];
assign desc_12_txn_type_wr_rd_f = desc_12_txn_type_reg[0];
assign desc_12_attr_axregion_f = desc_12_attr_reg[18:15];
assign desc_12_attr_axqos_f = desc_12_attr_reg[14:11];
assign desc_12_attr_axprot_f = desc_12_attr_reg[10:8];
assign desc_12_attr_axcache_f = desc_12_attr_reg[7:4];
assign desc_12_attr_axlock_f = desc_12_attr_reg[3:2];
assign desc_12_attr_axburst_f = desc_12_attr_reg[1:0];
assign desc_12_axid_0_axid_f = desc_12_axid_0_reg[31:0];
assign desc_12_axid_1_axid_f = desc_12_axid_1_reg[31:0];
assign desc_12_axid_2_axid_f = desc_12_axid_2_reg[31:0];
assign desc_12_axid_3_axid_f = desc_12_axid_3_reg[31:0];
assign desc_12_axuser_0_axuser_f = desc_12_axuser_0_reg[31:0];
assign desc_12_axuser_1_axuser_f = desc_12_axuser_1_reg[31:0];
assign desc_12_axuser_2_axuser_f = desc_12_axuser_2_reg[31:0];
assign desc_12_axuser_3_axuser_f = desc_12_axuser_3_reg[31:0];
assign desc_12_axuser_4_axuser_f = desc_12_axuser_4_reg[31:0];
assign desc_12_axuser_5_axuser_f = desc_12_axuser_5_reg[31:0];
assign desc_12_axuser_6_axuser_f = desc_12_axuser_6_reg[31:0];
assign desc_12_axuser_7_axuser_f = desc_12_axuser_7_reg[31:0];
assign desc_12_axuser_8_axuser_f = desc_12_axuser_8_reg[31:0];
assign desc_12_axuser_9_axuser_f = desc_12_axuser_9_reg[31:0];
assign desc_12_axuser_10_axuser_f = desc_12_axuser_10_reg[31:0];
assign desc_12_axuser_11_axuser_f = desc_12_axuser_11_reg[31:0];
assign desc_12_axuser_12_axuser_f = desc_12_axuser_12_reg[31:0];
assign desc_12_axuser_13_axuser_f = desc_12_axuser_13_reg[31:0];
assign desc_12_axuser_14_axuser_f = desc_12_axuser_14_reg[31:0];
assign desc_12_axuser_15_axuser_f = desc_12_axuser_15_reg[31:0];
assign desc_12_size_txn_size_f = desc_12_size_reg[15:0];
assign desc_12_axsize_axsize_f = desc_12_axsize_reg[2:0];
assign desc_12_axaddr_0_addr_f = desc_12_axaddr_0_reg[31:0];
assign desc_12_axaddr_1_addr_f = desc_12_axaddr_1_reg[31:0];
assign desc_12_axaddr_2_addr_f = desc_12_axaddr_2_reg[31:0];
assign desc_12_axaddr_3_addr_f = desc_12_axaddr_3_reg[31:0];
assign desc_12_data_offset_addr_f = desc_12_data_offset_reg[31:0];
assign desc_12_wuser_0_wuser_f = desc_12_wuser_0_reg[31:0];
assign desc_12_wuser_1_wuser_f = desc_12_wuser_1_reg[31:0];
assign desc_12_wuser_2_wuser_f = desc_12_wuser_2_reg[31:0];
assign desc_12_wuser_3_wuser_f = desc_12_wuser_3_reg[31:0];
assign desc_12_wuser_4_wuser_f = desc_12_wuser_4_reg[31:0];
assign desc_12_wuser_5_wuser_f = desc_12_wuser_5_reg[31:0];
assign desc_12_wuser_6_wuser_f = desc_12_wuser_6_reg[31:0];
assign desc_12_wuser_7_wuser_f = desc_12_wuser_7_reg[31:0];
assign desc_12_wuser_8_wuser_f = desc_12_wuser_8_reg[31:0];
assign desc_12_wuser_9_wuser_f = desc_12_wuser_9_reg[31:0];
assign desc_12_wuser_10_wuser_f = desc_12_wuser_10_reg[31:0];
assign desc_12_wuser_11_wuser_f = desc_12_wuser_11_reg[31:0];
assign desc_12_wuser_12_wuser_f = desc_12_wuser_12_reg[31:0];
assign desc_12_wuser_13_wuser_f = desc_12_wuser_13_reg[31:0];
assign desc_12_wuser_14_wuser_f = desc_12_wuser_14_reg[31:0];
assign desc_12_wuser_15_wuser_f = desc_12_wuser_15_reg[31:0];
assign desc_12_data_host_addr_0_addr_f = desc_12_data_host_addr_0_reg[31:0];
assign desc_12_data_host_addr_1_addr_f = desc_12_data_host_addr_1_reg[31:0];
assign desc_12_data_host_addr_2_addr_f = desc_12_data_host_addr_2_reg[31:0];
assign desc_12_data_host_addr_3_addr_f = desc_12_data_host_addr_3_reg[31:0];
assign desc_12_wstrb_host_addr_0_addr_f = desc_12_wstrb_host_addr_0_reg[31:0];
assign desc_12_wstrb_host_addr_1_addr_f = desc_12_wstrb_host_addr_1_reg[31:0];
assign desc_12_wstrb_host_addr_2_addr_f = desc_12_wstrb_host_addr_2_reg[31:0];
assign desc_12_wstrb_host_addr_3_addr_f = desc_12_wstrb_host_addr_3_reg[31:0];
assign desc_12_xuser_0_xuser_f = desc_12_xuser_0_reg[31:0];
assign desc_12_xuser_1_xuser_f = desc_12_xuser_1_reg[31:0];
assign desc_12_xuser_2_xuser_f = desc_12_xuser_2_reg[31:0];
assign desc_12_xuser_3_xuser_f = desc_12_xuser_3_reg[31:0];
assign desc_12_xuser_4_xuser_f = desc_12_xuser_4_reg[31:0];
assign desc_12_xuser_5_xuser_f = desc_12_xuser_5_reg[31:0];
assign desc_12_xuser_6_xuser_f = desc_12_xuser_6_reg[31:0];
assign desc_12_xuser_7_xuser_f = desc_12_xuser_7_reg[31:0];
assign desc_12_xuser_8_xuser_f = desc_12_xuser_8_reg[31:0];
assign desc_12_xuser_9_xuser_f = desc_12_xuser_9_reg[31:0];
assign desc_12_xuser_10_xuser_f = desc_12_xuser_10_reg[31:0];
assign desc_12_xuser_11_xuser_f = desc_12_xuser_11_reg[31:0];
assign desc_12_xuser_12_xuser_f = desc_12_xuser_12_reg[31:0];
assign desc_12_xuser_13_xuser_f = desc_12_xuser_13_reg[31:0];
assign desc_12_xuser_14_xuser_f = desc_12_xuser_14_reg[31:0];
assign desc_12_xuser_15_xuser_f = desc_12_xuser_15_reg[31:0];
assign desc_13_txn_type_wr_strb_f = desc_13_txn_type_reg[1];
assign desc_13_txn_type_wr_rd_f = desc_13_txn_type_reg[0];
assign desc_13_attr_axregion_f = desc_13_attr_reg[18:15];
assign desc_13_attr_axqos_f = desc_13_attr_reg[14:11];
assign desc_13_attr_axprot_f = desc_13_attr_reg[10:8];
assign desc_13_attr_axcache_f = desc_13_attr_reg[7:4];
assign desc_13_attr_axlock_f = desc_13_attr_reg[3:2];
assign desc_13_attr_axburst_f = desc_13_attr_reg[1:0];
assign desc_13_axid_0_axid_f = desc_13_axid_0_reg[31:0];
assign desc_13_axid_1_axid_f = desc_13_axid_1_reg[31:0];
assign desc_13_axid_2_axid_f = desc_13_axid_2_reg[31:0];
assign desc_13_axid_3_axid_f = desc_13_axid_3_reg[31:0];
assign desc_13_axuser_0_axuser_f = desc_13_axuser_0_reg[31:0];
assign desc_13_axuser_1_axuser_f = desc_13_axuser_1_reg[31:0];
assign desc_13_axuser_2_axuser_f = desc_13_axuser_2_reg[31:0];
assign desc_13_axuser_3_axuser_f = desc_13_axuser_3_reg[31:0];
assign desc_13_axuser_4_axuser_f = desc_13_axuser_4_reg[31:0];
assign desc_13_axuser_5_axuser_f = desc_13_axuser_5_reg[31:0];
assign desc_13_axuser_6_axuser_f = desc_13_axuser_6_reg[31:0];
assign desc_13_axuser_7_axuser_f = desc_13_axuser_7_reg[31:0];
assign desc_13_axuser_8_axuser_f = desc_13_axuser_8_reg[31:0];
assign desc_13_axuser_9_axuser_f = desc_13_axuser_9_reg[31:0];
assign desc_13_axuser_10_axuser_f = desc_13_axuser_10_reg[31:0];
assign desc_13_axuser_11_axuser_f = desc_13_axuser_11_reg[31:0];
assign desc_13_axuser_12_axuser_f = desc_13_axuser_12_reg[31:0];
assign desc_13_axuser_13_axuser_f = desc_13_axuser_13_reg[31:0];
assign desc_13_axuser_14_axuser_f = desc_13_axuser_14_reg[31:0];
assign desc_13_axuser_15_axuser_f = desc_13_axuser_15_reg[31:0];
assign desc_13_size_txn_size_f = desc_13_size_reg[15:0];
assign desc_13_axsize_axsize_f = desc_13_axsize_reg[2:0];
assign desc_13_axaddr_0_addr_f = desc_13_axaddr_0_reg[31:0];
assign desc_13_axaddr_1_addr_f = desc_13_axaddr_1_reg[31:0];
assign desc_13_axaddr_2_addr_f = desc_13_axaddr_2_reg[31:0];
assign desc_13_axaddr_3_addr_f = desc_13_axaddr_3_reg[31:0];
assign desc_13_data_offset_addr_f = desc_13_data_offset_reg[31:0];
assign desc_13_wuser_0_wuser_f = desc_13_wuser_0_reg[31:0];
assign desc_13_wuser_1_wuser_f = desc_13_wuser_1_reg[31:0];
assign desc_13_wuser_2_wuser_f = desc_13_wuser_2_reg[31:0];
assign desc_13_wuser_3_wuser_f = desc_13_wuser_3_reg[31:0];
assign desc_13_wuser_4_wuser_f = desc_13_wuser_4_reg[31:0];
assign desc_13_wuser_5_wuser_f = desc_13_wuser_5_reg[31:0];
assign desc_13_wuser_6_wuser_f = desc_13_wuser_6_reg[31:0];
assign desc_13_wuser_7_wuser_f = desc_13_wuser_7_reg[31:0];
assign desc_13_wuser_8_wuser_f = desc_13_wuser_8_reg[31:0];
assign desc_13_wuser_9_wuser_f = desc_13_wuser_9_reg[31:0];
assign desc_13_wuser_10_wuser_f = desc_13_wuser_10_reg[31:0];
assign desc_13_wuser_11_wuser_f = desc_13_wuser_11_reg[31:0];
assign desc_13_wuser_12_wuser_f = desc_13_wuser_12_reg[31:0];
assign desc_13_wuser_13_wuser_f = desc_13_wuser_13_reg[31:0];
assign desc_13_wuser_14_wuser_f = desc_13_wuser_14_reg[31:0];
assign desc_13_wuser_15_wuser_f = desc_13_wuser_15_reg[31:0];
assign desc_13_data_host_addr_0_addr_f = desc_13_data_host_addr_0_reg[31:0];
assign desc_13_data_host_addr_1_addr_f = desc_13_data_host_addr_1_reg[31:0];
assign desc_13_data_host_addr_2_addr_f = desc_13_data_host_addr_2_reg[31:0];
assign desc_13_data_host_addr_3_addr_f = desc_13_data_host_addr_3_reg[31:0];
assign desc_13_wstrb_host_addr_0_addr_f = desc_13_wstrb_host_addr_0_reg[31:0];
assign desc_13_wstrb_host_addr_1_addr_f = desc_13_wstrb_host_addr_1_reg[31:0];
assign desc_13_wstrb_host_addr_2_addr_f = desc_13_wstrb_host_addr_2_reg[31:0];
assign desc_13_wstrb_host_addr_3_addr_f = desc_13_wstrb_host_addr_3_reg[31:0];
assign desc_13_xuser_0_xuser_f = desc_13_xuser_0_reg[31:0];
assign desc_13_xuser_1_xuser_f = desc_13_xuser_1_reg[31:0];
assign desc_13_xuser_2_xuser_f = desc_13_xuser_2_reg[31:0];
assign desc_13_xuser_3_xuser_f = desc_13_xuser_3_reg[31:0];
assign desc_13_xuser_4_xuser_f = desc_13_xuser_4_reg[31:0];
assign desc_13_xuser_5_xuser_f = desc_13_xuser_5_reg[31:0];
assign desc_13_xuser_6_xuser_f = desc_13_xuser_6_reg[31:0];
assign desc_13_xuser_7_xuser_f = desc_13_xuser_7_reg[31:0];
assign desc_13_xuser_8_xuser_f = desc_13_xuser_8_reg[31:0];
assign desc_13_xuser_9_xuser_f = desc_13_xuser_9_reg[31:0];
assign desc_13_xuser_10_xuser_f = desc_13_xuser_10_reg[31:0];
assign desc_13_xuser_11_xuser_f = desc_13_xuser_11_reg[31:0];
assign desc_13_xuser_12_xuser_f = desc_13_xuser_12_reg[31:0];
assign desc_13_xuser_13_xuser_f = desc_13_xuser_13_reg[31:0];
assign desc_13_xuser_14_xuser_f = desc_13_xuser_14_reg[31:0];
assign desc_13_xuser_15_xuser_f = desc_13_xuser_15_reg[31:0];
assign desc_14_txn_type_wr_strb_f = desc_14_txn_type_reg[1];
assign desc_14_txn_type_wr_rd_f = desc_14_txn_type_reg[0];
assign desc_14_attr_axregion_f = desc_14_attr_reg[18:15];
assign desc_14_attr_axqos_f = desc_14_attr_reg[14:11];
assign desc_14_attr_axprot_f = desc_14_attr_reg[10:8];
assign desc_14_attr_axcache_f = desc_14_attr_reg[7:4];
assign desc_14_attr_axlock_f = desc_14_attr_reg[3:2];
assign desc_14_attr_axburst_f = desc_14_attr_reg[1:0];
assign desc_14_axid_0_axid_f = desc_14_axid_0_reg[31:0];
assign desc_14_axid_1_axid_f = desc_14_axid_1_reg[31:0];
assign desc_14_axid_2_axid_f = desc_14_axid_2_reg[31:0];
assign desc_14_axid_3_axid_f = desc_14_axid_3_reg[31:0];
assign desc_14_axuser_0_axuser_f = desc_14_axuser_0_reg[31:0];
assign desc_14_axuser_1_axuser_f = desc_14_axuser_1_reg[31:0];
assign desc_14_axuser_2_axuser_f = desc_14_axuser_2_reg[31:0];
assign desc_14_axuser_3_axuser_f = desc_14_axuser_3_reg[31:0];
assign desc_14_axuser_4_axuser_f = desc_14_axuser_4_reg[31:0];
assign desc_14_axuser_5_axuser_f = desc_14_axuser_5_reg[31:0];
assign desc_14_axuser_6_axuser_f = desc_14_axuser_6_reg[31:0];
assign desc_14_axuser_7_axuser_f = desc_14_axuser_7_reg[31:0];
assign desc_14_axuser_8_axuser_f = desc_14_axuser_8_reg[31:0];
assign desc_14_axuser_9_axuser_f = desc_14_axuser_9_reg[31:0];
assign desc_14_axuser_10_axuser_f = desc_14_axuser_10_reg[31:0];
assign desc_14_axuser_11_axuser_f = desc_14_axuser_11_reg[31:0];
assign desc_14_axuser_12_axuser_f = desc_14_axuser_12_reg[31:0];
assign desc_14_axuser_13_axuser_f = desc_14_axuser_13_reg[31:0];
assign desc_14_axuser_14_axuser_f = desc_14_axuser_14_reg[31:0];
assign desc_14_axuser_15_axuser_f = desc_14_axuser_15_reg[31:0];
assign desc_14_size_txn_size_f = desc_14_size_reg[15:0];
assign desc_14_axsize_axsize_f = desc_14_axsize_reg[2:0];
assign desc_14_axaddr_0_addr_f = desc_14_axaddr_0_reg[31:0];
assign desc_14_axaddr_1_addr_f = desc_14_axaddr_1_reg[31:0];
assign desc_14_axaddr_2_addr_f = desc_14_axaddr_2_reg[31:0];
assign desc_14_axaddr_3_addr_f = desc_14_axaddr_3_reg[31:0];
assign desc_14_data_offset_addr_f = desc_14_data_offset_reg[31:0];
assign desc_14_wuser_0_wuser_f = desc_14_wuser_0_reg[31:0];
assign desc_14_wuser_1_wuser_f = desc_14_wuser_1_reg[31:0];
assign desc_14_wuser_2_wuser_f = desc_14_wuser_2_reg[31:0];
assign desc_14_wuser_3_wuser_f = desc_14_wuser_3_reg[31:0];
assign desc_14_wuser_4_wuser_f = desc_14_wuser_4_reg[31:0];
assign desc_14_wuser_5_wuser_f = desc_14_wuser_5_reg[31:0];
assign desc_14_wuser_6_wuser_f = desc_14_wuser_6_reg[31:0];
assign desc_14_wuser_7_wuser_f = desc_14_wuser_7_reg[31:0];
assign desc_14_wuser_8_wuser_f = desc_14_wuser_8_reg[31:0];
assign desc_14_wuser_9_wuser_f = desc_14_wuser_9_reg[31:0];
assign desc_14_wuser_10_wuser_f = desc_14_wuser_10_reg[31:0];
assign desc_14_wuser_11_wuser_f = desc_14_wuser_11_reg[31:0];
assign desc_14_wuser_12_wuser_f = desc_14_wuser_12_reg[31:0];
assign desc_14_wuser_13_wuser_f = desc_14_wuser_13_reg[31:0];
assign desc_14_wuser_14_wuser_f = desc_14_wuser_14_reg[31:0];
assign desc_14_wuser_15_wuser_f = desc_14_wuser_15_reg[31:0];
assign desc_14_data_host_addr_0_addr_f = desc_14_data_host_addr_0_reg[31:0];
assign desc_14_data_host_addr_1_addr_f = desc_14_data_host_addr_1_reg[31:0];
assign desc_14_data_host_addr_2_addr_f = desc_14_data_host_addr_2_reg[31:0];
assign desc_14_data_host_addr_3_addr_f = desc_14_data_host_addr_3_reg[31:0];
assign desc_14_wstrb_host_addr_0_addr_f = desc_14_wstrb_host_addr_0_reg[31:0];
assign desc_14_wstrb_host_addr_1_addr_f = desc_14_wstrb_host_addr_1_reg[31:0];
assign desc_14_wstrb_host_addr_2_addr_f = desc_14_wstrb_host_addr_2_reg[31:0];
assign desc_14_wstrb_host_addr_3_addr_f = desc_14_wstrb_host_addr_3_reg[31:0];
assign desc_14_xuser_0_xuser_f = desc_14_xuser_0_reg[31:0];
assign desc_14_xuser_1_xuser_f = desc_14_xuser_1_reg[31:0];
assign desc_14_xuser_2_xuser_f = desc_14_xuser_2_reg[31:0];
assign desc_14_xuser_3_xuser_f = desc_14_xuser_3_reg[31:0];
assign desc_14_xuser_4_xuser_f = desc_14_xuser_4_reg[31:0];
assign desc_14_xuser_5_xuser_f = desc_14_xuser_5_reg[31:0];
assign desc_14_xuser_6_xuser_f = desc_14_xuser_6_reg[31:0];
assign desc_14_xuser_7_xuser_f = desc_14_xuser_7_reg[31:0];
assign desc_14_xuser_8_xuser_f = desc_14_xuser_8_reg[31:0];
assign desc_14_xuser_9_xuser_f = desc_14_xuser_9_reg[31:0];
assign desc_14_xuser_10_xuser_f = desc_14_xuser_10_reg[31:0];
assign desc_14_xuser_11_xuser_f = desc_14_xuser_11_reg[31:0];
assign desc_14_xuser_12_xuser_f = desc_14_xuser_12_reg[31:0];
assign desc_14_xuser_13_xuser_f = desc_14_xuser_13_reg[31:0];
assign desc_14_xuser_14_xuser_f = desc_14_xuser_14_reg[31:0];
assign desc_14_xuser_15_xuser_f = desc_14_xuser_15_reg[31:0];
assign desc_15_txn_type_wr_strb_f = desc_15_txn_type_reg[1];
assign desc_15_txn_type_wr_rd_f = desc_15_txn_type_reg[0];
assign desc_15_attr_axregion_f = desc_15_attr_reg[18:15];
assign desc_15_attr_axqos_f = desc_15_attr_reg[14:11];
assign desc_15_attr_axprot_f = desc_15_attr_reg[10:8];
assign desc_15_attr_axcache_f = desc_15_attr_reg[7:4];
assign desc_15_attr_axlock_f = desc_15_attr_reg[3:2];
assign desc_15_attr_axburst_f = desc_15_attr_reg[1:0];
assign desc_15_axid_0_axid_f = desc_15_axid_0_reg[31:0];
assign desc_15_axid_1_axid_f = desc_15_axid_1_reg[31:0];
assign desc_15_axid_2_axid_f = desc_15_axid_2_reg[31:0];
assign desc_15_axid_3_axid_f = desc_15_axid_3_reg[31:0];
assign desc_15_axuser_0_axuser_f = desc_15_axuser_0_reg[31:0];
assign desc_15_axuser_1_axuser_f = desc_15_axuser_1_reg[31:0];
assign desc_15_axuser_2_axuser_f = desc_15_axuser_2_reg[31:0];
assign desc_15_axuser_3_axuser_f = desc_15_axuser_3_reg[31:0];
assign desc_15_axuser_4_axuser_f = desc_15_axuser_4_reg[31:0];
assign desc_15_axuser_5_axuser_f = desc_15_axuser_5_reg[31:0];
assign desc_15_axuser_6_axuser_f = desc_15_axuser_6_reg[31:0];
assign desc_15_axuser_7_axuser_f = desc_15_axuser_7_reg[31:0];
assign desc_15_axuser_8_axuser_f = desc_15_axuser_8_reg[31:0];
assign desc_15_axuser_9_axuser_f = desc_15_axuser_9_reg[31:0];
assign desc_15_axuser_10_axuser_f = desc_15_axuser_10_reg[31:0];
assign desc_15_axuser_11_axuser_f = desc_15_axuser_11_reg[31:0];
assign desc_15_axuser_12_axuser_f = desc_15_axuser_12_reg[31:0];
assign desc_15_axuser_13_axuser_f = desc_15_axuser_13_reg[31:0];
assign desc_15_axuser_14_axuser_f = desc_15_axuser_14_reg[31:0];
assign desc_15_axuser_15_axuser_f = desc_15_axuser_15_reg[31:0];
assign desc_15_size_txn_size_f = desc_15_size_reg[15:0];
assign desc_15_axsize_axsize_f = desc_15_axsize_reg[2:0];
assign desc_15_axaddr_0_addr_f = desc_15_axaddr_0_reg[31:0];
assign desc_15_axaddr_1_addr_f = desc_15_axaddr_1_reg[31:0];
assign desc_15_axaddr_2_addr_f = desc_15_axaddr_2_reg[31:0];
assign desc_15_axaddr_3_addr_f = desc_15_axaddr_3_reg[31:0];
assign desc_15_data_offset_addr_f = desc_15_data_offset_reg[31:0];
assign desc_15_wuser_0_wuser_f = desc_15_wuser_0_reg[31:0];
assign desc_15_wuser_1_wuser_f = desc_15_wuser_1_reg[31:0];
assign desc_15_wuser_2_wuser_f = desc_15_wuser_2_reg[31:0];
assign desc_15_wuser_3_wuser_f = desc_15_wuser_3_reg[31:0];
assign desc_15_wuser_4_wuser_f = desc_15_wuser_4_reg[31:0];
assign desc_15_wuser_5_wuser_f = desc_15_wuser_5_reg[31:0];
assign desc_15_wuser_6_wuser_f = desc_15_wuser_6_reg[31:0];
assign desc_15_wuser_7_wuser_f = desc_15_wuser_7_reg[31:0];
assign desc_15_wuser_8_wuser_f = desc_15_wuser_8_reg[31:0];
assign desc_15_wuser_9_wuser_f = desc_15_wuser_9_reg[31:0];
assign desc_15_wuser_10_wuser_f = desc_15_wuser_10_reg[31:0];
assign desc_15_wuser_11_wuser_f = desc_15_wuser_11_reg[31:0];
assign desc_15_wuser_12_wuser_f = desc_15_wuser_12_reg[31:0];
assign desc_15_wuser_13_wuser_f = desc_15_wuser_13_reg[31:0];
assign desc_15_wuser_14_wuser_f = desc_15_wuser_14_reg[31:0];
assign desc_15_wuser_15_wuser_f = desc_15_wuser_15_reg[31:0];
assign desc_15_data_host_addr_0_addr_f = desc_15_data_host_addr_0_reg[31:0];
assign desc_15_data_host_addr_1_addr_f = desc_15_data_host_addr_1_reg[31:0];
assign desc_15_data_host_addr_2_addr_f = desc_15_data_host_addr_2_reg[31:0];
assign desc_15_data_host_addr_3_addr_f = desc_15_data_host_addr_3_reg[31:0];
assign desc_15_wstrb_host_addr_0_addr_f = desc_15_wstrb_host_addr_0_reg[31:0];
assign desc_15_wstrb_host_addr_1_addr_f = desc_15_wstrb_host_addr_1_reg[31:0];
assign desc_15_wstrb_host_addr_2_addr_f = desc_15_wstrb_host_addr_2_reg[31:0];
assign desc_15_wstrb_host_addr_3_addr_f = desc_15_wstrb_host_addr_3_reg[31:0];
assign desc_15_xuser_0_xuser_f = desc_15_xuser_0_reg[31:0];
assign desc_15_xuser_1_xuser_f = desc_15_xuser_1_reg[31:0];
assign desc_15_xuser_2_xuser_f = desc_15_xuser_2_reg[31:0];
assign desc_15_xuser_3_xuser_f = desc_15_xuser_3_reg[31:0];
assign desc_15_xuser_4_xuser_f = desc_15_xuser_4_reg[31:0];
assign desc_15_xuser_5_xuser_f = desc_15_xuser_5_reg[31:0];
assign desc_15_xuser_6_xuser_f = desc_15_xuser_6_reg[31:0];
assign desc_15_xuser_7_xuser_f = desc_15_xuser_7_reg[31:0];
assign desc_15_xuser_8_xuser_f = desc_15_xuser_8_reg[31:0];
assign desc_15_xuser_9_xuser_f = desc_15_xuser_9_reg[31:0];
assign desc_15_xuser_10_xuser_f = desc_15_xuser_10_reg[31:0];
assign desc_15_xuser_11_xuser_f = desc_15_xuser_11_reg[31:0];
assign desc_15_xuser_12_xuser_f = desc_15_xuser_12_reg[31:0];
assign desc_15_xuser_13_xuser_f = desc_15_xuser_13_reg[31:0];
assign desc_15_xuser_14_xuser_f = desc_15_xuser_14_reg[31:0];
assign desc_15_xuser_15_xuser_f = desc_15_xuser_15_reg[31:0];


//////////////////////
//Assign signals to use in entire slave RTL ( int_<reg>_<field> )
//////////////////////

assign int_version_major_ver = version_major_ver_f;
assign int_version_minor_ver = version_minor_ver_f;
assign int_bridge_type_type = bridge_type_type_f;
assign int_axi_bridge_config_user_width = axi_bridge_config_user_width_f;
assign int_axi_bridge_config_id_width = axi_bridge_config_id_width_f;
assign int_axi_bridge_config_data_width = axi_bridge_config_data_width_f;
assign int_reset_dut_srst_3 = reset_dut_srst_3_f;
assign int_reset_dut_srst_2 = reset_dut_srst_2_f;
assign int_reset_dut_srst_1 = reset_dut_srst_1_f;
assign int_reset_dut_srst_0 = reset_dut_srst_0_f;
assign int_reset_srst = reset_srst_f;
assign int_mode_select_imm_bresp = mode_select_imm_bresp_f;
assign int_mode_select_mode_2 = mode_select_mode_2_f;
assign int_mode_select_mode_0_1 = mode_select_mode_0_1_f;
assign int_ownership_flip_flip = ownership_flip_flip_f;
assign int_status_resp_comp_resp_comp = status_resp_comp_resp_comp_f;
assign int_status_resp_resp = status_resp_resp_f;
assign int_intr_status_comp = intr_status_comp_f;
assign int_intr_status_c2h = intr_status_c2h_f;
assign int_intr_status_error = intr_status_error_f;
assign int_intr_status_txn_avail = intr_status_txn_avail_f;
assign int_intr_txn_avail_clear_clr_avail = intr_txn_avail_clear_clr_avail_f;
assign int_intr_txn_avail_enable_en_avail = intr_txn_avail_enable_en_avail_f;
assign int_intr_comp_clear_clr_comp = intr_comp_clear_clr_comp_f;
assign int_intr_comp_enable_en_comp = intr_comp_enable_en_comp_f;
assign int_intr_error_clear_clr_err_2 = intr_error_clear_clr_err_2_f;
assign int_intr_error_clear_clr_err_1 = intr_error_clear_clr_err_1_f;
assign int_intr_error_clear_clr_err_0 = intr_error_clear_clr_err_0_f;
assign int_intr_error_enable_en_err_2 = intr_error_enable_en_err_2_f;
assign int_intr_error_enable_en_err_1 = intr_error_enable_en_err_1_f;
assign int_intr_error_enable_en_err_0 = intr_error_enable_en_err_0_f;
assign int_intr_h2c_0_h2c = intr_h2c_0_h2c_f;
assign int_intr_h2c_1_h2c = intr_h2c_1_h2c_f;
assign int_intr_c2h_0_status_c2h = intr_c2h_0_status_c2h_f;
assign int_intr_c2h_1_status_c2h = intr_c2h_1_status_c2h_f;
assign int_c2h_gpio_0_status_gpio = c2h_gpio_0_status_gpio_f;
assign int_c2h_gpio_1_status_gpio = c2h_gpio_1_status_gpio_f;
assign int_c2h_gpio_2_status_gpio = c2h_gpio_2_status_gpio_f;
assign int_c2h_gpio_3_status_gpio = c2h_gpio_3_status_gpio_f;
assign int_c2h_gpio_4_status_gpio = c2h_gpio_4_status_gpio_f;
assign int_c2h_gpio_5_status_gpio = c2h_gpio_5_status_gpio_f;
assign int_c2h_gpio_6_status_gpio = c2h_gpio_6_status_gpio_f;
assign int_c2h_gpio_7_status_gpio = c2h_gpio_7_status_gpio_f;
assign int_c2h_gpio_8_status_gpio = c2h_gpio_8_status_gpio_f;
assign int_c2h_gpio_9_status_gpio = c2h_gpio_9_status_gpio_f;
assign int_c2h_gpio_10_status_gpio = c2h_gpio_10_status_gpio_f;
assign int_c2h_gpio_11_status_gpio = c2h_gpio_11_status_gpio_f;
assign int_c2h_gpio_12_status_gpio = c2h_gpio_12_status_gpio_f;
assign int_c2h_gpio_13_status_gpio = c2h_gpio_13_status_gpio_f;
assign int_c2h_gpio_14_status_gpio = c2h_gpio_14_status_gpio_f;
assign int_c2h_gpio_15_status_gpio = c2h_gpio_15_status_gpio_f;
assign int_addr_in_0_addr = addr_in_0_addr_f;
assign int_addr_in_1_addr = addr_in_1_addr_f;
assign int_addr_in_2_addr = addr_in_2_addr_f;
assign int_addr_in_3_addr = addr_in_3_addr_f;
assign int_trans_mask_0_addr = trans_mask_0_addr_f;
assign int_trans_mask_1_addr = trans_mask_1_addr_f;
assign int_trans_mask_2_addr = trans_mask_2_addr_f;
assign int_trans_mask_3_addr = trans_mask_3_addr_f;
assign int_trans_addr_0_addr = trans_addr_0_addr_f;
assign int_trans_addr_1_addr = trans_addr_1_addr_f;
assign int_trans_addr_2_addr = trans_addr_2_addr_f;
assign int_trans_addr_3_addr = trans_addr_3_addr_f;
assign int_resp_order_field = resp_order_field_f;

assign int_desc_0_data_host_addr_0_addr = desc_0_data_host_addr_0_addr_f;
assign int_desc_0_data_host_addr_1_addr = desc_0_data_host_addr_1_addr_f;
assign int_desc_0_data_host_addr_2_addr = desc_0_data_host_addr_2_addr_f;
assign int_desc_0_data_host_addr_3_addr = desc_0_data_host_addr_3_addr_f;
assign int_desc_0_wstrb_host_addr_0_addr = desc_0_wstrb_host_addr_0_addr_f;
assign int_desc_0_wstrb_host_addr_1_addr = desc_0_wstrb_host_addr_1_addr_f;
assign int_desc_0_wstrb_host_addr_2_addr = desc_0_wstrb_host_addr_2_addr_f;
assign int_desc_0_wstrb_host_addr_3_addr = desc_0_wstrb_host_addr_3_addr_f;
assign int_desc_1_data_host_addr_0_addr = desc_1_data_host_addr_0_addr_f;
assign int_desc_1_data_host_addr_1_addr = desc_1_data_host_addr_1_addr_f;
assign int_desc_1_data_host_addr_2_addr = desc_1_data_host_addr_2_addr_f;
assign int_desc_1_data_host_addr_3_addr = desc_1_data_host_addr_3_addr_f;
assign int_desc_1_wstrb_host_addr_0_addr = desc_1_wstrb_host_addr_0_addr_f;
assign int_desc_1_wstrb_host_addr_1_addr = desc_1_wstrb_host_addr_1_addr_f;
assign int_desc_1_wstrb_host_addr_2_addr = desc_1_wstrb_host_addr_2_addr_f;
assign int_desc_1_wstrb_host_addr_3_addr = desc_1_wstrb_host_addr_3_addr_f;
assign int_desc_2_data_host_addr_0_addr = desc_2_data_host_addr_0_addr_f;
assign int_desc_2_data_host_addr_1_addr = desc_2_data_host_addr_1_addr_f;
assign int_desc_2_data_host_addr_2_addr = desc_2_data_host_addr_2_addr_f;
assign int_desc_2_data_host_addr_3_addr = desc_2_data_host_addr_3_addr_f;
assign int_desc_2_wstrb_host_addr_0_addr = desc_2_wstrb_host_addr_0_addr_f;
assign int_desc_2_wstrb_host_addr_1_addr = desc_2_wstrb_host_addr_1_addr_f;
assign int_desc_2_wstrb_host_addr_2_addr = desc_2_wstrb_host_addr_2_addr_f;
assign int_desc_2_wstrb_host_addr_3_addr = desc_2_wstrb_host_addr_3_addr_f;
assign int_desc_3_data_host_addr_0_addr = desc_3_data_host_addr_0_addr_f;
assign int_desc_3_data_host_addr_1_addr = desc_3_data_host_addr_1_addr_f;
assign int_desc_3_data_host_addr_2_addr = desc_3_data_host_addr_2_addr_f;
assign int_desc_3_data_host_addr_3_addr = desc_3_data_host_addr_3_addr_f;
assign int_desc_3_wstrb_host_addr_0_addr = desc_3_wstrb_host_addr_0_addr_f;
assign int_desc_3_wstrb_host_addr_1_addr = desc_3_wstrb_host_addr_1_addr_f;
assign int_desc_3_wstrb_host_addr_2_addr = desc_3_wstrb_host_addr_2_addr_f;
assign int_desc_3_wstrb_host_addr_3_addr = desc_3_wstrb_host_addr_3_addr_f;
assign int_desc_4_data_host_addr_0_addr = desc_4_data_host_addr_0_addr_f;
assign int_desc_4_data_host_addr_1_addr = desc_4_data_host_addr_1_addr_f;
assign int_desc_4_data_host_addr_2_addr = desc_4_data_host_addr_2_addr_f;
assign int_desc_4_data_host_addr_3_addr = desc_4_data_host_addr_3_addr_f;
assign int_desc_4_wstrb_host_addr_0_addr = desc_4_wstrb_host_addr_0_addr_f;
assign int_desc_4_wstrb_host_addr_1_addr = desc_4_wstrb_host_addr_1_addr_f;
assign int_desc_4_wstrb_host_addr_2_addr = desc_4_wstrb_host_addr_2_addr_f;
assign int_desc_4_wstrb_host_addr_3_addr = desc_4_wstrb_host_addr_3_addr_f;
assign int_desc_5_data_host_addr_0_addr = desc_5_data_host_addr_0_addr_f;
assign int_desc_5_data_host_addr_1_addr = desc_5_data_host_addr_1_addr_f;
assign int_desc_5_data_host_addr_2_addr = desc_5_data_host_addr_2_addr_f;
assign int_desc_5_data_host_addr_3_addr = desc_5_data_host_addr_3_addr_f;
assign int_desc_5_wstrb_host_addr_0_addr = desc_5_wstrb_host_addr_0_addr_f;
assign int_desc_5_wstrb_host_addr_1_addr = desc_5_wstrb_host_addr_1_addr_f;
assign int_desc_5_wstrb_host_addr_2_addr = desc_5_wstrb_host_addr_2_addr_f;
assign int_desc_5_wstrb_host_addr_3_addr = desc_5_wstrb_host_addr_3_addr_f;
assign int_desc_6_data_host_addr_0_addr = desc_6_data_host_addr_0_addr_f;
assign int_desc_6_data_host_addr_1_addr = desc_6_data_host_addr_1_addr_f;
assign int_desc_6_data_host_addr_2_addr = desc_6_data_host_addr_2_addr_f;
assign int_desc_6_data_host_addr_3_addr = desc_6_data_host_addr_3_addr_f;
assign int_desc_6_wstrb_host_addr_0_addr = desc_6_wstrb_host_addr_0_addr_f;
assign int_desc_6_wstrb_host_addr_1_addr = desc_6_wstrb_host_addr_1_addr_f;
assign int_desc_6_wstrb_host_addr_2_addr = desc_6_wstrb_host_addr_2_addr_f;
assign int_desc_6_wstrb_host_addr_3_addr = desc_6_wstrb_host_addr_3_addr_f;
assign int_desc_7_data_host_addr_0_addr = desc_7_data_host_addr_0_addr_f;
assign int_desc_7_data_host_addr_1_addr = desc_7_data_host_addr_1_addr_f;
assign int_desc_7_data_host_addr_2_addr = desc_7_data_host_addr_2_addr_f;
assign int_desc_7_data_host_addr_3_addr = desc_7_data_host_addr_3_addr_f;
assign int_desc_7_wstrb_host_addr_0_addr = desc_7_wstrb_host_addr_0_addr_f;
assign int_desc_7_wstrb_host_addr_1_addr = desc_7_wstrb_host_addr_1_addr_f;
assign int_desc_7_wstrb_host_addr_2_addr = desc_7_wstrb_host_addr_2_addr_f;
assign int_desc_7_wstrb_host_addr_3_addr = desc_7_wstrb_host_addr_3_addr_f;
assign int_desc_8_data_host_addr_0_addr = desc_8_data_host_addr_0_addr_f;
assign int_desc_8_data_host_addr_1_addr = desc_8_data_host_addr_1_addr_f;
assign int_desc_8_data_host_addr_2_addr = desc_8_data_host_addr_2_addr_f;
assign int_desc_8_data_host_addr_3_addr = desc_8_data_host_addr_3_addr_f;
assign int_desc_8_wstrb_host_addr_0_addr = desc_8_wstrb_host_addr_0_addr_f;
assign int_desc_8_wstrb_host_addr_1_addr = desc_8_wstrb_host_addr_1_addr_f;
assign int_desc_8_wstrb_host_addr_2_addr = desc_8_wstrb_host_addr_2_addr_f;
assign int_desc_8_wstrb_host_addr_3_addr = desc_8_wstrb_host_addr_3_addr_f;
assign int_desc_9_data_host_addr_0_addr = desc_9_data_host_addr_0_addr_f;
assign int_desc_9_data_host_addr_1_addr = desc_9_data_host_addr_1_addr_f;
assign int_desc_9_data_host_addr_2_addr = desc_9_data_host_addr_2_addr_f;
assign int_desc_9_data_host_addr_3_addr = desc_9_data_host_addr_3_addr_f;
assign int_desc_9_wstrb_host_addr_0_addr = desc_9_wstrb_host_addr_0_addr_f;
assign int_desc_9_wstrb_host_addr_1_addr = desc_9_wstrb_host_addr_1_addr_f;
assign int_desc_9_wstrb_host_addr_2_addr = desc_9_wstrb_host_addr_2_addr_f;
assign int_desc_9_wstrb_host_addr_3_addr = desc_9_wstrb_host_addr_3_addr_f;
assign int_desc_10_data_host_addr_0_addr = desc_10_data_host_addr_0_addr_f;
assign int_desc_10_data_host_addr_1_addr = desc_10_data_host_addr_1_addr_f;
assign int_desc_10_data_host_addr_2_addr = desc_10_data_host_addr_2_addr_f;
assign int_desc_10_data_host_addr_3_addr = desc_10_data_host_addr_3_addr_f;
assign int_desc_10_wstrb_host_addr_0_addr = desc_10_wstrb_host_addr_0_addr_f;
assign int_desc_10_wstrb_host_addr_1_addr = desc_10_wstrb_host_addr_1_addr_f;
assign int_desc_10_wstrb_host_addr_2_addr = desc_10_wstrb_host_addr_2_addr_f;
assign int_desc_10_wstrb_host_addr_3_addr = desc_10_wstrb_host_addr_3_addr_f;
assign int_desc_11_data_host_addr_0_addr = desc_11_data_host_addr_0_addr_f;
assign int_desc_11_data_host_addr_1_addr = desc_11_data_host_addr_1_addr_f;
assign int_desc_11_data_host_addr_2_addr = desc_11_data_host_addr_2_addr_f;
assign int_desc_11_data_host_addr_3_addr = desc_11_data_host_addr_3_addr_f;
assign int_desc_11_wstrb_host_addr_0_addr = desc_11_wstrb_host_addr_0_addr_f;
assign int_desc_11_wstrb_host_addr_1_addr = desc_11_wstrb_host_addr_1_addr_f;
assign int_desc_11_wstrb_host_addr_2_addr = desc_11_wstrb_host_addr_2_addr_f;
assign int_desc_11_wstrb_host_addr_3_addr = desc_11_wstrb_host_addr_3_addr_f;
assign int_desc_12_data_host_addr_0_addr = desc_12_data_host_addr_0_addr_f;
assign int_desc_12_data_host_addr_1_addr = desc_12_data_host_addr_1_addr_f;
assign int_desc_12_data_host_addr_2_addr = desc_12_data_host_addr_2_addr_f;
assign int_desc_12_data_host_addr_3_addr = desc_12_data_host_addr_3_addr_f;
assign int_desc_12_wstrb_host_addr_0_addr = desc_12_wstrb_host_addr_0_addr_f;
assign int_desc_12_wstrb_host_addr_1_addr = desc_12_wstrb_host_addr_1_addr_f;
assign int_desc_12_wstrb_host_addr_2_addr = desc_12_wstrb_host_addr_2_addr_f;
assign int_desc_12_wstrb_host_addr_3_addr = desc_12_wstrb_host_addr_3_addr_f;
assign int_desc_13_data_host_addr_0_addr = desc_13_data_host_addr_0_addr_f;
assign int_desc_13_data_host_addr_1_addr = desc_13_data_host_addr_1_addr_f;
assign int_desc_13_data_host_addr_2_addr = desc_13_data_host_addr_2_addr_f;
assign int_desc_13_data_host_addr_3_addr = desc_13_data_host_addr_3_addr_f;
assign int_desc_13_wstrb_host_addr_0_addr = desc_13_wstrb_host_addr_0_addr_f;
assign int_desc_13_wstrb_host_addr_1_addr = desc_13_wstrb_host_addr_1_addr_f;
assign int_desc_13_wstrb_host_addr_2_addr = desc_13_wstrb_host_addr_2_addr_f;
assign int_desc_13_wstrb_host_addr_3_addr = desc_13_wstrb_host_addr_3_addr_f;
assign int_desc_14_data_host_addr_0_addr = desc_14_data_host_addr_0_addr_f;
assign int_desc_14_data_host_addr_1_addr = desc_14_data_host_addr_1_addr_f;
assign int_desc_14_data_host_addr_2_addr = desc_14_data_host_addr_2_addr_f;
assign int_desc_14_data_host_addr_3_addr = desc_14_data_host_addr_3_addr_f;
assign int_desc_14_wstrb_host_addr_0_addr = desc_14_wstrb_host_addr_0_addr_f;
assign int_desc_14_wstrb_host_addr_1_addr = desc_14_wstrb_host_addr_1_addr_f;
assign int_desc_14_wstrb_host_addr_2_addr = desc_14_wstrb_host_addr_2_addr_f;
assign int_desc_14_wstrb_host_addr_3_addr = desc_14_wstrb_host_addr_3_addr_f;
assign int_desc_15_data_host_addr_0_addr = desc_15_data_host_addr_0_addr_f;
assign int_desc_15_data_host_addr_1_addr = desc_15_data_host_addr_1_addr_f;
assign int_desc_15_data_host_addr_2_addr = desc_15_data_host_addr_2_addr_f;
assign int_desc_15_data_host_addr_3_addr = desc_15_data_host_addr_3_addr_f;
assign int_desc_15_wstrb_host_addr_0_addr = desc_15_wstrb_host_addr_0_addr_f;
assign int_desc_15_wstrb_host_addr_1_addr = desc_15_wstrb_host_addr_1_addr_f;
assign int_desc_15_wstrb_host_addr_2_addr = desc_15_wstrb_host_addr_2_addr_f;
assign int_desc_15_wstrb_host_addr_3_addr = desc_15_wstrb_host_addr_3_addr_f;
assign int_desc_0_xuser_0_xuser = desc_0_xuser_0_xuser_f;
assign int_desc_0_xuser_1_xuser = desc_0_xuser_1_xuser_f;
assign int_desc_0_xuser_2_xuser = desc_0_xuser_2_xuser_f;
assign int_desc_0_xuser_3_xuser = desc_0_xuser_3_xuser_f;
assign int_desc_0_xuser_4_xuser = desc_0_xuser_4_xuser_f;
assign int_desc_0_xuser_5_xuser = desc_0_xuser_5_xuser_f;
assign int_desc_0_xuser_6_xuser = desc_0_xuser_6_xuser_f;
assign int_desc_0_xuser_7_xuser = desc_0_xuser_7_xuser_f;
assign int_desc_0_xuser_8_xuser = desc_0_xuser_8_xuser_f;
assign int_desc_0_xuser_9_xuser = desc_0_xuser_9_xuser_f;
assign int_desc_0_xuser_10_xuser = desc_0_xuser_10_xuser_f;
assign int_desc_0_xuser_11_xuser = desc_0_xuser_11_xuser_f;
assign int_desc_0_xuser_12_xuser = desc_0_xuser_12_xuser_f;
assign int_desc_0_xuser_13_xuser = desc_0_xuser_13_xuser_f;
assign int_desc_0_xuser_14_xuser = desc_0_xuser_14_xuser_f;
assign int_desc_0_xuser_15_xuser = desc_0_xuser_15_xuser_f;
assign int_desc_1_xuser_0_xuser = desc_1_xuser_0_xuser_f;
assign int_desc_1_xuser_1_xuser = desc_1_xuser_1_xuser_f;
assign int_desc_1_xuser_2_xuser = desc_1_xuser_2_xuser_f;
assign int_desc_1_xuser_3_xuser = desc_1_xuser_3_xuser_f;
assign int_desc_1_xuser_4_xuser = desc_1_xuser_4_xuser_f;
assign int_desc_1_xuser_5_xuser = desc_1_xuser_5_xuser_f;
assign int_desc_1_xuser_6_xuser = desc_1_xuser_6_xuser_f;
assign int_desc_1_xuser_7_xuser = desc_1_xuser_7_xuser_f;
assign int_desc_1_xuser_8_xuser = desc_1_xuser_8_xuser_f;
assign int_desc_1_xuser_9_xuser = desc_1_xuser_9_xuser_f;
assign int_desc_1_xuser_10_xuser = desc_1_xuser_10_xuser_f;
assign int_desc_1_xuser_11_xuser = desc_1_xuser_11_xuser_f;
assign int_desc_1_xuser_12_xuser = desc_1_xuser_12_xuser_f;
assign int_desc_1_xuser_13_xuser = desc_1_xuser_13_xuser_f;
assign int_desc_1_xuser_14_xuser = desc_1_xuser_14_xuser_f;
assign int_desc_1_xuser_15_xuser = desc_1_xuser_15_xuser_f;
assign int_desc_2_xuser_0_xuser = desc_2_xuser_0_xuser_f;
assign int_desc_2_xuser_1_xuser = desc_2_xuser_1_xuser_f;
assign int_desc_2_xuser_2_xuser = desc_2_xuser_2_xuser_f;
assign int_desc_2_xuser_3_xuser = desc_2_xuser_3_xuser_f;
assign int_desc_2_xuser_4_xuser = desc_2_xuser_4_xuser_f;
assign int_desc_2_xuser_5_xuser = desc_2_xuser_5_xuser_f;
assign int_desc_2_xuser_6_xuser = desc_2_xuser_6_xuser_f;
assign int_desc_2_xuser_7_xuser = desc_2_xuser_7_xuser_f;
assign int_desc_2_xuser_8_xuser = desc_2_xuser_8_xuser_f;
assign int_desc_2_xuser_9_xuser = desc_2_xuser_9_xuser_f;
assign int_desc_2_xuser_10_xuser = desc_2_xuser_10_xuser_f;
assign int_desc_2_xuser_11_xuser = desc_2_xuser_11_xuser_f;
assign int_desc_2_xuser_12_xuser = desc_2_xuser_12_xuser_f;
assign int_desc_2_xuser_13_xuser = desc_2_xuser_13_xuser_f;
assign int_desc_2_xuser_14_xuser = desc_2_xuser_14_xuser_f;
assign int_desc_2_xuser_15_xuser = desc_2_xuser_15_xuser_f;
assign int_desc_3_xuser_0_xuser = desc_3_xuser_0_xuser_f;
assign int_desc_3_xuser_1_xuser = desc_3_xuser_1_xuser_f;
assign int_desc_3_xuser_2_xuser = desc_3_xuser_2_xuser_f;
assign int_desc_3_xuser_3_xuser = desc_3_xuser_3_xuser_f;
assign int_desc_3_xuser_4_xuser = desc_3_xuser_4_xuser_f;
assign int_desc_3_xuser_5_xuser = desc_3_xuser_5_xuser_f;
assign int_desc_3_xuser_6_xuser = desc_3_xuser_6_xuser_f;
assign int_desc_3_xuser_7_xuser = desc_3_xuser_7_xuser_f;
assign int_desc_3_xuser_8_xuser = desc_3_xuser_8_xuser_f;
assign int_desc_3_xuser_9_xuser = desc_3_xuser_9_xuser_f;
assign int_desc_3_xuser_10_xuser = desc_3_xuser_10_xuser_f;
assign int_desc_3_xuser_11_xuser = desc_3_xuser_11_xuser_f;
assign int_desc_3_xuser_12_xuser = desc_3_xuser_12_xuser_f;
assign int_desc_3_xuser_13_xuser = desc_3_xuser_13_xuser_f;
assign int_desc_3_xuser_14_xuser = desc_3_xuser_14_xuser_f;
assign int_desc_3_xuser_15_xuser = desc_3_xuser_15_xuser_f;
assign int_desc_4_xuser_0_xuser = desc_4_xuser_0_xuser_f;
assign int_desc_4_xuser_1_xuser = desc_4_xuser_1_xuser_f;
assign int_desc_4_xuser_2_xuser = desc_4_xuser_2_xuser_f;
assign int_desc_4_xuser_3_xuser = desc_4_xuser_3_xuser_f;
assign int_desc_4_xuser_4_xuser = desc_4_xuser_4_xuser_f;
assign int_desc_4_xuser_5_xuser = desc_4_xuser_5_xuser_f;
assign int_desc_4_xuser_6_xuser = desc_4_xuser_6_xuser_f;
assign int_desc_4_xuser_7_xuser = desc_4_xuser_7_xuser_f;
assign int_desc_4_xuser_8_xuser = desc_4_xuser_8_xuser_f;
assign int_desc_4_xuser_9_xuser = desc_4_xuser_9_xuser_f;
assign int_desc_4_xuser_10_xuser = desc_4_xuser_10_xuser_f;
assign int_desc_4_xuser_11_xuser = desc_4_xuser_11_xuser_f;
assign int_desc_4_xuser_12_xuser = desc_4_xuser_12_xuser_f;
assign int_desc_4_xuser_13_xuser = desc_4_xuser_13_xuser_f;
assign int_desc_4_xuser_14_xuser = desc_4_xuser_14_xuser_f;
assign int_desc_4_xuser_15_xuser = desc_4_xuser_15_xuser_f;
assign int_desc_5_xuser_0_xuser = desc_5_xuser_0_xuser_f;
assign int_desc_5_xuser_1_xuser = desc_5_xuser_1_xuser_f;
assign int_desc_5_xuser_2_xuser = desc_5_xuser_2_xuser_f;
assign int_desc_5_xuser_3_xuser = desc_5_xuser_3_xuser_f;
assign int_desc_5_xuser_4_xuser = desc_5_xuser_4_xuser_f;
assign int_desc_5_xuser_5_xuser = desc_5_xuser_5_xuser_f;
assign int_desc_5_xuser_6_xuser = desc_5_xuser_6_xuser_f;
assign int_desc_5_xuser_7_xuser = desc_5_xuser_7_xuser_f;
assign int_desc_5_xuser_8_xuser = desc_5_xuser_8_xuser_f;
assign int_desc_5_xuser_9_xuser = desc_5_xuser_9_xuser_f;
assign int_desc_5_xuser_10_xuser = desc_5_xuser_10_xuser_f;
assign int_desc_5_xuser_11_xuser = desc_5_xuser_11_xuser_f;
assign int_desc_5_xuser_12_xuser = desc_5_xuser_12_xuser_f;
assign int_desc_5_xuser_13_xuser = desc_5_xuser_13_xuser_f;
assign int_desc_5_xuser_14_xuser = desc_5_xuser_14_xuser_f;
assign int_desc_5_xuser_15_xuser = desc_5_xuser_15_xuser_f;
assign int_desc_6_xuser_0_xuser = desc_6_xuser_0_xuser_f;
assign int_desc_6_xuser_1_xuser = desc_6_xuser_1_xuser_f;
assign int_desc_6_xuser_2_xuser = desc_6_xuser_2_xuser_f;
assign int_desc_6_xuser_3_xuser = desc_6_xuser_3_xuser_f;
assign int_desc_6_xuser_4_xuser = desc_6_xuser_4_xuser_f;
assign int_desc_6_xuser_5_xuser = desc_6_xuser_5_xuser_f;
assign int_desc_6_xuser_6_xuser = desc_6_xuser_6_xuser_f;
assign int_desc_6_xuser_7_xuser = desc_6_xuser_7_xuser_f;
assign int_desc_6_xuser_8_xuser = desc_6_xuser_8_xuser_f;
assign int_desc_6_xuser_9_xuser = desc_6_xuser_9_xuser_f;
assign int_desc_6_xuser_10_xuser = desc_6_xuser_10_xuser_f;
assign int_desc_6_xuser_11_xuser = desc_6_xuser_11_xuser_f;
assign int_desc_6_xuser_12_xuser = desc_6_xuser_12_xuser_f;
assign int_desc_6_xuser_13_xuser = desc_6_xuser_13_xuser_f;
assign int_desc_6_xuser_14_xuser = desc_6_xuser_14_xuser_f;
assign int_desc_6_xuser_15_xuser = desc_6_xuser_15_xuser_f;
assign int_desc_7_xuser_0_xuser = desc_7_xuser_0_xuser_f;
assign int_desc_7_xuser_1_xuser = desc_7_xuser_1_xuser_f;
assign int_desc_7_xuser_2_xuser = desc_7_xuser_2_xuser_f;
assign int_desc_7_xuser_3_xuser = desc_7_xuser_3_xuser_f;
assign int_desc_7_xuser_4_xuser = desc_7_xuser_4_xuser_f;
assign int_desc_7_xuser_5_xuser = desc_7_xuser_5_xuser_f;
assign int_desc_7_xuser_6_xuser = desc_7_xuser_6_xuser_f;
assign int_desc_7_xuser_7_xuser = desc_7_xuser_7_xuser_f;
assign int_desc_7_xuser_8_xuser = desc_7_xuser_8_xuser_f;
assign int_desc_7_xuser_9_xuser = desc_7_xuser_9_xuser_f;
assign int_desc_7_xuser_10_xuser = desc_7_xuser_10_xuser_f;
assign int_desc_7_xuser_11_xuser = desc_7_xuser_11_xuser_f;
assign int_desc_7_xuser_12_xuser = desc_7_xuser_12_xuser_f;
assign int_desc_7_xuser_13_xuser = desc_7_xuser_13_xuser_f;
assign int_desc_7_xuser_14_xuser = desc_7_xuser_14_xuser_f;
assign int_desc_7_xuser_15_xuser = desc_7_xuser_15_xuser_f;
assign int_desc_8_xuser_0_xuser = desc_8_xuser_0_xuser_f;
assign int_desc_8_xuser_1_xuser = desc_8_xuser_1_xuser_f;
assign int_desc_8_xuser_2_xuser = desc_8_xuser_2_xuser_f;
assign int_desc_8_xuser_3_xuser = desc_8_xuser_3_xuser_f;
assign int_desc_8_xuser_4_xuser = desc_8_xuser_4_xuser_f;
assign int_desc_8_xuser_5_xuser = desc_8_xuser_5_xuser_f;
assign int_desc_8_xuser_6_xuser = desc_8_xuser_6_xuser_f;
assign int_desc_8_xuser_7_xuser = desc_8_xuser_7_xuser_f;
assign int_desc_8_xuser_8_xuser = desc_8_xuser_8_xuser_f;
assign int_desc_8_xuser_9_xuser = desc_8_xuser_9_xuser_f;
assign int_desc_8_xuser_10_xuser = desc_8_xuser_10_xuser_f;
assign int_desc_8_xuser_11_xuser = desc_8_xuser_11_xuser_f;
assign int_desc_8_xuser_12_xuser = desc_8_xuser_12_xuser_f;
assign int_desc_8_xuser_13_xuser = desc_8_xuser_13_xuser_f;
assign int_desc_8_xuser_14_xuser = desc_8_xuser_14_xuser_f;
assign int_desc_8_xuser_15_xuser = desc_8_xuser_15_xuser_f;
assign int_desc_9_xuser_0_xuser = desc_9_xuser_0_xuser_f;
assign int_desc_9_xuser_1_xuser = desc_9_xuser_1_xuser_f;
assign int_desc_9_xuser_2_xuser = desc_9_xuser_2_xuser_f;
assign int_desc_9_xuser_3_xuser = desc_9_xuser_3_xuser_f;
assign int_desc_9_xuser_4_xuser = desc_9_xuser_4_xuser_f;
assign int_desc_9_xuser_5_xuser = desc_9_xuser_5_xuser_f;
assign int_desc_9_xuser_6_xuser = desc_9_xuser_6_xuser_f;
assign int_desc_9_xuser_7_xuser = desc_9_xuser_7_xuser_f;
assign int_desc_9_xuser_8_xuser = desc_9_xuser_8_xuser_f;
assign int_desc_9_xuser_9_xuser = desc_9_xuser_9_xuser_f;
assign int_desc_9_xuser_10_xuser = desc_9_xuser_10_xuser_f;
assign int_desc_9_xuser_11_xuser = desc_9_xuser_11_xuser_f;
assign int_desc_9_xuser_12_xuser = desc_9_xuser_12_xuser_f;
assign int_desc_9_xuser_13_xuser = desc_9_xuser_13_xuser_f;
assign int_desc_9_xuser_14_xuser = desc_9_xuser_14_xuser_f;
assign int_desc_9_xuser_15_xuser = desc_9_xuser_15_xuser_f;
assign int_desc_10_xuser_0_xuser = desc_10_xuser_0_xuser_f;
assign int_desc_10_xuser_1_xuser = desc_10_xuser_1_xuser_f;
assign int_desc_10_xuser_2_xuser = desc_10_xuser_2_xuser_f;
assign int_desc_10_xuser_3_xuser = desc_10_xuser_3_xuser_f;
assign int_desc_10_xuser_4_xuser = desc_10_xuser_4_xuser_f;
assign int_desc_10_xuser_5_xuser = desc_10_xuser_5_xuser_f;
assign int_desc_10_xuser_6_xuser = desc_10_xuser_6_xuser_f;
assign int_desc_10_xuser_7_xuser = desc_10_xuser_7_xuser_f;
assign int_desc_10_xuser_8_xuser = desc_10_xuser_8_xuser_f;
assign int_desc_10_xuser_9_xuser = desc_10_xuser_9_xuser_f;
assign int_desc_10_xuser_10_xuser = desc_10_xuser_10_xuser_f;
assign int_desc_10_xuser_11_xuser = desc_10_xuser_11_xuser_f;
assign int_desc_10_xuser_12_xuser = desc_10_xuser_12_xuser_f;
assign int_desc_10_xuser_13_xuser = desc_10_xuser_13_xuser_f;
assign int_desc_10_xuser_14_xuser = desc_10_xuser_14_xuser_f;
assign int_desc_10_xuser_15_xuser = desc_10_xuser_15_xuser_f;
assign int_desc_11_xuser_0_xuser = desc_11_xuser_0_xuser_f;
assign int_desc_11_xuser_1_xuser = desc_11_xuser_1_xuser_f;
assign int_desc_11_xuser_2_xuser = desc_11_xuser_2_xuser_f;
assign int_desc_11_xuser_3_xuser = desc_11_xuser_3_xuser_f;
assign int_desc_11_xuser_4_xuser = desc_11_xuser_4_xuser_f;
assign int_desc_11_xuser_5_xuser = desc_11_xuser_5_xuser_f;
assign int_desc_11_xuser_6_xuser = desc_11_xuser_6_xuser_f;
assign int_desc_11_xuser_7_xuser = desc_11_xuser_7_xuser_f;
assign int_desc_11_xuser_8_xuser = desc_11_xuser_8_xuser_f;
assign int_desc_11_xuser_9_xuser = desc_11_xuser_9_xuser_f;
assign int_desc_11_xuser_10_xuser = desc_11_xuser_10_xuser_f;
assign int_desc_11_xuser_11_xuser = desc_11_xuser_11_xuser_f;
assign int_desc_11_xuser_12_xuser = desc_11_xuser_12_xuser_f;
assign int_desc_11_xuser_13_xuser = desc_11_xuser_13_xuser_f;
assign int_desc_11_xuser_14_xuser = desc_11_xuser_14_xuser_f;
assign int_desc_11_xuser_15_xuser = desc_11_xuser_15_xuser_f;
assign int_desc_12_xuser_0_xuser = desc_12_xuser_0_xuser_f;
assign int_desc_12_xuser_1_xuser = desc_12_xuser_1_xuser_f;
assign int_desc_12_xuser_2_xuser = desc_12_xuser_2_xuser_f;
assign int_desc_12_xuser_3_xuser = desc_12_xuser_3_xuser_f;
assign int_desc_12_xuser_4_xuser = desc_12_xuser_4_xuser_f;
assign int_desc_12_xuser_5_xuser = desc_12_xuser_5_xuser_f;
assign int_desc_12_xuser_6_xuser = desc_12_xuser_6_xuser_f;
assign int_desc_12_xuser_7_xuser = desc_12_xuser_7_xuser_f;
assign int_desc_12_xuser_8_xuser = desc_12_xuser_8_xuser_f;
assign int_desc_12_xuser_9_xuser = desc_12_xuser_9_xuser_f;
assign int_desc_12_xuser_10_xuser = desc_12_xuser_10_xuser_f;
assign int_desc_12_xuser_11_xuser = desc_12_xuser_11_xuser_f;
assign int_desc_12_xuser_12_xuser = desc_12_xuser_12_xuser_f;
assign int_desc_12_xuser_13_xuser = desc_12_xuser_13_xuser_f;
assign int_desc_12_xuser_14_xuser = desc_12_xuser_14_xuser_f;
assign int_desc_12_xuser_15_xuser = desc_12_xuser_15_xuser_f;
assign int_desc_13_xuser_0_xuser = desc_13_xuser_0_xuser_f;
assign int_desc_13_xuser_1_xuser = desc_13_xuser_1_xuser_f;
assign int_desc_13_xuser_2_xuser = desc_13_xuser_2_xuser_f;
assign int_desc_13_xuser_3_xuser = desc_13_xuser_3_xuser_f;
assign int_desc_13_xuser_4_xuser = desc_13_xuser_4_xuser_f;
assign int_desc_13_xuser_5_xuser = desc_13_xuser_5_xuser_f;
assign int_desc_13_xuser_6_xuser = desc_13_xuser_6_xuser_f;
assign int_desc_13_xuser_7_xuser = desc_13_xuser_7_xuser_f;
assign int_desc_13_xuser_8_xuser = desc_13_xuser_8_xuser_f;
assign int_desc_13_xuser_9_xuser = desc_13_xuser_9_xuser_f;
assign int_desc_13_xuser_10_xuser = desc_13_xuser_10_xuser_f;
assign int_desc_13_xuser_11_xuser = desc_13_xuser_11_xuser_f;
assign int_desc_13_xuser_12_xuser = desc_13_xuser_12_xuser_f;
assign int_desc_13_xuser_13_xuser = desc_13_xuser_13_xuser_f;
assign int_desc_13_xuser_14_xuser = desc_13_xuser_14_xuser_f;
assign int_desc_13_xuser_15_xuser = desc_13_xuser_15_xuser_f;
assign int_desc_14_xuser_0_xuser = desc_14_xuser_0_xuser_f;
assign int_desc_14_xuser_1_xuser = desc_14_xuser_1_xuser_f;
assign int_desc_14_xuser_2_xuser = desc_14_xuser_2_xuser_f;
assign int_desc_14_xuser_3_xuser = desc_14_xuser_3_xuser_f;
assign int_desc_14_xuser_4_xuser = desc_14_xuser_4_xuser_f;
assign int_desc_14_xuser_5_xuser = desc_14_xuser_5_xuser_f;
assign int_desc_14_xuser_6_xuser = desc_14_xuser_6_xuser_f;
assign int_desc_14_xuser_7_xuser = desc_14_xuser_7_xuser_f;
assign int_desc_14_xuser_8_xuser = desc_14_xuser_8_xuser_f;
assign int_desc_14_xuser_9_xuser = desc_14_xuser_9_xuser_f;
assign int_desc_14_xuser_10_xuser = desc_14_xuser_10_xuser_f;
assign int_desc_14_xuser_11_xuser = desc_14_xuser_11_xuser_f;
assign int_desc_14_xuser_12_xuser = desc_14_xuser_12_xuser_f;
assign int_desc_14_xuser_13_xuser = desc_14_xuser_13_xuser_f;
assign int_desc_14_xuser_14_xuser = desc_14_xuser_14_xuser_f;
assign int_desc_14_xuser_15_xuser = desc_14_xuser_15_xuser_f;
assign int_desc_15_xuser_0_xuser = desc_15_xuser_0_xuser_f;
assign int_desc_15_xuser_1_xuser = desc_15_xuser_1_xuser_f;
assign int_desc_15_xuser_2_xuser = desc_15_xuser_2_xuser_f;
assign int_desc_15_xuser_3_xuser = desc_15_xuser_3_xuser_f;
assign int_desc_15_xuser_4_xuser = desc_15_xuser_4_xuser_f;
assign int_desc_15_xuser_5_xuser = desc_15_xuser_5_xuser_f;
assign int_desc_15_xuser_6_xuser = desc_15_xuser_6_xuser_f;
assign int_desc_15_xuser_7_xuser = desc_15_xuser_7_xuser_f;
assign int_desc_15_xuser_8_xuser = desc_15_xuser_8_xuser_f;
assign int_desc_15_xuser_9_xuser = desc_15_xuser_9_xuser_f;
assign int_desc_15_xuser_10_xuser = desc_15_xuser_10_xuser_f;
assign int_desc_15_xuser_11_xuser = desc_15_xuser_11_xuser_f;
assign int_desc_15_xuser_12_xuser = desc_15_xuser_12_xuser_f;
assign int_desc_15_xuser_13_xuser = desc_15_xuser_13_xuser_f;
assign int_desc_15_xuser_14_xuser = desc_15_xuser_14_xuser_f;
assign int_desc_15_xuser_15_xuser = desc_15_xuser_15_xuser_f;

//////////////////////
//Signals to be given as input to RB  
//////////////////////

assign uc2rb_ownership_reg[31:MAX_DESC] = {(32-MAX_DESC){1'b0}};
assign uc2rb_ownership_reg[MAX_DESC-1:0] = int_ownership_own;
assign uc2rb_intr_txn_avail_status_reg[31:MAX_DESC] = {(32-MAX_DESC){1'b0}};				
assign uc2rb_intr_txn_avail_status_reg[MAX_DESC-1:0] = int_intr_txn_avail_status_avail;				
assign uc2rb_intr_comp_status_reg[31:MAX_DESC] = {(32-MAX_DESC){1'b0}};				
assign uc2rb_intr_comp_status_reg[MAX_DESC-1:0] = int_intr_comp_status_comp;				
assign uc2rb_intr_error_status_reg[31:1] = 31'h0;	
assign uc2rb_intr_error_status_reg[0] = int_intr_error_status_err_0;	

assign uc2rb_status_busy_reg[31:MAX_DESC] = {(32-MAX_DESC){1'b0}};
assign uc2rb_status_busy_reg[MAX_DESC-1:0] = int_status_busy_busy;

assign uc2rb_resp_fifo_free_level_reg[31:(DESC_IDX_WIDTH+1)] = {(32-DESC_IDX_WIDTH-1){1'b0}};
assign uc2rb_resp_fifo_free_level_reg[DESC_IDX_WIDTH:0] = int_resp_fifo_free_level_level;

assign uc2rb_desc_0_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_0_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_0_size_reg[31:16] = 16'h0;
assign uc2rb_desc_0_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_0_txn_type_reg[1] = int_desc_0_txn_type_wr_strb;
assign uc2rb_desc_0_txn_type_reg[0] = int_desc_0_txn_type_wr_rd;
assign uc2rb_desc_0_attr_reg[18:15] = int_desc_0_attr_axregion;
assign uc2rb_desc_0_attr_reg[14:11] = int_desc_0_attr_axqos;
assign uc2rb_desc_0_attr_reg[10:8] = int_desc_0_attr_axprot;
assign uc2rb_desc_0_attr_reg[7:4] = int_desc_0_attr_axcache;
assign uc2rb_desc_0_attr_reg[3:2] = int_desc_0_attr_axlock;
assign uc2rb_desc_0_attr_reg[1:0] = int_desc_0_attr_axburst;
assign uc2rb_desc_0_axid_0_reg[31:0] = int_desc_0_axid_0_axid;
assign uc2rb_desc_0_axid_1_reg[31:0] = int_desc_0_axid_1_axid;
assign uc2rb_desc_0_axid_2_reg[31:0] = int_desc_0_axid_2_axid;
assign uc2rb_desc_0_axid_3_reg[31:0] = int_desc_0_axid_3_axid;
assign uc2rb_desc_0_axuser_0_reg[31:0] = int_desc_0_axuser_0_axuser;
assign uc2rb_desc_0_axuser_1_reg[31:0] = int_desc_0_axuser_1_axuser;
assign uc2rb_desc_0_axuser_2_reg[31:0] = int_desc_0_axuser_2_axuser;
assign uc2rb_desc_0_axuser_3_reg[31:0] = int_desc_0_axuser_3_axuser;
assign uc2rb_desc_0_axuser_4_reg[31:0] = int_desc_0_axuser_4_axuser;
assign uc2rb_desc_0_axuser_5_reg[31:0] = int_desc_0_axuser_5_axuser;
assign uc2rb_desc_0_axuser_6_reg[31:0] = int_desc_0_axuser_6_axuser;
assign uc2rb_desc_0_axuser_7_reg[31:0] = int_desc_0_axuser_7_axuser;
assign uc2rb_desc_0_axuser_8_reg[31:0] = int_desc_0_axuser_8_axuser;
assign uc2rb_desc_0_axuser_9_reg[31:0] = int_desc_0_axuser_9_axuser;
assign uc2rb_desc_0_axuser_10_reg[31:0] = int_desc_0_axuser_10_axuser;
assign uc2rb_desc_0_axuser_11_reg[31:0] = int_desc_0_axuser_11_axuser;
assign uc2rb_desc_0_axuser_12_reg[31:0] = int_desc_0_axuser_12_axuser;
assign uc2rb_desc_0_axuser_13_reg[31:0] = int_desc_0_axuser_13_axuser;
assign uc2rb_desc_0_axuser_14_reg[31:0] = int_desc_0_axuser_14_axuser;
assign uc2rb_desc_0_axuser_15_reg[31:0] = int_desc_0_axuser_15_axuser;
assign uc2rb_desc_0_size_reg[15:0] = int_desc_0_size_txn_size;
assign uc2rb_desc_0_axsize_reg[2:0] = int_desc_0_axsize_axsize;
assign uc2rb_desc_0_axaddr_0_reg[31:0] = int_desc_0_axaddr_0_addr;
assign uc2rb_desc_0_axaddr_1_reg[31:0] = int_desc_0_axaddr_1_addr;
assign uc2rb_desc_0_axaddr_2_reg[31:0] = int_desc_0_axaddr_2_addr;
assign uc2rb_desc_0_axaddr_3_reg[31:0] = int_desc_0_axaddr_3_addr;
assign uc2rb_desc_0_data_offset_reg[31:0] = int_desc_0_data_offset_addr;
assign uc2rb_desc_0_wuser_0_reg[31:0] = int_desc_0_wuser_0_wuser;
assign uc2rb_desc_0_wuser_1_reg[31:0] = int_desc_0_wuser_1_wuser;
assign uc2rb_desc_0_wuser_2_reg[31:0] = int_desc_0_wuser_2_wuser;
assign uc2rb_desc_0_wuser_3_reg[31:0] = int_desc_0_wuser_3_wuser;
assign uc2rb_desc_0_wuser_4_reg[31:0] = int_desc_0_wuser_4_wuser;
assign uc2rb_desc_0_wuser_5_reg[31:0] = int_desc_0_wuser_5_wuser;
assign uc2rb_desc_0_wuser_6_reg[31:0] = int_desc_0_wuser_6_wuser;
assign uc2rb_desc_0_wuser_7_reg[31:0] = int_desc_0_wuser_7_wuser;
assign uc2rb_desc_0_wuser_8_reg[31:0] = int_desc_0_wuser_8_wuser;
assign uc2rb_desc_0_wuser_9_reg[31:0] = int_desc_0_wuser_9_wuser;
assign uc2rb_desc_0_wuser_10_reg[31:0] = int_desc_0_wuser_10_wuser;
assign uc2rb_desc_0_wuser_11_reg[31:0] = int_desc_0_wuser_11_wuser;
assign uc2rb_desc_0_wuser_12_reg[31:0] = int_desc_0_wuser_12_wuser;
assign uc2rb_desc_0_wuser_13_reg[31:0] = int_desc_0_wuser_13_wuser;
assign uc2rb_desc_0_wuser_14_reg[31:0] = int_desc_0_wuser_14_wuser;
assign uc2rb_desc_0_wuser_15_reg[31:0] = int_desc_0_wuser_15_wuser;
assign uc2rb_desc_1_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_1_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_1_size_reg[31:16] = 16'h0;
assign uc2rb_desc_1_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_1_txn_type_reg[1] = int_desc_1_txn_type_wr_strb;
assign uc2rb_desc_1_txn_type_reg[0] = int_desc_1_txn_type_wr_rd;
assign uc2rb_desc_1_attr_reg[18:15] = int_desc_1_attr_axregion;
assign uc2rb_desc_1_attr_reg[14:11] = int_desc_1_attr_axqos;
assign uc2rb_desc_1_attr_reg[10:8] = int_desc_1_attr_axprot;
assign uc2rb_desc_1_attr_reg[7:4] = int_desc_1_attr_axcache;
assign uc2rb_desc_1_attr_reg[3:2] = int_desc_1_attr_axlock;
assign uc2rb_desc_1_attr_reg[1:0] = int_desc_1_attr_axburst;
assign uc2rb_desc_1_axid_0_reg[31:0] = int_desc_1_axid_0_axid;
assign uc2rb_desc_1_axid_1_reg[31:0] = int_desc_1_axid_1_axid;
assign uc2rb_desc_1_axid_2_reg[31:0] = int_desc_1_axid_2_axid;
assign uc2rb_desc_1_axid_3_reg[31:0] = int_desc_1_axid_3_axid;
assign uc2rb_desc_1_axuser_0_reg[31:0] = int_desc_1_axuser_0_axuser;
assign uc2rb_desc_1_axuser_1_reg[31:0] = int_desc_1_axuser_1_axuser;
assign uc2rb_desc_1_axuser_2_reg[31:0] = int_desc_1_axuser_2_axuser;
assign uc2rb_desc_1_axuser_3_reg[31:0] = int_desc_1_axuser_3_axuser;
assign uc2rb_desc_1_axuser_4_reg[31:0] = int_desc_1_axuser_4_axuser;
assign uc2rb_desc_1_axuser_5_reg[31:0] = int_desc_1_axuser_5_axuser;
assign uc2rb_desc_1_axuser_6_reg[31:0] = int_desc_1_axuser_6_axuser;
assign uc2rb_desc_1_axuser_7_reg[31:0] = int_desc_1_axuser_7_axuser;
assign uc2rb_desc_1_axuser_8_reg[31:0] = int_desc_1_axuser_8_axuser;
assign uc2rb_desc_1_axuser_9_reg[31:0] = int_desc_1_axuser_9_axuser;
assign uc2rb_desc_1_axuser_10_reg[31:0] = int_desc_1_axuser_10_axuser;
assign uc2rb_desc_1_axuser_11_reg[31:0] = int_desc_1_axuser_11_axuser;
assign uc2rb_desc_1_axuser_12_reg[31:0] = int_desc_1_axuser_12_axuser;
assign uc2rb_desc_1_axuser_13_reg[31:0] = int_desc_1_axuser_13_axuser;
assign uc2rb_desc_1_axuser_14_reg[31:0] = int_desc_1_axuser_14_axuser;
assign uc2rb_desc_1_axuser_15_reg[31:0] = int_desc_1_axuser_15_axuser;
assign uc2rb_desc_1_size_reg[15:0] = int_desc_1_size_txn_size;
assign uc2rb_desc_1_axsize_reg[2:0] = int_desc_1_axsize_axsize;
assign uc2rb_desc_1_axaddr_0_reg[31:0] = int_desc_1_axaddr_0_addr;
assign uc2rb_desc_1_axaddr_1_reg[31:0] = int_desc_1_axaddr_1_addr;
assign uc2rb_desc_1_axaddr_2_reg[31:0] = int_desc_1_axaddr_2_addr;
assign uc2rb_desc_1_axaddr_3_reg[31:0] = int_desc_1_axaddr_3_addr;
assign uc2rb_desc_1_data_offset_reg[31:0] = int_desc_1_data_offset_addr;
assign uc2rb_desc_1_wuser_0_reg[31:0] = int_desc_1_wuser_0_wuser;
assign uc2rb_desc_1_wuser_1_reg[31:0] = int_desc_1_wuser_1_wuser;
assign uc2rb_desc_1_wuser_2_reg[31:0] = int_desc_1_wuser_2_wuser;
assign uc2rb_desc_1_wuser_3_reg[31:0] = int_desc_1_wuser_3_wuser;
assign uc2rb_desc_1_wuser_4_reg[31:0] = int_desc_1_wuser_4_wuser;
assign uc2rb_desc_1_wuser_5_reg[31:0] = int_desc_1_wuser_5_wuser;
assign uc2rb_desc_1_wuser_6_reg[31:0] = int_desc_1_wuser_6_wuser;
assign uc2rb_desc_1_wuser_7_reg[31:0] = int_desc_1_wuser_7_wuser;
assign uc2rb_desc_1_wuser_8_reg[31:0] = int_desc_1_wuser_8_wuser;
assign uc2rb_desc_1_wuser_9_reg[31:0] = int_desc_1_wuser_9_wuser;
assign uc2rb_desc_1_wuser_10_reg[31:0] = int_desc_1_wuser_10_wuser;
assign uc2rb_desc_1_wuser_11_reg[31:0] = int_desc_1_wuser_11_wuser;
assign uc2rb_desc_1_wuser_12_reg[31:0] = int_desc_1_wuser_12_wuser;
assign uc2rb_desc_1_wuser_13_reg[31:0] = int_desc_1_wuser_13_wuser;
assign uc2rb_desc_1_wuser_14_reg[31:0] = int_desc_1_wuser_14_wuser;
assign uc2rb_desc_1_wuser_15_reg[31:0] = int_desc_1_wuser_15_wuser;
assign uc2rb_desc_2_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_2_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_2_size_reg[31:16] = 16'h0;
assign uc2rb_desc_2_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_2_txn_type_reg[1] = int_desc_2_txn_type_wr_strb;
assign uc2rb_desc_2_txn_type_reg[0] = int_desc_2_txn_type_wr_rd;
assign uc2rb_desc_2_attr_reg[18:15] = int_desc_2_attr_axregion;
assign uc2rb_desc_2_attr_reg[14:11] = int_desc_2_attr_axqos;
assign uc2rb_desc_2_attr_reg[10:8] = int_desc_2_attr_axprot;
assign uc2rb_desc_2_attr_reg[7:4] = int_desc_2_attr_axcache;
assign uc2rb_desc_2_attr_reg[3:2] = int_desc_2_attr_axlock;
assign uc2rb_desc_2_attr_reg[1:0] = int_desc_2_attr_axburst;
assign uc2rb_desc_2_axid_0_reg[31:0] = int_desc_2_axid_0_axid;
assign uc2rb_desc_2_axid_1_reg[31:0] = int_desc_2_axid_1_axid;
assign uc2rb_desc_2_axid_2_reg[31:0] = int_desc_2_axid_2_axid;
assign uc2rb_desc_2_axid_3_reg[31:0] = int_desc_2_axid_3_axid;
assign uc2rb_desc_2_axuser_0_reg[31:0] = int_desc_2_axuser_0_axuser;
assign uc2rb_desc_2_axuser_1_reg[31:0] = int_desc_2_axuser_1_axuser;
assign uc2rb_desc_2_axuser_2_reg[31:0] = int_desc_2_axuser_2_axuser;
assign uc2rb_desc_2_axuser_3_reg[31:0] = int_desc_2_axuser_3_axuser;
assign uc2rb_desc_2_axuser_4_reg[31:0] = int_desc_2_axuser_4_axuser;
assign uc2rb_desc_2_axuser_5_reg[31:0] = int_desc_2_axuser_5_axuser;
assign uc2rb_desc_2_axuser_6_reg[31:0] = int_desc_2_axuser_6_axuser;
assign uc2rb_desc_2_axuser_7_reg[31:0] = int_desc_2_axuser_7_axuser;
assign uc2rb_desc_2_axuser_8_reg[31:0] = int_desc_2_axuser_8_axuser;
assign uc2rb_desc_2_axuser_9_reg[31:0] = int_desc_2_axuser_9_axuser;
assign uc2rb_desc_2_axuser_10_reg[31:0] = int_desc_2_axuser_10_axuser;
assign uc2rb_desc_2_axuser_11_reg[31:0] = int_desc_2_axuser_11_axuser;
assign uc2rb_desc_2_axuser_12_reg[31:0] = int_desc_2_axuser_12_axuser;
assign uc2rb_desc_2_axuser_13_reg[31:0] = int_desc_2_axuser_13_axuser;
assign uc2rb_desc_2_axuser_14_reg[31:0] = int_desc_2_axuser_14_axuser;
assign uc2rb_desc_2_axuser_15_reg[31:0] = int_desc_2_axuser_15_axuser;
assign uc2rb_desc_2_size_reg[15:0] = int_desc_2_size_txn_size;
assign uc2rb_desc_2_axsize_reg[2:0] = int_desc_2_axsize_axsize;
assign uc2rb_desc_2_axaddr_0_reg[31:0] = int_desc_2_axaddr_0_addr;
assign uc2rb_desc_2_axaddr_1_reg[31:0] = int_desc_2_axaddr_1_addr;
assign uc2rb_desc_2_axaddr_2_reg[31:0] = int_desc_2_axaddr_2_addr;
assign uc2rb_desc_2_axaddr_3_reg[31:0] = int_desc_2_axaddr_3_addr;
assign uc2rb_desc_2_data_offset_reg[31:0] = int_desc_2_data_offset_addr;
assign uc2rb_desc_2_wuser_0_reg[31:0] = int_desc_2_wuser_0_wuser;
assign uc2rb_desc_2_wuser_1_reg[31:0] = int_desc_2_wuser_1_wuser;
assign uc2rb_desc_2_wuser_2_reg[31:0] = int_desc_2_wuser_2_wuser;
assign uc2rb_desc_2_wuser_3_reg[31:0] = int_desc_2_wuser_3_wuser;
assign uc2rb_desc_2_wuser_4_reg[31:0] = int_desc_2_wuser_4_wuser;
assign uc2rb_desc_2_wuser_5_reg[31:0] = int_desc_2_wuser_5_wuser;
assign uc2rb_desc_2_wuser_6_reg[31:0] = int_desc_2_wuser_6_wuser;
assign uc2rb_desc_2_wuser_7_reg[31:0] = int_desc_2_wuser_7_wuser;
assign uc2rb_desc_2_wuser_8_reg[31:0] = int_desc_2_wuser_8_wuser;
assign uc2rb_desc_2_wuser_9_reg[31:0] = int_desc_2_wuser_9_wuser;
assign uc2rb_desc_2_wuser_10_reg[31:0] = int_desc_2_wuser_10_wuser;
assign uc2rb_desc_2_wuser_11_reg[31:0] = int_desc_2_wuser_11_wuser;
assign uc2rb_desc_2_wuser_12_reg[31:0] = int_desc_2_wuser_12_wuser;
assign uc2rb_desc_2_wuser_13_reg[31:0] = int_desc_2_wuser_13_wuser;
assign uc2rb_desc_2_wuser_14_reg[31:0] = int_desc_2_wuser_14_wuser;
assign uc2rb_desc_2_wuser_15_reg[31:0] = int_desc_2_wuser_15_wuser;
assign uc2rb_desc_3_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_3_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_3_size_reg[31:16] = 16'h0;
assign uc2rb_desc_3_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_3_txn_type_reg[1] = int_desc_3_txn_type_wr_strb;
assign uc2rb_desc_3_txn_type_reg[0] = int_desc_3_txn_type_wr_rd;
assign uc2rb_desc_3_attr_reg[18:15] = int_desc_3_attr_axregion;
assign uc2rb_desc_3_attr_reg[14:11] = int_desc_3_attr_axqos;
assign uc2rb_desc_3_attr_reg[10:8] = int_desc_3_attr_axprot;
assign uc2rb_desc_3_attr_reg[7:4] = int_desc_3_attr_axcache;
assign uc2rb_desc_3_attr_reg[3:2] = int_desc_3_attr_axlock;
assign uc2rb_desc_3_attr_reg[1:0] = int_desc_3_attr_axburst;
assign uc2rb_desc_3_axid_0_reg[31:0] = int_desc_3_axid_0_axid;
assign uc2rb_desc_3_axid_1_reg[31:0] = int_desc_3_axid_1_axid;
assign uc2rb_desc_3_axid_2_reg[31:0] = int_desc_3_axid_2_axid;
assign uc2rb_desc_3_axid_3_reg[31:0] = int_desc_3_axid_3_axid;
assign uc2rb_desc_3_axuser_0_reg[31:0] = int_desc_3_axuser_0_axuser;
assign uc2rb_desc_3_axuser_1_reg[31:0] = int_desc_3_axuser_1_axuser;
assign uc2rb_desc_3_axuser_2_reg[31:0] = int_desc_3_axuser_2_axuser;
assign uc2rb_desc_3_axuser_3_reg[31:0] = int_desc_3_axuser_3_axuser;
assign uc2rb_desc_3_axuser_4_reg[31:0] = int_desc_3_axuser_4_axuser;
assign uc2rb_desc_3_axuser_5_reg[31:0] = int_desc_3_axuser_5_axuser;
assign uc2rb_desc_3_axuser_6_reg[31:0] = int_desc_3_axuser_6_axuser;
assign uc2rb_desc_3_axuser_7_reg[31:0] = int_desc_3_axuser_7_axuser;
assign uc2rb_desc_3_axuser_8_reg[31:0] = int_desc_3_axuser_8_axuser;
assign uc2rb_desc_3_axuser_9_reg[31:0] = int_desc_3_axuser_9_axuser;
assign uc2rb_desc_3_axuser_10_reg[31:0] = int_desc_3_axuser_10_axuser;
assign uc2rb_desc_3_axuser_11_reg[31:0] = int_desc_3_axuser_11_axuser;
assign uc2rb_desc_3_axuser_12_reg[31:0] = int_desc_3_axuser_12_axuser;
assign uc2rb_desc_3_axuser_13_reg[31:0] = int_desc_3_axuser_13_axuser;
assign uc2rb_desc_3_axuser_14_reg[31:0] = int_desc_3_axuser_14_axuser;
assign uc2rb_desc_3_axuser_15_reg[31:0] = int_desc_3_axuser_15_axuser;
assign uc2rb_desc_3_size_reg[15:0] = int_desc_3_size_txn_size;
assign uc2rb_desc_3_axsize_reg[2:0] = int_desc_3_axsize_axsize;
assign uc2rb_desc_3_axaddr_0_reg[31:0] = int_desc_3_axaddr_0_addr;
assign uc2rb_desc_3_axaddr_1_reg[31:0] = int_desc_3_axaddr_1_addr;
assign uc2rb_desc_3_axaddr_2_reg[31:0] = int_desc_3_axaddr_2_addr;
assign uc2rb_desc_3_axaddr_3_reg[31:0] = int_desc_3_axaddr_3_addr;
assign uc2rb_desc_3_data_offset_reg[31:0] = int_desc_3_data_offset_addr;
assign uc2rb_desc_3_wuser_0_reg[31:0] = int_desc_3_wuser_0_wuser;
assign uc2rb_desc_3_wuser_1_reg[31:0] = int_desc_3_wuser_1_wuser;
assign uc2rb_desc_3_wuser_2_reg[31:0] = int_desc_3_wuser_2_wuser;
assign uc2rb_desc_3_wuser_3_reg[31:0] = int_desc_3_wuser_3_wuser;
assign uc2rb_desc_3_wuser_4_reg[31:0] = int_desc_3_wuser_4_wuser;
assign uc2rb_desc_3_wuser_5_reg[31:0] = int_desc_3_wuser_5_wuser;
assign uc2rb_desc_3_wuser_6_reg[31:0] = int_desc_3_wuser_6_wuser;
assign uc2rb_desc_3_wuser_7_reg[31:0] = int_desc_3_wuser_7_wuser;
assign uc2rb_desc_3_wuser_8_reg[31:0] = int_desc_3_wuser_8_wuser;
assign uc2rb_desc_3_wuser_9_reg[31:0] = int_desc_3_wuser_9_wuser;
assign uc2rb_desc_3_wuser_10_reg[31:0] = int_desc_3_wuser_10_wuser;
assign uc2rb_desc_3_wuser_11_reg[31:0] = int_desc_3_wuser_11_wuser;
assign uc2rb_desc_3_wuser_12_reg[31:0] = int_desc_3_wuser_12_wuser;
assign uc2rb_desc_3_wuser_13_reg[31:0] = int_desc_3_wuser_13_wuser;
assign uc2rb_desc_3_wuser_14_reg[31:0] = int_desc_3_wuser_14_wuser;
assign uc2rb_desc_3_wuser_15_reg[31:0] = int_desc_3_wuser_15_wuser;
assign uc2rb_desc_4_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_4_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_4_size_reg[31:16] = 16'h0;
assign uc2rb_desc_4_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_4_txn_type_reg[1] = int_desc_4_txn_type_wr_strb;
assign uc2rb_desc_4_txn_type_reg[0] = int_desc_4_txn_type_wr_rd;
assign uc2rb_desc_4_attr_reg[18:15] = int_desc_4_attr_axregion;
assign uc2rb_desc_4_attr_reg[14:11] = int_desc_4_attr_axqos;
assign uc2rb_desc_4_attr_reg[10:8] = int_desc_4_attr_axprot;
assign uc2rb_desc_4_attr_reg[7:4] = int_desc_4_attr_axcache;
assign uc2rb_desc_4_attr_reg[3:2] = int_desc_4_attr_axlock;
assign uc2rb_desc_4_attr_reg[1:0] = int_desc_4_attr_axburst;
assign uc2rb_desc_4_axid_0_reg[31:0] = int_desc_4_axid_0_axid;
assign uc2rb_desc_4_axid_1_reg[31:0] = int_desc_4_axid_1_axid;
assign uc2rb_desc_4_axid_2_reg[31:0] = int_desc_4_axid_2_axid;
assign uc2rb_desc_4_axid_3_reg[31:0] = int_desc_4_axid_3_axid;
assign uc2rb_desc_4_axuser_0_reg[31:0] = int_desc_4_axuser_0_axuser;
assign uc2rb_desc_4_axuser_1_reg[31:0] = int_desc_4_axuser_1_axuser;
assign uc2rb_desc_4_axuser_2_reg[31:0] = int_desc_4_axuser_2_axuser;
assign uc2rb_desc_4_axuser_3_reg[31:0] = int_desc_4_axuser_3_axuser;
assign uc2rb_desc_4_axuser_4_reg[31:0] = int_desc_4_axuser_4_axuser;
assign uc2rb_desc_4_axuser_5_reg[31:0] = int_desc_4_axuser_5_axuser;
assign uc2rb_desc_4_axuser_6_reg[31:0] = int_desc_4_axuser_6_axuser;
assign uc2rb_desc_4_axuser_7_reg[31:0] = int_desc_4_axuser_7_axuser;
assign uc2rb_desc_4_axuser_8_reg[31:0] = int_desc_4_axuser_8_axuser;
assign uc2rb_desc_4_axuser_9_reg[31:0] = int_desc_4_axuser_9_axuser;
assign uc2rb_desc_4_axuser_10_reg[31:0] = int_desc_4_axuser_10_axuser;
assign uc2rb_desc_4_axuser_11_reg[31:0] = int_desc_4_axuser_11_axuser;
assign uc2rb_desc_4_axuser_12_reg[31:0] = int_desc_4_axuser_12_axuser;
assign uc2rb_desc_4_axuser_13_reg[31:0] = int_desc_4_axuser_13_axuser;
assign uc2rb_desc_4_axuser_14_reg[31:0] = int_desc_4_axuser_14_axuser;
assign uc2rb_desc_4_axuser_15_reg[31:0] = int_desc_4_axuser_15_axuser;
assign uc2rb_desc_4_size_reg[15:0] = int_desc_4_size_txn_size;
assign uc2rb_desc_4_axsize_reg[2:0] = int_desc_4_axsize_axsize;
assign uc2rb_desc_4_axaddr_0_reg[31:0] = int_desc_4_axaddr_0_addr;
assign uc2rb_desc_4_axaddr_1_reg[31:0] = int_desc_4_axaddr_1_addr;
assign uc2rb_desc_4_axaddr_2_reg[31:0] = int_desc_4_axaddr_2_addr;
assign uc2rb_desc_4_axaddr_3_reg[31:0] = int_desc_4_axaddr_3_addr;
assign uc2rb_desc_4_data_offset_reg[31:0] = int_desc_4_data_offset_addr;
assign uc2rb_desc_4_wuser_0_reg[31:0] = int_desc_4_wuser_0_wuser;
assign uc2rb_desc_4_wuser_1_reg[31:0] = int_desc_4_wuser_1_wuser;
assign uc2rb_desc_4_wuser_2_reg[31:0] = int_desc_4_wuser_2_wuser;
assign uc2rb_desc_4_wuser_3_reg[31:0] = int_desc_4_wuser_3_wuser;
assign uc2rb_desc_4_wuser_4_reg[31:0] = int_desc_4_wuser_4_wuser;
assign uc2rb_desc_4_wuser_5_reg[31:0] = int_desc_4_wuser_5_wuser;
assign uc2rb_desc_4_wuser_6_reg[31:0] = int_desc_4_wuser_6_wuser;
assign uc2rb_desc_4_wuser_7_reg[31:0] = int_desc_4_wuser_7_wuser;
assign uc2rb_desc_4_wuser_8_reg[31:0] = int_desc_4_wuser_8_wuser;
assign uc2rb_desc_4_wuser_9_reg[31:0] = int_desc_4_wuser_9_wuser;
assign uc2rb_desc_4_wuser_10_reg[31:0] = int_desc_4_wuser_10_wuser;
assign uc2rb_desc_4_wuser_11_reg[31:0] = int_desc_4_wuser_11_wuser;
assign uc2rb_desc_4_wuser_12_reg[31:0] = int_desc_4_wuser_12_wuser;
assign uc2rb_desc_4_wuser_13_reg[31:0] = int_desc_4_wuser_13_wuser;
assign uc2rb_desc_4_wuser_14_reg[31:0] = int_desc_4_wuser_14_wuser;
assign uc2rb_desc_4_wuser_15_reg[31:0] = int_desc_4_wuser_15_wuser;
assign uc2rb_desc_5_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_5_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_5_size_reg[31:16] = 16'h0;
assign uc2rb_desc_5_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_5_txn_type_reg[1] = int_desc_5_txn_type_wr_strb;
assign uc2rb_desc_5_txn_type_reg[0] = int_desc_5_txn_type_wr_rd;
assign uc2rb_desc_5_attr_reg[18:15] = int_desc_5_attr_axregion;
assign uc2rb_desc_5_attr_reg[14:11] = int_desc_5_attr_axqos;
assign uc2rb_desc_5_attr_reg[10:8] = int_desc_5_attr_axprot;
assign uc2rb_desc_5_attr_reg[7:4] = int_desc_5_attr_axcache;
assign uc2rb_desc_5_attr_reg[3:2] = int_desc_5_attr_axlock;
assign uc2rb_desc_5_attr_reg[1:0] = int_desc_5_attr_axburst;
assign uc2rb_desc_5_axid_0_reg[31:0] = int_desc_5_axid_0_axid;
assign uc2rb_desc_5_axid_1_reg[31:0] = int_desc_5_axid_1_axid;
assign uc2rb_desc_5_axid_2_reg[31:0] = int_desc_5_axid_2_axid;
assign uc2rb_desc_5_axid_3_reg[31:0] = int_desc_5_axid_3_axid;
assign uc2rb_desc_5_axuser_0_reg[31:0] = int_desc_5_axuser_0_axuser;
assign uc2rb_desc_5_axuser_1_reg[31:0] = int_desc_5_axuser_1_axuser;
assign uc2rb_desc_5_axuser_2_reg[31:0] = int_desc_5_axuser_2_axuser;
assign uc2rb_desc_5_axuser_3_reg[31:0] = int_desc_5_axuser_3_axuser;
assign uc2rb_desc_5_axuser_4_reg[31:0] = int_desc_5_axuser_4_axuser;
assign uc2rb_desc_5_axuser_5_reg[31:0] = int_desc_5_axuser_5_axuser;
assign uc2rb_desc_5_axuser_6_reg[31:0] = int_desc_5_axuser_6_axuser;
assign uc2rb_desc_5_axuser_7_reg[31:0] = int_desc_5_axuser_7_axuser;
assign uc2rb_desc_5_axuser_8_reg[31:0] = int_desc_5_axuser_8_axuser;
assign uc2rb_desc_5_axuser_9_reg[31:0] = int_desc_5_axuser_9_axuser;
assign uc2rb_desc_5_axuser_10_reg[31:0] = int_desc_5_axuser_10_axuser;
assign uc2rb_desc_5_axuser_11_reg[31:0] = int_desc_5_axuser_11_axuser;
assign uc2rb_desc_5_axuser_12_reg[31:0] = int_desc_5_axuser_12_axuser;
assign uc2rb_desc_5_axuser_13_reg[31:0] = int_desc_5_axuser_13_axuser;
assign uc2rb_desc_5_axuser_14_reg[31:0] = int_desc_5_axuser_14_axuser;
assign uc2rb_desc_5_axuser_15_reg[31:0] = int_desc_5_axuser_15_axuser;
assign uc2rb_desc_5_size_reg[15:0] = int_desc_5_size_txn_size;
assign uc2rb_desc_5_axsize_reg[2:0] = int_desc_5_axsize_axsize;
assign uc2rb_desc_5_axaddr_0_reg[31:0] = int_desc_5_axaddr_0_addr;
assign uc2rb_desc_5_axaddr_1_reg[31:0] = int_desc_5_axaddr_1_addr;
assign uc2rb_desc_5_axaddr_2_reg[31:0] = int_desc_5_axaddr_2_addr;
assign uc2rb_desc_5_axaddr_3_reg[31:0] = int_desc_5_axaddr_3_addr;
assign uc2rb_desc_5_data_offset_reg[31:0] = int_desc_5_data_offset_addr;
assign uc2rb_desc_5_wuser_0_reg[31:0] = int_desc_5_wuser_0_wuser;
assign uc2rb_desc_5_wuser_1_reg[31:0] = int_desc_5_wuser_1_wuser;
assign uc2rb_desc_5_wuser_2_reg[31:0] = int_desc_5_wuser_2_wuser;
assign uc2rb_desc_5_wuser_3_reg[31:0] = int_desc_5_wuser_3_wuser;
assign uc2rb_desc_5_wuser_4_reg[31:0] = int_desc_5_wuser_4_wuser;
assign uc2rb_desc_5_wuser_5_reg[31:0] = int_desc_5_wuser_5_wuser;
assign uc2rb_desc_5_wuser_6_reg[31:0] = int_desc_5_wuser_6_wuser;
assign uc2rb_desc_5_wuser_7_reg[31:0] = int_desc_5_wuser_7_wuser;
assign uc2rb_desc_5_wuser_8_reg[31:0] = int_desc_5_wuser_8_wuser;
assign uc2rb_desc_5_wuser_9_reg[31:0] = int_desc_5_wuser_9_wuser;
assign uc2rb_desc_5_wuser_10_reg[31:0] = int_desc_5_wuser_10_wuser;
assign uc2rb_desc_5_wuser_11_reg[31:0] = int_desc_5_wuser_11_wuser;
assign uc2rb_desc_5_wuser_12_reg[31:0] = int_desc_5_wuser_12_wuser;
assign uc2rb_desc_5_wuser_13_reg[31:0] = int_desc_5_wuser_13_wuser;
assign uc2rb_desc_5_wuser_14_reg[31:0] = int_desc_5_wuser_14_wuser;
assign uc2rb_desc_5_wuser_15_reg[31:0] = int_desc_5_wuser_15_wuser;
assign uc2rb_desc_6_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_6_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_6_size_reg[31:16] = 16'h0;
assign uc2rb_desc_6_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_6_txn_type_reg[1] = int_desc_6_txn_type_wr_strb;
assign uc2rb_desc_6_txn_type_reg[0] = int_desc_6_txn_type_wr_rd;
assign uc2rb_desc_6_attr_reg[18:15] = int_desc_6_attr_axregion;
assign uc2rb_desc_6_attr_reg[14:11] = int_desc_6_attr_axqos;
assign uc2rb_desc_6_attr_reg[10:8] = int_desc_6_attr_axprot;
assign uc2rb_desc_6_attr_reg[7:4] = int_desc_6_attr_axcache;
assign uc2rb_desc_6_attr_reg[3:2] = int_desc_6_attr_axlock;
assign uc2rb_desc_6_attr_reg[1:0] = int_desc_6_attr_axburst;
assign uc2rb_desc_6_axid_0_reg[31:0] = int_desc_6_axid_0_axid;
assign uc2rb_desc_6_axid_1_reg[31:0] = int_desc_6_axid_1_axid;
assign uc2rb_desc_6_axid_2_reg[31:0] = int_desc_6_axid_2_axid;
assign uc2rb_desc_6_axid_3_reg[31:0] = int_desc_6_axid_3_axid;
assign uc2rb_desc_6_axuser_0_reg[31:0] = int_desc_6_axuser_0_axuser;
assign uc2rb_desc_6_axuser_1_reg[31:0] = int_desc_6_axuser_1_axuser;
assign uc2rb_desc_6_axuser_2_reg[31:0] = int_desc_6_axuser_2_axuser;
assign uc2rb_desc_6_axuser_3_reg[31:0] = int_desc_6_axuser_3_axuser;
assign uc2rb_desc_6_axuser_4_reg[31:0] = int_desc_6_axuser_4_axuser;
assign uc2rb_desc_6_axuser_5_reg[31:0] = int_desc_6_axuser_5_axuser;
assign uc2rb_desc_6_axuser_6_reg[31:0] = int_desc_6_axuser_6_axuser;
assign uc2rb_desc_6_axuser_7_reg[31:0] = int_desc_6_axuser_7_axuser;
assign uc2rb_desc_6_axuser_8_reg[31:0] = int_desc_6_axuser_8_axuser;
assign uc2rb_desc_6_axuser_9_reg[31:0] = int_desc_6_axuser_9_axuser;
assign uc2rb_desc_6_axuser_10_reg[31:0] = int_desc_6_axuser_10_axuser;
assign uc2rb_desc_6_axuser_11_reg[31:0] = int_desc_6_axuser_11_axuser;
assign uc2rb_desc_6_axuser_12_reg[31:0] = int_desc_6_axuser_12_axuser;
assign uc2rb_desc_6_axuser_13_reg[31:0] = int_desc_6_axuser_13_axuser;
assign uc2rb_desc_6_axuser_14_reg[31:0] = int_desc_6_axuser_14_axuser;
assign uc2rb_desc_6_axuser_15_reg[31:0] = int_desc_6_axuser_15_axuser;
assign uc2rb_desc_6_size_reg[15:0] = int_desc_6_size_txn_size;
assign uc2rb_desc_6_axsize_reg[2:0] = int_desc_6_axsize_axsize;
assign uc2rb_desc_6_axaddr_0_reg[31:0] = int_desc_6_axaddr_0_addr;
assign uc2rb_desc_6_axaddr_1_reg[31:0] = int_desc_6_axaddr_1_addr;
assign uc2rb_desc_6_axaddr_2_reg[31:0] = int_desc_6_axaddr_2_addr;
assign uc2rb_desc_6_axaddr_3_reg[31:0] = int_desc_6_axaddr_3_addr;
assign uc2rb_desc_6_data_offset_reg[31:0] = int_desc_6_data_offset_addr;
assign uc2rb_desc_6_wuser_0_reg[31:0] = int_desc_6_wuser_0_wuser;
assign uc2rb_desc_6_wuser_1_reg[31:0] = int_desc_6_wuser_1_wuser;
assign uc2rb_desc_6_wuser_2_reg[31:0] = int_desc_6_wuser_2_wuser;
assign uc2rb_desc_6_wuser_3_reg[31:0] = int_desc_6_wuser_3_wuser;
assign uc2rb_desc_6_wuser_4_reg[31:0] = int_desc_6_wuser_4_wuser;
assign uc2rb_desc_6_wuser_5_reg[31:0] = int_desc_6_wuser_5_wuser;
assign uc2rb_desc_6_wuser_6_reg[31:0] = int_desc_6_wuser_6_wuser;
assign uc2rb_desc_6_wuser_7_reg[31:0] = int_desc_6_wuser_7_wuser;
assign uc2rb_desc_6_wuser_8_reg[31:0] = int_desc_6_wuser_8_wuser;
assign uc2rb_desc_6_wuser_9_reg[31:0] = int_desc_6_wuser_9_wuser;
assign uc2rb_desc_6_wuser_10_reg[31:0] = int_desc_6_wuser_10_wuser;
assign uc2rb_desc_6_wuser_11_reg[31:0] = int_desc_6_wuser_11_wuser;
assign uc2rb_desc_6_wuser_12_reg[31:0] = int_desc_6_wuser_12_wuser;
assign uc2rb_desc_6_wuser_13_reg[31:0] = int_desc_6_wuser_13_wuser;
assign uc2rb_desc_6_wuser_14_reg[31:0] = int_desc_6_wuser_14_wuser;
assign uc2rb_desc_6_wuser_15_reg[31:0] = int_desc_6_wuser_15_wuser;
assign uc2rb_desc_7_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_7_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_7_size_reg[31:16] = 16'h0;
assign uc2rb_desc_7_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_7_txn_type_reg[1] = int_desc_7_txn_type_wr_strb;
assign uc2rb_desc_7_txn_type_reg[0] = int_desc_7_txn_type_wr_rd;
assign uc2rb_desc_7_attr_reg[18:15] = int_desc_7_attr_axregion;
assign uc2rb_desc_7_attr_reg[14:11] = int_desc_7_attr_axqos;
assign uc2rb_desc_7_attr_reg[10:8] = int_desc_7_attr_axprot;
assign uc2rb_desc_7_attr_reg[7:4] = int_desc_7_attr_axcache;
assign uc2rb_desc_7_attr_reg[3:2] = int_desc_7_attr_axlock;
assign uc2rb_desc_7_attr_reg[1:0] = int_desc_7_attr_axburst;
assign uc2rb_desc_7_axid_0_reg[31:0] = int_desc_7_axid_0_axid;
assign uc2rb_desc_7_axid_1_reg[31:0] = int_desc_7_axid_1_axid;
assign uc2rb_desc_7_axid_2_reg[31:0] = int_desc_7_axid_2_axid;
assign uc2rb_desc_7_axid_3_reg[31:0] = int_desc_7_axid_3_axid;
assign uc2rb_desc_7_axuser_0_reg[31:0] = int_desc_7_axuser_0_axuser;
assign uc2rb_desc_7_axuser_1_reg[31:0] = int_desc_7_axuser_1_axuser;
assign uc2rb_desc_7_axuser_2_reg[31:0] = int_desc_7_axuser_2_axuser;
assign uc2rb_desc_7_axuser_3_reg[31:0] = int_desc_7_axuser_3_axuser;
assign uc2rb_desc_7_axuser_4_reg[31:0] = int_desc_7_axuser_4_axuser;
assign uc2rb_desc_7_axuser_5_reg[31:0] = int_desc_7_axuser_5_axuser;
assign uc2rb_desc_7_axuser_6_reg[31:0] = int_desc_7_axuser_6_axuser;
assign uc2rb_desc_7_axuser_7_reg[31:0] = int_desc_7_axuser_7_axuser;
assign uc2rb_desc_7_axuser_8_reg[31:0] = int_desc_7_axuser_8_axuser;
assign uc2rb_desc_7_axuser_9_reg[31:0] = int_desc_7_axuser_9_axuser;
assign uc2rb_desc_7_axuser_10_reg[31:0] = int_desc_7_axuser_10_axuser;
assign uc2rb_desc_7_axuser_11_reg[31:0] = int_desc_7_axuser_11_axuser;
assign uc2rb_desc_7_axuser_12_reg[31:0] = int_desc_7_axuser_12_axuser;
assign uc2rb_desc_7_axuser_13_reg[31:0] = int_desc_7_axuser_13_axuser;
assign uc2rb_desc_7_axuser_14_reg[31:0] = int_desc_7_axuser_14_axuser;
assign uc2rb_desc_7_axuser_15_reg[31:0] = int_desc_7_axuser_15_axuser;
assign uc2rb_desc_7_size_reg[15:0] = int_desc_7_size_txn_size;
assign uc2rb_desc_7_axsize_reg[2:0] = int_desc_7_axsize_axsize;
assign uc2rb_desc_7_axaddr_0_reg[31:0] = int_desc_7_axaddr_0_addr;
assign uc2rb_desc_7_axaddr_1_reg[31:0] = int_desc_7_axaddr_1_addr;
assign uc2rb_desc_7_axaddr_2_reg[31:0] = int_desc_7_axaddr_2_addr;
assign uc2rb_desc_7_axaddr_3_reg[31:0] = int_desc_7_axaddr_3_addr;
assign uc2rb_desc_7_data_offset_reg[31:0] = int_desc_7_data_offset_addr;
assign uc2rb_desc_7_wuser_0_reg[31:0] = int_desc_7_wuser_0_wuser;
assign uc2rb_desc_7_wuser_1_reg[31:0] = int_desc_7_wuser_1_wuser;
assign uc2rb_desc_7_wuser_2_reg[31:0] = int_desc_7_wuser_2_wuser;
assign uc2rb_desc_7_wuser_3_reg[31:0] = int_desc_7_wuser_3_wuser;
assign uc2rb_desc_7_wuser_4_reg[31:0] = int_desc_7_wuser_4_wuser;
assign uc2rb_desc_7_wuser_5_reg[31:0] = int_desc_7_wuser_5_wuser;
assign uc2rb_desc_7_wuser_6_reg[31:0] = int_desc_7_wuser_6_wuser;
assign uc2rb_desc_7_wuser_7_reg[31:0] = int_desc_7_wuser_7_wuser;
assign uc2rb_desc_7_wuser_8_reg[31:0] = int_desc_7_wuser_8_wuser;
assign uc2rb_desc_7_wuser_9_reg[31:0] = int_desc_7_wuser_9_wuser;
assign uc2rb_desc_7_wuser_10_reg[31:0] = int_desc_7_wuser_10_wuser;
assign uc2rb_desc_7_wuser_11_reg[31:0] = int_desc_7_wuser_11_wuser;
assign uc2rb_desc_7_wuser_12_reg[31:0] = int_desc_7_wuser_12_wuser;
assign uc2rb_desc_7_wuser_13_reg[31:0] = int_desc_7_wuser_13_wuser;
assign uc2rb_desc_7_wuser_14_reg[31:0] = int_desc_7_wuser_14_wuser;
assign uc2rb_desc_7_wuser_15_reg[31:0] = int_desc_7_wuser_15_wuser;
assign uc2rb_desc_8_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_8_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_8_size_reg[31:16] = 16'h0;
assign uc2rb_desc_8_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_8_txn_type_reg[1] = int_desc_8_txn_type_wr_strb;
assign uc2rb_desc_8_txn_type_reg[0] = int_desc_8_txn_type_wr_rd;
assign uc2rb_desc_8_attr_reg[18:15] = int_desc_8_attr_axregion;
assign uc2rb_desc_8_attr_reg[14:11] = int_desc_8_attr_axqos;
assign uc2rb_desc_8_attr_reg[10:8] = int_desc_8_attr_axprot;
assign uc2rb_desc_8_attr_reg[7:4] = int_desc_8_attr_axcache;
assign uc2rb_desc_8_attr_reg[3:2] = int_desc_8_attr_axlock;
assign uc2rb_desc_8_attr_reg[1:0] = int_desc_8_attr_axburst;
assign uc2rb_desc_8_axid_0_reg[31:0] = int_desc_8_axid_0_axid;
assign uc2rb_desc_8_axid_1_reg[31:0] = int_desc_8_axid_1_axid;
assign uc2rb_desc_8_axid_2_reg[31:0] = int_desc_8_axid_2_axid;
assign uc2rb_desc_8_axid_3_reg[31:0] = int_desc_8_axid_3_axid;
assign uc2rb_desc_8_axuser_0_reg[31:0] = int_desc_8_axuser_0_axuser;
assign uc2rb_desc_8_axuser_1_reg[31:0] = int_desc_8_axuser_1_axuser;
assign uc2rb_desc_8_axuser_2_reg[31:0] = int_desc_8_axuser_2_axuser;
assign uc2rb_desc_8_axuser_3_reg[31:0] = int_desc_8_axuser_3_axuser;
assign uc2rb_desc_8_axuser_4_reg[31:0] = int_desc_8_axuser_4_axuser;
assign uc2rb_desc_8_axuser_5_reg[31:0] = int_desc_8_axuser_5_axuser;
assign uc2rb_desc_8_axuser_6_reg[31:0] = int_desc_8_axuser_6_axuser;
assign uc2rb_desc_8_axuser_7_reg[31:0] = int_desc_8_axuser_7_axuser;
assign uc2rb_desc_8_axuser_8_reg[31:0] = int_desc_8_axuser_8_axuser;
assign uc2rb_desc_8_axuser_9_reg[31:0] = int_desc_8_axuser_9_axuser;
assign uc2rb_desc_8_axuser_10_reg[31:0] = int_desc_8_axuser_10_axuser;
assign uc2rb_desc_8_axuser_11_reg[31:0] = int_desc_8_axuser_11_axuser;
assign uc2rb_desc_8_axuser_12_reg[31:0] = int_desc_8_axuser_12_axuser;
assign uc2rb_desc_8_axuser_13_reg[31:0] = int_desc_8_axuser_13_axuser;
assign uc2rb_desc_8_axuser_14_reg[31:0] = int_desc_8_axuser_14_axuser;
assign uc2rb_desc_8_axuser_15_reg[31:0] = int_desc_8_axuser_15_axuser;
assign uc2rb_desc_8_size_reg[15:0] = int_desc_8_size_txn_size;
assign uc2rb_desc_8_axsize_reg[2:0] = int_desc_8_axsize_axsize;
assign uc2rb_desc_8_axaddr_0_reg[31:0] = int_desc_8_axaddr_0_addr;
assign uc2rb_desc_8_axaddr_1_reg[31:0] = int_desc_8_axaddr_1_addr;
assign uc2rb_desc_8_axaddr_2_reg[31:0] = int_desc_8_axaddr_2_addr;
assign uc2rb_desc_8_axaddr_3_reg[31:0] = int_desc_8_axaddr_3_addr;
assign uc2rb_desc_8_data_offset_reg[31:0] = int_desc_8_data_offset_addr;
assign uc2rb_desc_8_wuser_0_reg[31:0] = int_desc_8_wuser_0_wuser;
assign uc2rb_desc_8_wuser_1_reg[31:0] = int_desc_8_wuser_1_wuser;
assign uc2rb_desc_8_wuser_2_reg[31:0] = int_desc_8_wuser_2_wuser;
assign uc2rb_desc_8_wuser_3_reg[31:0] = int_desc_8_wuser_3_wuser;
assign uc2rb_desc_8_wuser_4_reg[31:0] = int_desc_8_wuser_4_wuser;
assign uc2rb_desc_8_wuser_5_reg[31:0] = int_desc_8_wuser_5_wuser;
assign uc2rb_desc_8_wuser_6_reg[31:0] = int_desc_8_wuser_6_wuser;
assign uc2rb_desc_8_wuser_7_reg[31:0] = int_desc_8_wuser_7_wuser;
assign uc2rb_desc_8_wuser_8_reg[31:0] = int_desc_8_wuser_8_wuser;
assign uc2rb_desc_8_wuser_9_reg[31:0] = int_desc_8_wuser_9_wuser;
assign uc2rb_desc_8_wuser_10_reg[31:0] = int_desc_8_wuser_10_wuser;
assign uc2rb_desc_8_wuser_11_reg[31:0] = int_desc_8_wuser_11_wuser;
assign uc2rb_desc_8_wuser_12_reg[31:0] = int_desc_8_wuser_12_wuser;
assign uc2rb_desc_8_wuser_13_reg[31:0] = int_desc_8_wuser_13_wuser;
assign uc2rb_desc_8_wuser_14_reg[31:0] = int_desc_8_wuser_14_wuser;
assign uc2rb_desc_8_wuser_15_reg[31:0] = int_desc_8_wuser_15_wuser;
assign uc2rb_desc_9_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_9_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_9_size_reg[31:16] = 16'h0;
assign uc2rb_desc_9_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_9_txn_type_reg[1] = int_desc_9_txn_type_wr_strb;
assign uc2rb_desc_9_txn_type_reg[0] = int_desc_9_txn_type_wr_rd;
assign uc2rb_desc_9_attr_reg[18:15] = int_desc_9_attr_axregion;
assign uc2rb_desc_9_attr_reg[14:11] = int_desc_9_attr_axqos;
assign uc2rb_desc_9_attr_reg[10:8] = int_desc_9_attr_axprot;
assign uc2rb_desc_9_attr_reg[7:4] = int_desc_9_attr_axcache;
assign uc2rb_desc_9_attr_reg[3:2] = int_desc_9_attr_axlock;
assign uc2rb_desc_9_attr_reg[1:0] = int_desc_9_attr_axburst;
assign uc2rb_desc_9_axid_0_reg[31:0] = int_desc_9_axid_0_axid;
assign uc2rb_desc_9_axid_1_reg[31:0] = int_desc_9_axid_1_axid;
assign uc2rb_desc_9_axid_2_reg[31:0] = int_desc_9_axid_2_axid;
assign uc2rb_desc_9_axid_3_reg[31:0] = int_desc_9_axid_3_axid;
assign uc2rb_desc_9_axuser_0_reg[31:0] = int_desc_9_axuser_0_axuser;
assign uc2rb_desc_9_axuser_1_reg[31:0] = int_desc_9_axuser_1_axuser;
assign uc2rb_desc_9_axuser_2_reg[31:0] = int_desc_9_axuser_2_axuser;
assign uc2rb_desc_9_axuser_3_reg[31:0] = int_desc_9_axuser_3_axuser;
assign uc2rb_desc_9_axuser_4_reg[31:0] = int_desc_9_axuser_4_axuser;
assign uc2rb_desc_9_axuser_5_reg[31:0] = int_desc_9_axuser_5_axuser;
assign uc2rb_desc_9_axuser_6_reg[31:0] = int_desc_9_axuser_6_axuser;
assign uc2rb_desc_9_axuser_7_reg[31:0] = int_desc_9_axuser_7_axuser;
assign uc2rb_desc_9_axuser_8_reg[31:0] = int_desc_9_axuser_8_axuser;
assign uc2rb_desc_9_axuser_9_reg[31:0] = int_desc_9_axuser_9_axuser;
assign uc2rb_desc_9_axuser_10_reg[31:0] = int_desc_9_axuser_10_axuser;
assign uc2rb_desc_9_axuser_11_reg[31:0] = int_desc_9_axuser_11_axuser;
assign uc2rb_desc_9_axuser_12_reg[31:0] = int_desc_9_axuser_12_axuser;
assign uc2rb_desc_9_axuser_13_reg[31:0] = int_desc_9_axuser_13_axuser;
assign uc2rb_desc_9_axuser_14_reg[31:0] = int_desc_9_axuser_14_axuser;
assign uc2rb_desc_9_axuser_15_reg[31:0] = int_desc_9_axuser_15_axuser;
assign uc2rb_desc_9_size_reg[15:0] = int_desc_9_size_txn_size;
assign uc2rb_desc_9_axsize_reg[2:0] = int_desc_9_axsize_axsize;
assign uc2rb_desc_9_axaddr_0_reg[31:0] = int_desc_9_axaddr_0_addr;
assign uc2rb_desc_9_axaddr_1_reg[31:0] = int_desc_9_axaddr_1_addr;
assign uc2rb_desc_9_axaddr_2_reg[31:0] = int_desc_9_axaddr_2_addr;
assign uc2rb_desc_9_axaddr_3_reg[31:0] = int_desc_9_axaddr_3_addr;
assign uc2rb_desc_9_data_offset_reg[31:0] = int_desc_9_data_offset_addr;
assign uc2rb_desc_9_wuser_0_reg[31:0] = int_desc_9_wuser_0_wuser;
assign uc2rb_desc_9_wuser_1_reg[31:0] = int_desc_9_wuser_1_wuser;
assign uc2rb_desc_9_wuser_2_reg[31:0] = int_desc_9_wuser_2_wuser;
assign uc2rb_desc_9_wuser_3_reg[31:0] = int_desc_9_wuser_3_wuser;
assign uc2rb_desc_9_wuser_4_reg[31:0] = int_desc_9_wuser_4_wuser;
assign uc2rb_desc_9_wuser_5_reg[31:0] = int_desc_9_wuser_5_wuser;
assign uc2rb_desc_9_wuser_6_reg[31:0] = int_desc_9_wuser_6_wuser;
assign uc2rb_desc_9_wuser_7_reg[31:0] = int_desc_9_wuser_7_wuser;
assign uc2rb_desc_9_wuser_8_reg[31:0] = int_desc_9_wuser_8_wuser;
assign uc2rb_desc_9_wuser_9_reg[31:0] = int_desc_9_wuser_9_wuser;
assign uc2rb_desc_9_wuser_10_reg[31:0] = int_desc_9_wuser_10_wuser;
assign uc2rb_desc_9_wuser_11_reg[31:0] = int_desc_9_wuser_11_wuser;
assign uc2rb_desc_9_wuser_12_reg[31:0] = int_desc_9_wuser_12_wuser;
assign uc2rb_desc_9_wuser_13_reg[31:0] = int_desc_9_wuser_13_wuser;
assign uc2rb_desc_9_wuser_14_reg[31:0] = int_desc_9_wuser_14_wuser;
assign uc2rb_desc_9_wuser_15_reg[31:0] = int_desc_9_wuser_15_wuser;
assign uc2rb_desc_10_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_10_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_10_size_reg[31:16] = 16'h0;
assign uc2rb_desc_10_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_10_txn_type_reg[1] = int_desc_10_txn_type_wr_strb;
assign uc2rb_desc_10_txn_type_reg[0] = int_desc_10_txn_type_wr_rd;
assign uc2rb_desc_10_attr_reg[18:15] = int_desc_10_attr_axregion;
assign uc2rb_desc_10_attr_reg[14:11] = int_desc_10_attr_axqos;
assign uc2rb_desc_10_attr_reg[10:8] = int_desc_10_attr_axprot;
assign uc2rb_desc_10_attr_reg[7:4] = int_desc_10_attr_axcache;
assign uc2rb_desc_10_attr_reg[3:2] = int_desc_10_attr_axlock;
assign uc2rb_desc_10_attr_reg[1:0] = int_desc_10_attr_axburst;
assign uc2rb_desc_10_axid_0_reg[31:0] = int_desc_10_axid_0_axid;
assign uc2rb_desc_10_axid_1_reg[31:0] = int_desc_10_axid_1_axid;
assign uc2rb_desc_10_axid_2_reg[31:0] = int_desc_10_axid_2_axid;
assign uc2rb_desc_10_axid_3_reg[31:0] = int_desc_10_axid_3_axid;
assign uc2rb_desc_10_axuser_0_reg[31:0] = int_desc_10_axuser_0_axuser;
assign uc2rb_desc_10_axuser_1_reg[31:0] = int_desc_10_axuser_1_axuser;
assign uc2rb_desc_10_axuser_2_reg[31:0] = int_desc_10_axuser_2_axuser;
assign uc2rb_desc_10_axuser_3_reg[31:0] = int_desc_10_axuser_3_axuser;
assign uc2rb_desc_10_axuser_4_reg[31:0] = int_desc_10_axuser_4_axuser;
assign uc2rb_desc_10_axuser_5_reg[31:0] = int_desc_10_axuser_5_axuser;
assign uc2rb_desc_10_axuser_6_reg[31:0] = int_desc_10_axuser_6_axuser;
assign uc2rb_desc_10_axuser_7_reg[31:0] = int_desc_10_axuser_7_axuser;
assign uc2rb_desc_10_axuser_8_reg[31:0] = int_desc_10_axuser_8_axuser;
assign uc2rb_desc_10_axuser_9_reg[31:0] = int_desc_10_axuser_9_axuser;
assign uc2rb_desc_10_axuser_10_reg[31:0] = int_desc_10_axuser_10_axuser;
assign uc2rb_desc_10_axuser_11_reg[31:0] = int_desc_10_axuser_11_axuser;
assign uc2rb_desc_10_axuser_12_reg[31:0] = int_desc_10_axuser_12_axuser;
assign uc2rb_desc_10_axuser_13_reg[31:0] = int_desc_10_axuser_13_axuser;
assign uc2rb_desc_10_axuser_14_reg[31:0] = int_desc_10_axuser_14_axuser;
assign uc2rb_desc_10_axuser_15_reg[31:0] = int_desc_10_axuser_15_axuser;
assign uc2rb_desc_10_size_reg[15:0] = int_desc_10_size_txn_size;
assign uc2rb_desc_10_axsize_reg[2:0] = int_desc_10_axsize_axsize;
assign uc2rb_desc_10_axaddr_0_reg[31:0] = int_desc_10_axaddr_0_addr;
assign uc2rb_desc_10_axaddr_1_reg[31:0] = int_desc_10_axaddr_1_addr;
assign uc2rb_desc_10_axaddr_2_reg[31:0] = int_desc_10_axaddr_2_addr;
assign uc2rb_desc_10_axaddr_3_reg[31:0] = int_desc_10_axaddr_3_addr;
assign uc2rb_desc_10_data_offset_reg[31:0] = int_desc_10_data_offset_addr;
assign uc2rb_desc_10_wuser_0_reg[31:0] = int_desc_10_wuser_0_wuser;
assign uc2rb_desc_10_wuser_1_reg[31:0] = int_desc_10_wuser_1_wuser;
assign uc2rb_desc_10_wuser_2_reg[31:0] = int_desc_10_wuser_2_wuser;
assign uc2rb_desc_10_wuser_3_reg[31:0] = int_desc_10_wuser_3_wuser;
assign uc2rb_desc_10_wuser_4_reg[31:0] = int_desc_10_wuser_4_wuser;
assign uc2rb_desc_10_wuser_5_reg[31:0] = int_desc_10_wuser_5_wuser;
assign uc2rb_desc_10_wuser_6_reg[31:0] = int_desc_10_wuser_6_wuser;
assign uc2rb_desc_10_wuser_7_reg[31:0] = int_desc_10_wuser_7_wuser;
assign uc2rb_desc_10_wuser_8_reg[31:0] = int_desc_10_wuser_8_wuser;
assign uc2rb_desc_10_wuser_9_reg[31:0] = int_desc_10_wuser_9_wuser;
assign uc2rb_desc_10_wuser_10_reg[31:0] = int_desc_10_wuser_10_wuser;
assign uc2rb_desc_10_wuser_11_reg[31:0] = int_desc_10_wuser_11_wuser;
assign uc2rb_desc_10_wuser_12_reg[31:0] = int_desc_10_wuser_12_wuser;
assign uc2rb_desc_10_wuser_13_reg[31:0] = int_desc_10_wuser_13_wuser;
assign uc2rb_desc_10_wuser_14_reg[31:0] = int_desc_10_wuser_14_wuser;
assign uc2rb_desc_10_wuser_15_reg[31:0] = int_desc_10_wuser_15_wuser;
assign uc2rb_desc_11_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_11_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_11_size_reg[31:16] = 16'h0;
assign uc2rb_desc_11_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_11_txn_type_reg[1] = int_desc_11_txn_type_wr_strb;
assign uc2rb_desc_11_txn_type_reg[0] = int_desc_11_txn_type_wr_rd;
assign uc2rb_desc_11_attr_reg[18:15] = int_desc_11_attr_axregion;
assign uc2rb_desc_11_attr_reg[14:11] = int_desc_11_attr_axqos;
assign uc2rb_desc_11_attr_reg[10:8] = int_desc_11_attr_axprot;
assign uc2rb_desc_11_attr_reg[7:4] = int_desc_11_attr_axcache;
assign uc2rb_desc_11_attr_reg[3:2] = int_desc_11_attr_axlock;
assign uc2rb_desc_11_attr_reg[1:0] = int_desc_11_attr_axburst;
assign uc2rb_desc_11_axid_0_reg[31:0] = int_desc_11_axid_0_axid;
assign uc2rb_desc_11_axid_1_reg[31:0] = int_desc_11_axid_1_axid;
assign uc2rb_desc_11_axid_2_reg[31:0] = int_desc_11_axid_2_axid;
assign uc2rb_desc_11_axid_3_reg[31:0] = int_desc_11_axid_3_axid;
assign uc2rb_desc_11_axuser_0_reg[31:0] = int_desc_11_axuser_0_axuser;
assign uc2rb_desc_11_axuser_1_reg[31:0] = int_desc_11_axuser_1_axuser;
assign uc2rb_desc_11_axuser_2_reg[31:0] = int_desc_11_axuser_2_axuser;
assign uc2rb_desc_11_axuser_3_reg[31:0] = int_desc_11_axuser_3_axuser;
assign uc2rb_desc_11_axuser_4_reg[31:0] = int_desc_11_axuser_4_axuser;
assign uc2rb_desc_11_axuser_5_reg[31:0] = int_desc_11_axuser_5_axuser;
assign uc2rb_desc_11_axuser_6_reg[31:0] = int_desc_11_axuser_6_axuser;
assign uc2rb_desc_11_axuser_7_reg[31:0] = int_desc_11_axuser_7_axuser;
assign uc2rb_desc_11_axuser_8_reg[31:0] = int_desc_11_axuser_8_axuser;
assign uc2rb_desc_11_axuser_9_reg[31:0] = int_desc_11_axuser_9_axuser;
assign uc2rb_desc_11_axuser_10_reg[31:0] = int_desc_11_axuser_10_axuser;
assign uc2rb_desc_11_axuser_11_reg[31:0] = int_desc_11_axuser_11_axuser;
assign uc2rb_desc_11_axuser_12_reg[31:0] = int_desc_11_axuser_12_axuser;
assign uc2rb_desc_11_axuser_13_reg[31:0] = int_desc_11_axuser_13_axuser;
assign uc2rb_desc_11_axuser_14_reg[31:0] = int_desc_11_axuser_14_axuser;
assign uc2rb_desc_11_axuser_15_reg[31:0] = int_desc_11_axuser_15_axuser;
assign uc2rb_desc_11_size_reg[15:0] = int_desc_11_size_txn_size;
assign uc2rb_desc_11_axsize_reg[2:0] = int_desc_11_axsize_axsize;
assign uc2rb_desc_11_axaddr_0_reg[31:0] = int_desc_11_axaddr_0_addr;
assign uc2rb_desc_11_axaddr_1_reg[31:0] = int_desc_11_axaddr_1_addr;
assign uc2rb_desc_11_axaddr_2_reg[31:0] = int_desc_11_axaddr_2_addr;
assign uc2rb_desc_11_axaddr_3_reg[31:0] = int_desc_11_axaddr_3_addr;
assign uc2rb_desc_11_data_offset_reg[31:0] = int_desc_11_data_offset_addr;
assign uc2rb_desc_11_wuser_0_reg[31:0] = int_desc_11_wuser_0_wuser;
assign uc2rb_desc_11_wuser_1_reg[31:0] = int_desc_11_wuser_1_wuser;
assign uc2rb_desc_11_wuser_2_reg[31:0] = int_desc_11_wuser_2_wuser;
assign uc2rb_desc_11_wuser_3_reg[31:0] = int_desc_11_wuser_3_wuser;
assign uc2rb_desc_11_wuser_4_reg[31:0] = int_desc_11_wuser_4_wuser;
assign uc2rb_desc_11_wuser_5_reg[31:0] = int_desc_11_wuser_5_wuser;
assign uc2rb_desc_11_wuser_6_reg[31:0] = int_desc_11_wuser_6_wuser;
assign uc2rb_desc_11_wuser_7_reg[31:0] = int_desc_11_wuser_7_wuser;
assign uc2rb_desc_11_wuser_8_reg[31:0] = int_desc_11_wuser_8_wuser;
assign uc2rb_desc_11_wuser_9_reg[31:0] = int_desc_11_wuser_9_wuser;
assign uc2rb_desc_11_wuser_10_reg[31:0] = int_desc_11_wuser_10_wuser;
assign uc2rb_desc_11_wuser_11_reg[31:0] = int_desc_11_wuser_11_wuser;
assign uc2rb_desc_11_wuser_12_reg[31:0] = int_desc_11_wuser_12_wuser;
assign uc2rb_desc_11_wuser_13_reg[31:0] = int_desc_11_wuser_13_wuser;
assign uc2rb_desc_11_wuser_14_reg[31:0] = int_desc_11_wuser_14_wuser;
assign uc2rb_desc_11_wuser_15_reg[31:0] = int_desc_11_wuser_15_wuser;
assign uc2rb_desc_12_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_12_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_12_size_reg[31:16] = 16'h0;
assign uc2rb_desc_12_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_12_txn_type_reg[1] = int_desc_12_txn_type_wr_strb;
assign uc2rb_desc_12_txn_type_reg[0] = int_desc_12_txn_type_wr_rd;
assign uc2rb_desc_12_attr_reg[18:15] = int_desc_12_attr_axregion;
assign uc2rb_desc_12_attr_reg[14:11] = int_desc_12_attr_axqos;
assign uc2rb_desc_12_attr_reg[10:8] = int_desc_12_attr_axprot;
assign uc2rb_desc_12_attr_reg[7:4] = int_desc_12_attr_axcache;
assign uc2rb_desc_12_attr_reg[3:2] = int_desc_12_attr_axlock;
assign uc2rb_desc_12_attr_reg[1:0] = int_desc_12_attr_axburst;
assign uc2rb_desc_12_axid_0_reg[31:0] = int_desc_12_axid_0_axid;
assign uc2rb_desc_12_axid_1_reg[31:0] = int_desc_12_axid_1_axid;
assign uc2rb_desc_12_axid_2_reg[31:0] = int_desc_12_axid_2_axid;
assign uc2rb_desc_12_axid_3_reg[31:0] = int_desc_12_axid_3_axid;
assign uc2rb_desc_12_axuser_0_reg[31:0] = int_desc_12_axuser_0_axuser;
assign uc2rb_desc_12_axuser_1_reg[31:0] = int_desc_12_axuser_1_axuser;
assign uc2rb_desc_12_axuser_2_reg[31:0] = int_desc_12_axuser_2_axuser;
assign uc2rb_desc_12_axuser_3_reg[31:0] = int_desc_12_axuser_3_axuser;
assign uc2rb_desc_12_axuser_4_reg[31:0] = int_desc_12_axuser_4_axuser;
assign uc2rb_desc_12_axuser_5_reg[31:0] = int_desc_12_axuser_5_axuser;
assign uc2rb_desc_12_axuser_6_reg[31:0] = int_desc_12_axuser_6_axuser;
assign uc2rb_desc_12_axuser_7_reg[31:0] = int_desc_12_axuser_7_axuser;
assign uc2rb_desc_12_axuser_8_reg[31:0] = int_desc_12_axuser_8_axuser;
assign uc2rb_desc_12_axuser_9_reg[31:0] = int_desc_12_axuser_9_axuser;
assign uc2rb_desc_12_axuser_10_reg[31:0] = int_desc_12_axuser_10_axuser;
assign uc2rb_desc_12_axuser_11_reg[31:0] = int_desc_12_axuser_11_axuser;
assign uc2rb_desc_12_axuser_12_reg[31:0] = int_desc_12_axuser_12_axuser;
assign uc2rb_desc_12_axuser_13_reg[31:0] = int_desc_12_axuser_13_axuser;
assign uc2rb_desc_12_axuser_14_reg[31:0] = int_desc_12_axuser_14_axuser;
assign uc2rb_desc_12_axuser_15_reg[31:0] = int_desc_12_axuser_15_axuser;
assign uc2rb_desc_12_size_reg[15:0] = int_desc_12_size_txn_size;
assign uc2rb_desc_12_axsize_reg[2:0] = int_desc_12_axsize_axsize;
assign uc2rb_desc_12_axaddr_0_reg[31:0] = int_desc_12_axaddr_0_addr;
assign uc2rb_desc_12_axaddr_1_reg[31:0] = int_desc_12_axaddr_1_addr;
assign uc2rb_desc_12_axaddr_2_reg[31:0] = int_desc_12_axaddr_2_addr;
assign uc2rb_desc_12_axaddr_3_reg[31:0] = int_desc_12_axaddr_3_addr;
assign uc2rb_desc_12_data_offset_reg[31:0] = int_desc_12_data_offset_addr;
assign uc2rb_desc_12_wuser_0_reg[31:0] = int_desc_12_wuser_0_wuser;
assign uc2rb_desc_12_wuser_1_reg[31:0] = int_desc_12_wuser_1_wuser;
assign uc2rb_desc_12_wuser_2_reg[31:0] = int_desc_12_wuser_2_wuser;
assign uc2rb_desc_12_wuser_3_reg[31:0] = int_desc_12_wuser_3_wuser;
assign uc2rb_desc_12_wuser_4_reg[31:0] = int_desc_12_wuser_4_wuser;
assign uc2rb_desc_12_wuser_5_reg[31:0] = int_desc_12_wuser_5_wuser;
assign uc2rb_desc_12_wuser_6_reg[31:0] = int_desc_12_wuser_6_wuser;
assign uc2rb_desc_12_wuser_7_reg[31:0] = int_desc_12_wuser_7_wuser;
assign uc2rb_desc_12_wuser_8_reg[31:0] = int_desc_12_wuser_8_wuser;
assign uc2rb_desc_12_wuser_9_reg[31:0] = int_desc_12_wuser_9_wuser;
assign uc2rb_desc_12_wuser_10_reg[31:0] = int_desc_12_wuser_10_wuser;
assign uc2rb_desc_12_wuser_11_reg[31:0] = int_desc_12_wuser_11_wuser;
assign uc2rb_desc_12_wuser_12_reg[31:0] = int_desc_12_wuser_12_wuser;
assign uc2rb_desc_12_wuser_13_reg[31:0] = int_desc_12_wuser_13_wuser;
assign uc2rb_desc_12_wuser_14_reg[31:0] = int_desc_12_wuser_14_wuser;
assign uc2rb_desc_12_wuser_15_reg[31:0] = int_desc_12_wuser_15_wuser;
assign uc2rb_desc_13_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_13_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_13_size_reg[31:16] = 16'h0;
assign uc2rb_desc_13_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_13_txn_type_reg[1] = int_desc_13_txn_type_wr_strb;
assign uc2rb_desc_13_txn_type_reg[0] = int_desc_13_txn_type_wr_rd;
assign uc2rb_desc_13_attr_reg[18:15] = int_desc_13_attr_axregion;
assign uc2rb_desc_13_attr_reg[14:11] = int_desc_13_attr_axqos;
assign uc2rb_desc_13_attr_reg[10:8] = int_desc_13_attr_axprot;
assign uc2rb_desc_13_attr_reg[7:4] = int_desc_13_attr_axcache;
assign uc2rb_desc_13_attr_reg[3:2] = int_desc_13_attr_axlock;
assign uc2rb_desc_13_attr_reg[1:0] = int_desc_13_attr_axburst;
assign uc2rb_desc_13_axid_0_reg[31:0] = int_desc_13_axid_0_axid;
assign uc2rb_desc_13_axid_1_reg[31:0] = int_desc_13_axid_1_axid;
assign uc2rb_desc_13_axid_2_reg[31:0] = int_desc_13_axid_2_axid;
assign uc2rb_desc_13_axid_3_reg[31:0] = int_desc_13_axid_3_axid;
assign uc2rb_desc_13_axuser_0_reg[31:0] = int_desc_13_axuser_0_axuser;
assign uc2rb_desc_13_axuser_1_reg[31:0] = int_desc_13_axuser_1_axuser;
assign uc2rb_desc_13_axuser_2_reg[31:0] = int_desc_13_axuser_2_axuser;
assign uc2rb_desc_13_axuser_3_reg[31:0] = int_desc_13_axuser_3_axuser;
assign uc2rb_desc_13_axuser_4_reg[31:0] = int_desc_13_axuser_4_axuser;
assign uc2rb_desc_13_axuser_5_reg[31:0] = int_desc_13_axuser_5_axuser;
assign uc2rb_desc_13_axuser_6_reg[31:0] = int_desc_13_axuser_6_axuser;
assign uc2rb_desc_13_axuser_7_reg[31:0] = int_desc_13_axuser_7_axuser;
assign uc2rb_desc_13_axuser_8_reg[31:0] = int_desc_13_axuser_8_axuser;
assign uc2rb_desc_13_axuser_9_reg[31:0] = int_desc_13_axuser_9_axuser;
assign uc2rb_desc_13_axuser_10_reg[31:0] = int_desc_13_axuser_10_axuser;
assign uc2rb_desc_13_axuser_11_reg[31:0] = int_desc_13_axuser_11_axuser;
assign uc2rb_desc_13_axuser_12_reg[31:0] = int_desc_13_axuser_12_axuser;
assign uc2rb_desc_13_axuser_13_reg[31:0] = int_desc_13_axuser_13_axuser;
assign uc2rb_desc_13_axuser_14_reg[31:0] = int_desc_13_axuser_14_axuser;
assign uc2rb_desc_13_axuser_15_reg[31:0] = int_desc_13_axuser_15_axuser;
assign uc2rb_desc_13_size_reg[15:0] = int_desc_13_size_txn_size;
assign uc2rb_desc_13_axsize_reg[2:0] = int_desc_13_axsize_axsize;
assign uc2rb_desc_13_axaddr_0_reg[31:0] = int_desc_13_axaddr_0_addr;
assign uc2rb_desc_13_axaddr_1_reg[31:0] = int_desc_13_axaddr_1_addr;
assign uc2rb_desc_13_axaddr_2_reg[31:0] = int_desc_13_axaddr_2_addr;
assign uc2rb_desc_13_axaddr_3_reg[31:0] = int_desc_13_axaddr_3_addr;
assign uc2rb_desc_13_data_offset_reg[31:0] = int_desc_13_data_offset_addr;
assign uc2rb_desc_13_wuser_0_reg[31:0] = int_desc_13_wuser_0_wuser;
assign uc2rb_desc_13_wuser_1_reg[31:0] = int_desc_13_wuser_1_wuser;
assign uc2rb_desc_13_wuser_2_reg[31:0] = int_desc_13_wuser_2_wuser;
assign uc2rb_desc_13_wuser_3_reg[31:0] = int_desc_13_wuser_3_wuser;
assign uc2rb_desc_13_wuser_4_reg[31:0] = int_desc_13_wuser_4_wuser;
assign uc2rb_desc_13_wuser_5_reg[31:0] = int_desc_13_wuser_5_wuser;
assign uc2rb_desc_13_wuser_6_reg[31:0] = int_desc_13_wuser_6_wuser;
assign uc2rb_desc_13_wuser_7_reg[31:0] = int_desc_13_wuser_7_wuser;
assign uc2rb_desc_13_wuser_8_reg[31:0] = int_desc_13_wuser_8_wuser;
assign uc2rb_desc_13_wuser_9_reg[31:0] = int_desc_13_wuser_9_wuser;
assign uc2rb_desc_13_wuser_10_reg[31:0] = int_desc_13_wuser_10_wuser;
assign uc2rb_desc_13_wuser_11_reg[31:0] = int_desc_13_wuser_11_wuser;
assign uc2rb_desc_13_wuser_12_reg[31:0] = int_desc_13_wuser_12_wuser;
assign uc2rb_desc_13_wuser_13_reg[31:0] = int_desc_13_wuser_13_wuser;
assign uc2rb_desc_13_wuser_14_reg[31:0] = int_desc_13_wuser_14_wuser;
assign uc2rb_desc_13_wuser_15_reg[31:0] = int_desc_13_wuser_15_wuser;
assign uc2rb_desc_14_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_14_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_14_size_reg[31:16] = 16'h0;
assign uc2rb_desc_14_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_14_txn_type_reg[1] = int_desc_14_txn_type_wr_strb;
assign uc2rb_desc_14_txn_type_reg[0] = int_desc_14_txn_type_wr_rd;
assign uc2rb_desc_14_attr_reg[18:15] = int_desc_14_attr_axregion;
assign uc2rb_desc_14_attr_reg[14:11] = int_desc_14_attr_axqos;
assign uc2rb_desc_14_attr_reg[10:8] = int_desc_14_attr_axprot;
assign uc2rb_desc_14_attr_reg[7:4] = int_desc_14_attr_axcache;
assign uc2rb_desc_14_attr_reg[3:2] = int_desc_14_attr_axlock;
assign uc2rb_desc_14_attr_reg[1:0] = int_desc_14_attr_axburst;
assign uc2rb_desc_14_axid_0_reg[31:0] = int_desc_14_axid_0_axid;
assign uc2rb_desc_14_axid_1_reg[31:0] = int_desc_14_axid_1_axid;
assign uc2rb_desc_14_axid_2_reg[31:0] = int_desc_14_axid_2_axid;
assign uc2rb_desc_14_axid_3_reg[31:0] = int_desc_14_axid_3_axid;
assign uc2rb_desc_14_axuser_0_reg[31:0] = int_desc_14_axuser_0_axuser;
assign uc2rb_desc_14_axuser_1_reg[31:0] = int_desc_14_axuser_1_axuser;
assign uc2rb_desc_14_axuser_2_reg[31:0] = int_desc_14_axuser_2_axuser;
assign uc2rb_desc_14_axuser_3_reg[31:0] = int_desc_14_axuser_3_axuser;
assign uc2rb_desc_14_axuser_4_reg[31:0] = int_desc_14_axuser_4_axuser;
assign uc2rb_desc_14_axuser_5_reg[31:0] = int_desc_14_axuser_5_axuser;
assign uc2rb_desc_14_axuser_6_reg[31:0] = int_desc_14_axuser_6_axuser;
assign uc2rb_desc_14_axuser_7_reg[31:0] = int_desc_14_axuser_7_axuser;
assign uc2rb_desc_14_axuser_8_reg[31:0] = int_desc_14_axuser_8_axuser;
assign uc2rb_desc_14_axuser_9_reg[31:0] = int_desc_14_axuser_9_axuser;
assign uc2rb_desc_14_axuser_10_reg[31:0] = int_desc_14_axuser_10_axuser;
assign uc2rb_desc_14_axuser_11_reg[31:0] = int_desc_14_axuser_11_axuser;
assign uc2rb_desc_14_axuser_12_reg[31:0] = int_desc_14_axuser_12_axuser;
assign uc2rb_desc_14_axuser_13_reg[31:0] = int_desc_14_axuser_13_axuser;
assign uc2rb_desc_14_axuser_14_reg[31:0] = int_desc_14_axuser_14_axuser;
assign uc2rb_desc_14_axuser_15_reg[31:0] = int_desc_14_axuser_15_axuser;
assign uc2rb_desc_14_size_reg[15:0] = int_desc_14_size_txn_size;
assign uc2rb_desc_14_axsize_reg[2:0] = int_desc_14_axsize_axsize;
assign uc2rb_desc_14_axaddr_0_reg[31:0] = int_desc_14_axaddr_0_addr;
assign uc2rb_desc_14_axaddr_1_reg[31:0] = int_desc_14_axaddr_1_addr;
assign uc2rb_desc_14_axaddr_2_reg[31:0] = int_desc_14_axaddr_2_addr;
assign uc2rb_desc_14_axaddr_3_reg[31:0] = int_desc_14_axaddr_3_addr;
assign uc2rb_desc_14_data_offset_reg[31:0] = int_desc_14_data_offset_addr;
assign uc2rb_desc_14_wuser_0_reg[31:0] = int_desc_14_wuser_0_wuser;
assign uc2rb_desc_14_wuser_1_reg[31:0] = int_desc_14_wuser_1_wuser;
assign uc2rb_desc_14_wuser_2_reg[31:0] = int_desc_14_wuser_2_wuser;
assign uc2rb_desc_14_wuser_3_reg[31:0] = int_desc_14_wuser_3_wuser;
assign uc2rb_desc_14_wuser_4_reg[31:0] = int_desc_14_wuser_4_wuser;
assign uc2rb_desc_14_wuser_5_reg[31:0] = int_desc_14_wuser_5_wuser;
assign uc2rb_desc_14_wuser_6_reg[31:0] = int_desc_14_wuser_6_wuser;
assign uc2rb_desc_14_wuser_7_reg[31:0] = int_desc_14_wuser_7_wuser;
assign uc2rb_desc_14_wuser_8_reg[31:0] = int_desc_14_wuser_8_wuser;
assign uc2rb_desc_14_wuser_9_reg[31:0] = int_desc_14_wuser_9_wuser;
assign uc2rb_desc_14_wuser_10_reg[31:0] = int_desc_14_wuser_10_wuser;
assign uc2rb_desc_14_wuser_11_reg[31:0] = int_desc_14_wuser_11_wuser;
assign uc2rb_desc_14_wuser_12_reg[31:0] = int_desc_14_wuser_12_wuser;
assign uc2rb_desc_14_wuser_13_reg[31:0] = int_desc_14_wuser_13_wuser;
assign uc2rb_desc_14_wuser_14_reg[31:0] = int_desc_14_wuser_14_wuser;
assign uc2rb_desc_14_wuser_15_reg[31:0] = int_desc_14_wuser_15_wuser;
assign uc2rb_desc_15_txn_type_reg[31:2] = 30'h0;
assign uc2rb_desc_15_attr_reg[31:19] = 13'h0;
assign uc2rb_desc_15_size_reg[31:16] = 16'h0;
assign uc2rb_desc_15_axsize_reg[31:3] = 29'h0;
assign uc2rb_desc_15_txn_type_reg[1] = int_desc_15_txn_type_wr_strb;
assign uc2rb_desc_15_txn_type_reg[0] = int_desc_15_txn_type_wr_rd;
assign uc2rb_desc_15_attr_reg[18:15] = int_desc_15_attr_axregion;
assign uc2rb_desc_15_attr_reg[14:11] = int_desc_15_attr_axqos;
assign uc2rb_desc_15_attr_reg[10:8] = int_desc_15_attr_axprot;
assign uc2rb_desc_15_attr_reg[7:4] = int_desc_15_attr_axcache;
assign uc2rb_desc_15_attr_reg[3:2] = int_desc_15_attr_axlock;
assign uc2rb_desc_15_attr_reg[1:0] = int_desc_15_attr_axburst;
assign uc2rb_desc_15_axid_0_reg[31:0] = int_desc_15_axid_0_axid;
assign uc2rb_desc_15_axid_1_reg[31:0] = int_desc_15_axid_1_axid;
assign uc2rb_desc_15_axid_2_reg[31:0] = int_desc_15_axid_2_axid;
assign uc2rb_desc_15_axid_3_reg[31:0] = int_desc_15_axid_3_axid;
assign uc2rb_desc_15_axuser_0_reg[31:0] = int_desc_15_axuser_0_axuser;
assign uc2rb_desc_15_axuser_1_reg[31:0] = int_desc_15_axuser_1_axuser;
assign uc2rb_desc_15_axuser_2_reg[31:0] = int_desc_15_axuser_2_axuser;
assign uc2rb_desc_15_axuser_3_reg[31:0] = int_desc_15_axuser_3_axuser;
assign uc2rb_desc_15_axuser_4_reg[31:0] = int_desc_15_axuser_4_axuser;
assign uc2rb_desc_15_axuser_5_reg[31:0] = int_desc_15_axuser_5_axuser;
assign uc2rb_desc_15_axuser_6_reg[31:0] = int_desc_15_axuser_6_axuser;
assign uc2rb_desc_15_axuser_7_reg[31:0] = int_desc_15_axuser_7_axuser;
assign uc2rb_desc_15_axuser_8_reg[31:0] = int_desc_15_axuser_8_axuser;
assign uc2rb_desc_15_axuser_9_reg[31:0] = int_desc_15_axuser_9_axuser;
assign uc2rb_desc_15_axuser_10_reg[31:0] = int_desc_15_axuser_10_axuser;
assign uc2rb_desc_15_axuser_11_reg[31:0] = int_desc_15_axuser_11_axuser;
assign uc2rb_desc_15_axuser_12_reg[31:0] = int_desc_15_axuser_12_axuser;
assign uc2rb_desc_15_axuser_13_reg[31:0] = int_desc_15_axuser_13_axuser;
assign uc2rb_desc_15_axuser_14_reg[31:0] = int_desc_15_axuser_14_axuser;
assign uc2rb_desc_15_axuser_15_reg[31:0] = int_desc_15_axuser_15_axuser;
assign uc2rb_desc_15_size_reg[15:0] = int_desc_15_size_txn_size;
assign uc2rb_desc_15_axsize_reg[2:0] = int_desc_15_axsize_axsize;
assign uc2rb_desc_15_axaddr_0_reg[31:0] = int_desc_15_axaddr_0_addr;
assign uc2rb_desc_15_axaddr_1_reg[31:0] = int_desc_15_axaddr_1_addr;
assign uc2rb_desc_15_axaddr_2_reg[31:0] = int_desc_15_axaddr_2_addr;
assign uc2rb_desc_15_axaddr_3_reg[31:0] = int_desc_15_axaddr_3_addr;
assign uc2rb_desc_15_data_offset_reg[31:0] = int_desc_15_data_offset_addr;
assign uc2rb_desc_15_wuser_0_reg[31:0] = int_desc_15_wuser_0_wuser;
assign uc2rb_desc_15_wuser_1_reg[31:0] = int_desc_15_wuser_1_wuser;
assign uc2rb_desc_15_wuser_2_reg[31:0] = int_desc_15_wuser_2_wuser;
assign uc2rb_desc_15_wuser_3_reg[31:0] = int_desc_15_wuser_3_wuser;
assign uc2rb_desc_15_wuser_4_reg[31:0] = int_desc_15_wuser_4_wuser;
assign uc2rb_desc_15_wuser_5_reg[31:0] = int_desc_15_wuser_5_wuser;
assign uc2rb_desc_15_wuser_6_reg[31:0] = int_desc_15_wuser_6_wuser;
assign uc2rb_desc_15_wuser_7_reg[31:0] = int_desc_15_wuser_7_wuser;
assign uc2rb_desc_15_wuser_8_reg[31:0] = int_desc_15_wuser_8_wuser;
assign uc2rb_desc_15_wuser_9_reg[31:0] = int_desc_15_wuser_9_wuser;
assign uc2rb_desc_15_wuser_10_reg[31:0] = int_desc_15_wuser_10_wuser;
assign uc2rb_desc_15_wuser_11_reg[31:0] = int_desc_15_wuser_11_wuser;
assign uc2rb_desc_15_wuser_12_reg[31:0] = int_desc_15_wuser_12_wuser;
assign uc2rb_desc_15_wuser_13_reg[31:0] = int_desc_15_wuser_13_wuser;
assign uc2rb_desc_15_wuser_14_reg[31:0] = int_desc_15_wuser_14_wuser;
assign uc2rb_desc_15_wuser_15_reg[31:0] = int_desc_15_wuser_15_wuser;

//////////////////////
//Instantiate slave_inf 
//////////////////////
slave_inf #(
         .EN_INTFS_AXI4(EN_INTFS_AXI4)
        ,.EN_INTFS_AXI4LITE(EN_INTFS_AXI4LITE)
        ,.EN_INTFS_AXI3(EN_INTFS_AXI3)
	,.ADDR_WIDTH(ADDR_WIDTH)
	,.DATA_WIDTH(DATA_WIDTH)
	,.ID_WIDTH(ID_WIDTH)
	,.AWUSER_WIDTH(AWUSER_WIDTH)
	,.WUSER_WIDTH(WUSER_WIDTH)
	,.BUSER_WIDTH(BUSER_WIDTH)
	,.ARUSER_WIDTH(ARUSER_WIDTH)
	,.RUSER_WIDTH(RUSER_WIDTH)
	,.RAM_SIZE(RAM_SIZE)
	,.MAX_DESC(MAX_DESC)
	,.FORCE_RESP_ORDER(FORCE_RESP_ORDER)        
) i_slave_inf(
	.axi_aclk(axi_aclk)
	,.axi_aresetn(axi_aresetn)
	,.s_axi_usr_awready(s_axi_usr_awready)
	,.s_axi_usr_wready(s_axi_usr_wready)
	,.s_axi_usr_bid(s_axi_usr_bid)
	,.s_axi_usr_bresp(s_axi_usr_bresp)
	,.s_axi_usr_buser(s_axi_usr_buser)
	,.s_axi_usr_bvalid(s_axi_usr_bvalid)
	,.s_axi_usr_arready(s_axi_usr_arready)
	,.s_axi_usr_rid(s_axi_usr_rid)
	,.s_axi_usr_rdata(s_axi_usr_rdata)
	,.s_axi_usr_rresp(s_axi_usr_rresp)
	,.s_axi_usr_rlast(s_axi_usr_rlast)
	,.s_axi_usr_ruser(s_axi_usr_ruser)
	,.s_axi_usr_rvalid(s_axi_usr_rvalid)
	,.s_axi_usr_awid(s_axi_usr_awid)
	,.s_axi_usr_awaddr(s_axi_usr_awaddr)
	,.s_axi_usr_awlen(s_axi_usr_awlen)
	,.s_axi_usr_awsize(s_axi_usr_awsize)
	,.s_axi_usr_awburst(s_axi_usr_awburst)
	,.s_axi_usr_awlock(s_axi_usr_awlock)
	,.s_axi_usr_awcache(s_axi_usr_awcache)
	,.s_axi_usr_awprot(s_axi_usr_awprot)
	,.s_axi_usr_awqos(s_axi_usr_awqos)
	,.s_axi_usr_awregion(s_axi_usr_awregion)
	,.s_axi_usr_awuser(s_axi_usr_awuser)
	,.s_axi_usr_awvalid(s_axi_usr_awvalid)
	,.s_axi_usr_wdata(s_axi_usr_wdata)
	,.s_axi_usr_wstrb(s_axi_usr_wstrb)
	,.s_axi_usr_wlast(s_axi_usr_wlast)
	,.s_axi_usr_wid(s_axi_usr_wid)
	,.s_axi_usr_wuser(s_axi_usr_wuser)
	,.s_axi_usr_wvalid(s_axi_usr_wvalid)
	,.s_axi_usr_bready(s_axi_usr_bready)
	,.s_axi_usr_arid(s_axi_usr_arid)
	,.s_axi_usr_araddr(s_axi_usr_araddr)
	,.s_axi_usr_arlen(s_axi_usr_arlen)
	,.s_axi_usr_arsize(s_axi_usr_arsize)
	,.s_axi_usr_arburst(s_axi_usr_arburst)
	,.s_axi_usr_arlock(s_axi_usr_arlock)
	,.s_axi_usr_arcache(s_axi_usr_arcache)
	,.s_axi_usr_arprot(s_axi_usr_arprot)
	,.s_axi_usr_arqos(s_axi_usr_arqos)
	,.s_axi_usr_arregion(s_axi_usr_arregion)
	,.s_axi_usr_aruser(s_axi_usr_aruser)
	,.s_axi_usr_arvalid(s_axi_usr_arvalid)
	,.s_axi_usr_rready(s_axi_usr_rready)
        ,.int_ownership_own(int_ownership_own)
	,.int_status_busy_busy(int_status_busy_busy)
	,.int_resp_fifo_free_level_level(int_resp_fifo_free_level_level)
	,.int_intr_txn_avail_status_avail(int_intr_txn_avail_status_avail)
	,.int_intr_comp_status_comp(int_intr_comp_status_comp)
	,.int_intr_error_status_err_0(int_intr_error_status_err_0)
        ,.int_resp_order_field(int_resp_order_field)
	,.int_desc_0_txn_type_wr_strb(int_desc_0_txn_type_wr_strb)
	,.int_desc_0_txn_type_wr_rd(int_desc_0_txn_type_wr_rd)
	,.int_desc_0_attr_axregion(int_desc_0_attr_axregion)
	,.int_desc_0_attr_axqos(int_desc_0_attr_axqos)
	,.int_desc_0_attr_axprot(int_desc_0_attr_axprot)
	,.int_desc_0_attr_axcache(int_desc_0_attr_axcache)
	,.int_desc_0_attr_axlock(int_desc_0_attr_axlock)
	,.int_desc_0_attr_axburst(int_desc_0_attr_axburst)
	,.int_desc_0_axid_0_axid(int_desc_0_axid_0_axid)
	,.int_desc_0_axid_1_axid(int_desc_0_axid_1_axid)
	,.int_desc_0_axid_2_axid(int_desc_0_axid_2_axid)
	,.int_desc_0_axid_3_axid(int_desc_0_axid_3_axid)
	,.int_desc_0_axuser_0_axuser(int_desc_0_axuser_0_axuser)
	,.int_desc_0_axuser_1_axuser(int_desc_0_axuser_1_axuser)
	,.int_desc_0_axuser_2_axuser(int_desc_0_axuser_2_axuser)
	,.int_desc_0_axuser_3_axuser(int_desc_0_axuser_3_axuser)
	,.int_desc_0_axuser_4_axuser(int_desc_0_axuser_4_axuser)
	,.int_desc_0_axuser_5_axuser(int_desc_0_axuser_5_axuser)
	,.int_desc_0_axuser_6_axuser(int_desc_0_axuser_6_axuser)
	,.int_desc_0_axuser_7_axuser(int_desc_0_axuser_7_axuser)
	,.int_desc_0_axuser_8_axuser(int_desc_0_axuser_8_axuser)
	,.int_desc_0_axuser_9_axuser(int_desc_0_axuser_9_axuser)
	,.int_desc_0_axuser_10_axuser(int_desc_0_axuser_10_axuser)
	,.int_desc_0_axuser_11_axuser(int_desc_0_axuser_11_axuser)
	,.int_desc_0_axuser_12_axuser(int_desc_0_axuser_12_axuser)
	,.int_desc_0_axuser_13_axuser(int_desc_0_axuser_13_axuser)
	,.int_desc_0_axuser_14_axuser(int_desc_0_axuser_14_axuser)
	,.int_desc_0_axuser_15_axuser(int_desc_0_axuser_15_axuser)
	,.int_desc_0_size_txn_size(int_desc_0_size_txn_size)
	,.int_desc_0_axsize_axsize(int_desc_0_axsize_axsize)
	,.int_desc_0_axaddr_0_addr(int_desc_0_axaddr_0_addr)
	,.int_desc_0_axaddr_1_addr(int_desc_0_axaddr_1_addr)
	,.int_desc_0_axaddr_2_addr(int_desc_0_axaddr_2_addr)
	,.int_desc_0_axaddr_3_addr(int_desc_0_axaddr_3_addr)
	,.int_desc_0_data_offset_addr(int_desc_0_data_offset_addr)
	,.int_desc_0_wuser_0_wuser(int_desc_0_wuser_0_wuser)
	,.int_desc_0_wuser_1_wuser(int_desc_0_wuser_1_wuser)
	,.int_desc_0_wuser_2_wuser(int_desc_0_wuser_2_wuser)
	,.int_desc_0_wuser_3_wuser(int_desc_0_wuser_3_wuser)
	,.int_desc_0_wuser_4_wuser(int_desc_0_wuser_4_wuser)
	,.int_desc_0_wuser_5_wuser(int_desc_0_wuser_5_wuser)
	,.int_desc_0_wuser_6_wuser(int_desc_0_wuser_6_wuser)
	,.int_desc_0_wuser_7_wuser(int_desc_0_wuser_7_wuser)
	,.int_desc_0_wuser_8_wuser(int_desc_0_wuser_8_wuser)
	,.int_desc_0_wuser_9_wuser(int_desc_0_wuser_9_wuser)
	,.int_desc_0_wuser_10_wuser(int_desc_0_wuser_10_wuser)
	,.int_desc_0_wuser_11_wuser(int_desc_0_wuser_11_wuser)
	,.int_desc_0_wuser_12_wuser(int_desc_0_wuser_12_wuser)
	,.int_desc_0_wuser_13_wuser(int_desc_0_wuser_13_wuser)
	,.int_desc_0_wuser_14_wuser(int_desc_0_wuser_14_wuser)
	,.int_desc_0_wuser_15_wuser(int_desc_0_wuser_15_wuser)
	,.int_desc_1_txn_type_wr_strb(int_desc_1_txn_type_wr_strb)
	,.int_desc_1_txn_type_wr_rd(int_desc_1_txn_type_wr_rd)
	,.int_desc_1_attr_axregion(int_desc_1_attr_axregion)
	,.int_desc_1_attr_axqos(int_desc_1_attr_axqos)
	,.int_desc_1_attr_axprot(int_desc_1_attr_axprot)
	,.int_desc_1_attr_axcache(int_desc_1_attr_axcache)
	,.int_desc_1_attr_axlock(int_desc_1_attr_axlock)
	,.int_desc_1_attr_axburst(int_desc_1_attr_axburst)
	,.int_desc_1_axid_0_axid(int_desc_1_axid_0_axid)
	,.int_desc_1_axid_1_axid(int_desc_1_axid_1_axid)
	,.int_desc_1_axid_2_axid(int_desc_1_axid_2_axid)
	,.int_desc_1_axid_3_axid(int_desc_1_axid_3_axid)
	,.int_desc_1_axuser_0_axuser(int_desc_1_axuser_0_axuser)
	,.int_desc_1_axuser_1_axuser(int_desc_1_axuser_1_axuser)
	,.int_desc_1_axuser_2_axuser(int_desc_1_axuser_2_axuser)
	,.int_desc_1_axuser_3_axuser(int_desc_1_axuser_3_axuser)
	,.int_desc_1_axuser_4_axuser(int_desc_1_axuser_4_axuser)
	,.int_desc_1_axuser_5_axuser(int_desc_1_axuser_5_axuser)
	,.int_desc_1_axuser_6_axuser(int_desc_1_axuser_6_axuser)
	,.int_desc_1_axuser_7_axuser(int_desc_1_axuser_7_axuser)
	,.int_desc_1_axuser_8_axuser(int_desc_1_axuser_8_axuser)
	,.int_desc_1_axuser_9_axuser(int_desc_1_axuser_9_axuser)
	,.int_desc_1_axuser_10_axuser(int_desc_1_axuser_10_axuser)
	,.int_desc_1_axuser_11_axuser(int_desc_1_axuser_11_axuser)
	,.int_desc_1_axuser_12_axuser(int_desc_1_axuser_12_axuser)
	,.int_desc_1_axuser_13_axuser(int_desc_1_axuser_13_axuser)
	,.int_desc_1_axuser_14_axuser(int_desc_1_axuser_14_axuser)
	,.int_desc_1_axuser_15_axuser(int_desc_1_axuser_15_axuser)
	,.int_desc_1_size_txn_size(int_desc_1_size_txn_size)
	,.int_desc_1_axsize_axsize(int_desc_1_axsize_axsize)
	,.int_desc_1_axaddr_0_addr(int_desc_1_axaddr_0_addr)
	,.int_desc_1_axaddr_1_addr(int_desc_1_axaddr_1_addr)
	,.int_desc_1_axaddr_2_addr(int_desc_1_axaddr_2_addr)
	,.int_desc_1_axaddr_3_addr(int_desc_1_axaddr_3_addr)
	,.int_desc_1_data_offset_addr(int_desc_1_data_offset_addr)
	,.int_desc_1_wuser_0_wuser(int_desc_1_wuser_0_wuser)
	,.int_desc_1_wuser_1_wuser(int_desc_1_wuser_1_wuser)
	,.int_desc_1_wuser_2_wuser(int_desc_1_wuser_2_wuser)
	,.int_desc_1_wuser_3_wuser(int_desc_1_wuser_3_wuser)
	,.int_desc_1_wuser_4_wuser(int_desc_1_wuser_4_wuser)
	,.int_desc_1_wuser_5_wuser(int_desc_1_wuser_5_wuser)
	,.int_desc_1_wuser_6_wuser(int_desc_1_wuser_6_wuser)
	,.int_desc_1_wuser_7_wuser(int_desc_1_wuser_7_wuser)
	,.int_desc_1_wuser_8_wuser(int_desc_1_wuser_8_wuser)
	,.int_desc_1_wuser_9_wuser(int_desc_1_wuser_9_wuser)
	,.int_desc_1_wuser_10_wuser(int_desc_1_wuser_10_wuser)
	,.int_desc_1_wuser_11_wuser(int_desc_1_wuser_11_wuser)
	,.int_desc_1_wuser_12_wuser(int_desc_1_wuser_12_wuser)
	,.int_desc_1_wuser_13_wuser(int_desc_1_wuser_13_wuser)
	,.int_desc_1_wuser_14_wuser(int_desc_1_wuser_14_wuser)
	,.int_desc_1_wuser_15_wuser(int_desc_1_wuser_15_wuser)
	,.int_desc_2_txn_type_wr_strb(int_desc_2_txn_type_wr_strb)
	,.int_desc_2_txn_type_wr_rd(int_desc_2_txn_type_wr_rd)
	,.int_desc_2_attr_axregion(int_desc_2_attr_axregion)
	,.int_desc_2_attr_axqos(int_desc_2_attr_axqos)
	,.int_desc_2_attr_axprot(int_desc_2_attr_axprot)
	,.int_desc_2_attr_axcache(int_desc_2_attr_axcache)
	,.int_desc_2_attr_axlock(int_desc_2_attr_axlock)
	,.int_desc_2_attr_axburst(int_desc_2_attr_axburst)
	,.int_desc_2_axid_0_axid(int_desc_2_axid_0_axid)
	,.int_desc_2_axid_1_axid(int_desc_2_axid_1_axid)
	,.int_desc_2_axid_2_axid(int_desc_2_axid_2_axid)
	,.int_desc_2_axid_3_axid(int_desc_2_axid_3_axid)
	,.int_desc_2_axuser_0_axuser(int_desc_2_axuser_0_axuser)
	,.int_desc_2_axuser_1_axuser(int_desc_2_axuser_1_axuser)
	,.int_desc_2_axuser_2_axuser(int_desc_2_axuser_2_axuser)
	,.int_desc_2_axuser_3_axuser(int_desc_2_axuser_3_axuser)
	,.int_desc_2_axuser_4_axuser(int_desc_2_axuser_4_axuser)
	,.int_desc_2_axuser_5_axuser(int_desc_2_axuser_5_axuser)
	,.int_desc_2_axuser_6_axuser(int_desc_2_axuser_6_axuser)
	,.int_desc_2_axuser_7_axuser(int_desc_2_axuser_7_axuser)
	,.int_desc_2_axuser_8_axuser(int_desc_2_axuser_8_axuser)
	,.int_desc_2_axuser_9_axuser(int_desc_2_axuser_9_axuser)
	,.int_desc_2_axuser_10_axuser(int_desc_2_axuser_10_axuser)
	,.int_desc_2_axuser_11_axuser(int_desc_2_axuser_11_axuser)
	,.int_desc_2_axuser_12_axuser(int_desc_2_axuser_12_axuser)
	,.int_desc_2_axuser_13_axuser(int_desc_2_axuser_13_axuser)
	,.int_desc_2_axuser_14_axuser(int_desc_2_axuser_14_axuser)
	,.int_desc_2_axuser_15_axuser(int_desc_2_axuser_15_axuser)
	,.int_desc_2_size_txn_size(int_desc_2_size_txn_size)
	,.int_desc_2_axsize_axsize(int_desc_2_axsize_axsize)
	,.int_desc_2_axaddr_0_addr(int_desc_2_axaddr_0_addr)
	,.int_desc_2_axaddr_1_addr(int_desc_2_axaddr_1_addr)
	,.int_desc_2_axaddr_2_addr(int_desc_2_axaddr_2_addr)
	,.int_desc_2_axaddr_3_addr(int_desc_2_axaddr_3_addr)
	,.int_desc_2_data_offset_addr(int_desc_2_data_offset_addr)
	,.int_desc_2_wuser_0_wuser(int_desc_2_wuser_0_wuser)
	,.int_desc_2_wuser_1_wuser(int_desc_2_wuser_1_wuser)
	,.int_desc_2_wuser_2_wuser(int_desc_2_wuser_2_wuser)
	,.int_desc_2_wuser_3_wuser(int_desc_2_wuser_3_wuser)
	,.int_desc_2_wuser_4_wuser(int_desc_2_wuser_4_wuser)
	,.int_desc_2_wuser_5_wuser(int_desc_2_wuser_5_wuser)
	,.int_desc_2_wuser_6_wuser(int_desc_2_wuser_6_wuser)
	,.int_desc_2_wuser_7_wuser(int_desc_2_wuser_7_wuser)
	,.int_desc_2_wuser_8_wuser(int_desc_2_wuser_8_wuser)
	,.int_desc_2_wuser_9_wuser(int_desc_2_wuser_9_wuser)
	,.int_desc_2_wuser_10_wuser(int_desc_2_wuser_10_wuser)
	,.int_desc_2_wuser_11_wuser(int_desc_2_wuser_11_wuser)
	,.int_desc_2_wuser_12_wuser(int_desc_2_wuser_12_wuser)
	,.int_desc_2_wuser_13_wuser(int_desc_2_wuser_13_wuser)
	,.int_desc_2_wuser_14_wuser(int_desc_2_wuser_14_wuser)
	,.int_desc_2_wuser_15_wuser(int_desc_2_wuser_15_wuser)
	,.int_desc_3_txn_type_wr_strb(int_desc_3_txn_type_wr_strb)
	,.int_desc_3_txn_type_wr_rd(int_desc_3_txn_type_wr_rd)
	,.int_desc_3_attr_axregion(int_desc_3_attr_axregion)
	,.int_desc_3_attr_axqos(int_desc_3_attr_axqos)
	,.int_desc_3_attr_axprot(int_desc_3_attr_axprot)
	,.int_desc_3_attr_axcache(int_desc_3_attr_axcache)
	,.int_desc_3_attr_axlock(int_desc_3_attr_axlock)
	,.int_desc_3_attr_axburst(int_desc_3_attr_axburst)
	,.int_desc_3_axid_0_axid(int_desc_3_axid_0_axid)
	,.int_desc_3_axid_1_axid(int_desc_3_axid_1_axid)
	,.int_desc_3_axid_2_axid(int_desc_3_axid_2_axid)
	,.int_desc_3_axid_3_axid(int_desc_3_axid_3_axid)
	,.int_desc_3_axuser_0_axuser(int_desc_3_axuser_0_axuser)
	,.int_desc_3_axuser_1_axuser(int_desc_3_axuser_1_axuser)
	,.int_desc_3_axuser_2_axuser(int_desc_3_axuser_2_axuser)
	,.int_desc_3_axuser_3_axuser(int_desc_3_axuser_3_axuser)
	,.int_desc_3_axuser_4_axuser(int_desc_3_axuser_4_axuser)
	,.int_desc_3_axuser_5_axuser(int_desc_3_axuser_5_axuser)
	,.int_desc_3_axuser_6_axuser(int_desc_3_axuser_6_axuser)
	,.int_desc_3_axuser_7_axuser(int_desc_3_axuser_7_axuser)
	,.int_desc_3_axuser_8_axuser(int_desc_3_axuser_8_axuser)
	,.int_desc_3_axuser_9_axuser(int_desc_3_axuser_9_axuser)
	,.int_desc_3_axuser_10_axuser(int_desc_3_axuser_10_axuser)
	,.int_desc_3_axuser_11_axuser(int_desc_3_axuser_11_axuser)
	,.int_desc_3_axuser_12_axuser(int_desc_3_axuser_12_axuser)
	,.int_desc_3_axuser_13_axuser(int_desc_3_axuser_13_axuser)
	,.int_desc_3_axuser_14_axuser(int_desc_3_axuser_14_axuser)
	,.int_desc_3_axuser_15_axuser(int_desc_3_axuser_15_axuser)
	,.int_desc_3_size_txn_size(int_desc_3_size_txn_size)
	,.int_desc_3_axsize_axsize(int_desc_3_axsize_axsize)
	,.int_desc_3_axaddr_0_addr(int_desc_3_axaddr_0_addr)
	,.int_desc_3_axaddr_1_addr(int_desc_3_axaddr_1_addr)
	,.int_desc_3_axaddr_2_addr(int_desc_3_axaddr_2_addr)
	,.int_desc_3_axaddr_3_addr(int_desc_3_axaddr_3_addr)
	,.int_desc_3_data_offset_addr(int_desc_3_data_offset_addr)
	,.int_desc_3_wuser_0_wuser(int_desc_3_wuser_0_wuser)
	,.int_desc_3_wuser_1_wuser(int_desc_3_wuser_1_wuser)
	,.int_desc_3_wuser_2_wuser(int_desc_3_wuser_2_wuser)
	,.int_desc_3_wuser_3_wuser(int_desc_3_wuser_3_wuser)
	,.int_desc_3_wuser_4_wuser(int_desc_3_wuser_4_wuser)
	,.int_desc_3_wuser_5_wuser(int_desc_3_wuser_5_wuser)
	,.int_desc_3_wuser_6_wuser(int_desc_3_wuser_6_wuser)
	,.int_desc_3_wuser_7_wuser(int_desc_3_wuser_7_wuser)
	,.int_desc_3_wuser_8_wuser(int_desc_3_wuser_8_wuser)
	,.int_desc_3_wuser_9_wuser(int_desc_3_wuser_9_wuser)
	,.int_desc_3_wuser_10_wuser(int_desc_3_wuser_10_wuser)
	,.int_desc_3_wuser_11_wuser(int_desc_3_wuser_11_wuser)
	,.int_desc_3_wuser_12_wuser(int_desc_3_wuser_12_wuser)
	,.int_desc_3_wuser_13_wuser(int_desc_3_wuser_13_wuser)
	,.int_desc_3_wuser_14_wuser(int_desc_3_wuser_14_wuser)
	,.int_desc_3_wuser_15_wuser(int_desc_3_wuser_15_wuser)
	,.int_desc_4_txn_type_wr_strb(int_desc_4_txn_type_wr_strb)
	,.int_desc_4_txn_type_wr_rd(int_desc_4_txn_type_wr_rd)
	,.int_desc_4_attr_axregion(int_desc_4_attr_axregion)
	,.int_desc_4_attr_axqos(int_desc_4_attr_axqos)
	,.int_desc_4_attr_axprot(int_desc_4_attr_axprot)
	,.int_desc_4_attr_axcache(int_desc_4_attr_axcache)
	,.int_desc_4_attr_axlock(int_desc_4_attr_axlock)
	,.int_desc_4_attr_axburst(int_desc_4_attr_axburst)
	,.int_desc_4_axid_0_axid(int_desc_4_axid_0_axid)
	,.int_desc_4_axid_1_axid(int_desc_4_axid_1_axid)
	,.int_desc_4_axid_2_axid(int_desc_4_axid_2_axid)
	,.int_desc_4_axid_3_axid(int_desc_4_axid_3_axid)
	,.int_desc_4_axuser_0_axuser(int_desc_4_axuser_0_axuser)
	,.int_desc_4_axuser_1_axuser(int_desc_4_axuser_1_axuser)
	,.int_desc_4_axuser_2_axuser(int_desc_4_axuser_2_axuser)
	,.int_desc_4_axuser_3_axuser(int_desc_4_axuser_3_axuser)
	,.int_desc_4_axuser_4_axuser(int_desc_4_axuser_4_axuser)
	,.int_desc_4_axuser_5_axuser(int_desc_4_axuser_5_axuser)
	,.int_desc_4_axuser_6_axuser(int_desc_4_axuser_6_axuser)
	,.int_desc_4_axuser_7_axuser(int_desc_4_axuser_7_axuser)
	,.int_desc_4_axuser_8_axuser(int_desc_4_axuser_8_axuser)
	,.int_desc_4_axuser_9_axuser(int_desc_4_axuser_9_axuser)
	,.int_desc_4_axuser_10_axuser(int_desc_4_axuser_10_axuser)
	,.int_desc_4_axuser_11_axuser(int_desc_4_axuser_11_axuser)
	,.int_desc_4_axuser_12_axuser(int_desc_4_axuser_12_axuser)
	,.int_desc_4_axuser_13_axuser(int_desc_4_axuser_13_axuser)
	,.int_desc_4_axuser_14_axuser(int_desc_4_axuser_14_axuser)
	,.int_desc_4_axuser_15_axuser(int_desc_4_axuser_15_axuser)
	,.int_desc_4_size_txn_size(int_desc_4_size_txn_size)
	,.int_desc_4_axsize_axsize(int_desc_4_axsize_axsize)
	,.int_desc_4_axaddr_0_addr(int_desc_4_axaddr_0_addr)
	,.int_desc_4_axaddr_1_addr(int_desc_4_axaddr_1_addr)
	,.int_desc_4_axaddr_2_addr(int_desc_4_axaddr_2_addr)
	,.int_desc_4_axaddr_3_addr(int_desc_4_axaddr_3_addr)
	,.int_desc_4_data_offset_addr(int_desc_4_data_offset_addr)
	,.int_desc_4_wuser_0_wuser(int_desc_4_wuser_0_wuser)
	,.int_desc_4_wuser_1_wuser(int_desc_4_wuser_1_wuser)
	,.int_desc_4_wuser_2_wuser(int_desc_4_wuser_2_wuser)
	,.int_desc_4_wuser_3_wuser(int_desc_4_wuser_3_wuser)
	,.int_desc_4_wuser_4_wuser(int_desc_4_wuser_4_wuser)
	,.int_desc_4_wuser_5_wuser(int_desc_4_wuser_5_wuser)
	,.int_desc_4_wuser_6_wuser(int_desc_4_wuser_6_wuser)
	,.int_desc_4_wuser_7_wuser(int_desc_4_wuser_7_wuser)
	,.int_desc_4_wuser_8_wuser(int_desc_4_wuser_8_wuser)
	,.int_desc_4_wuser_9_wuser(int_desc_4_wuser_9_wuser)
	,.int_desc_4_wuser_10_wuser(int_desc_4_wuser_10_wuser)
	,.int_desc_4_wuser_11_wuser(int_desc_4_wuser_11_wuser)
	,.int_desc_4_wuser_12_wuser(int_desc_4_wuser_12_wuser)
	,.int_desc_4_wuser_13_wuser(int_desc_4_wuser_13_wuser)
	,.int_desc_4_wuser_14_wuser(int_desc_4_wuser_14_wuser)
	,.int_desc_4_wuser_15_wuser(int_desc_4_wuser_15_wuser)
	,.int_desc_5_txn_type_wr_strb(int_desc_5_txn_type_wr_strb)
	,.int_desc_5_txn_type_wr_rd(int_desc_5_txn_type_wr_rd)
	,.int_desc_5_attr_axregion(int_desc_5_attr_axregion)
	,.int_desc_5_attr_axqos(int_desc_5_attr_axqos)
	,.int_desc_5_attr_axprot(int_desc_5_attr_axprot)
	,.int_desc_5_attr_axcache(int_desc_5_attr_axcache)
	,.int_desc_5_attr_axlock(int_desc_5_attr_axlock)
	,.int_desc_5_attr_axburst(int_desc_5_attr_axburst)
	,.int_desc_5_axid_0_axid(int_desc_5_axid_0_axid)
	,.int_desc_5_axid_1_axid(int_desc_5_axid_1_axid)
	,.int_desc_5_axid_2_axid(int_desc_5_axid_2_axid)
	,.int_desc_5_axid_3_axid(int_desc_5_axid_3_axid)
	,.int_desc_5_axuser_0_axuser(int_desc_5_axuser_0_axuser)
	,.int_desc_5_axuser_1_axuser(int_desc_5_axuser_1_axuser)
	,.int_desc_5_axuser_2_axuser(int_desc_5_axuser_2_axuser)
	,.int_desc_5_axuser_3_axuser(int_desc_5_axuser_3_axuser)
	,.int_desc_5_axuser_4_axuser(int_desc_5_axuser_4_axuser)
	,.int_desc_5_axuser_5_axuser(int_desc_5_axuser_5_axuser)
	,.int_desc_5_axuser_6_axuser(int_desc_5_axuser_6_axuser)
	,.int_desc_5_axuser_7_axuser(int_desc_5_axuser_7_axuser)
	,.int_desc_5_axuser_8_axuser(int_desc_5_axuser_8_axuser)
	,.int_desc_5_axuser_9_axuser(int_desc_5_axuser_9_axuser)
	,.int_desc_5_axuser_10_axuser(int_desc_5_axuser_10_axuser)
	,.int_desc_5_axuser_11_axuser(int_desc_5_axuser_11_axuser)
	,.int_desc_5_axuser_12_axuser(int_desc_5_axuser_12_axuser)
	,.int_desc_5_axuser_13_axuser(int_desc_5_axuser_13_axuser)
	,.int_desc_5_axuser_14_axuser(int_desc_5_axuser_14_axuser)
	,.int_desc_5_axuser_15_axuser(int_desc_5_axuser_15_axuser)
	,.int_desc_5_size_txn_size(int_desc_5_size_txn_size)
	,.int_desc_5_axsize_axsize(int_desc_5_axsize_axsize)
	,.int_desc_5_axaddr_0_addr(int_desc_5_axaddr_0_addr)
	,.int_desc_5_axaddr_1_addr(int_desc_5_axaddr_1_addr)
	,.int_desc_5_axaddr_2_addr(int_desc_5_axaddr_2_addr)
	,.int_desc_5_axaddr_3_addr(int_desc_5_axaddr_3_addr)
	,.int_desc_5_data_offset_addr(int_desc_5_data_offset_addr)
	,.int_desc_5_wuser_0_wuser(int_desc_5_wuser_0_wuser)
	,.int_desc_5_wuser_1_wuser(int_desc_5_wuser_1_wuser)
	,.int_desc_5_wuser_2_wuser(int_desc_5_wuser_2_wuser)
	,.int_desc_5_wuser_3_wuser(int_desc_5_wuser_3_wuser)
	,.int_desc_5_wuser_4_wuser(int_desc_5_wuser_4_wuser)
	,.int_desc_5_wuser_5_wuser(int_desc_5_wuser_5_wuser)
	,.int_desc_5_wuser_6_wuser(int_desc_5_wuser_6_wuser)
	,.int_desc_5_wuser_7_wuser(int_desc_5_wuser_7_wuser)
	,.int_desc_5_wuser_8_wuser(int_desc_5_wuser_8_wuser)
	,.int_desc_5_wuser_9_wuser(int_desc_5_wuser_9_wuser)
	,.int_desc_5_wuser_10_wuser(int_desc_5_wuser_10_wuser)
	,.int_desc_5_wuser_11_wuser(int_desc_5_wuser_11_wuser)
	,.int_desc_5_wuser_12_wuser(int_desc_5_wuser_12_wuser)
	,.int_desc_5_wuser_13_wuser(int_desc_5_wuser_13_wuser)
	,.int_desc_5_wuser_14_wuser(int_desc_5_wuser_14_wuser)
	,.int_desc_5_wuser_15_wuser(int_desc_5_wuser_15_wuser)
	,.int_desc_6_txn_type_wr_strb(int_desc_6_txn_type_wr_strb)
	,.int_desc_6_txn_type_wr_rd(int_desc_6_txn_type_wr_rd)
	,.int_desc_6_attr_axregion(int_desc_6_attr_axregion)
	,.int_desc_6_attr_axqos(int_desc_6_attr_axqos)
	,.int_desc_6_attr_axprot(int_desc_6_attr_axprot)
	,.int_desc_6_attr_axcache(int_desc_6_attr_axcache)
	,.int_desc_6_attr_axlock(int_desc_6_attr_axlock)
	,.int_desc_6_attr_axburst(int_desc_6_attr_axburst)
	,.int_desc_6_axid_0_axid(int_desc_6_axid_0_axid)
	,.int_desc_6_axid_1_axid(int_desc_6_axid_1_axid)
	,.int_desc_6_axid_2_axid(int_desc_6_axid_2_axid)
	,.int_desc_6_axid_3_axid(int_desc_6_axid_3_axid)
	,.int_desc_6_axuser_0_axuser(int_desc_6_axuser_0_axuser)
	,.int_desc_6_axuser_1_axuser(int_desc_6_axuser_1_axuser)
	,.int_desc_6_axuser_2_axuser(int_desc_6_axuser_2_axuser)
	,.int_desc_6_axuser_3_axuser(int_desc_6_axuser_3_axuser)
	,.int_desc_6_axuser_4_axuser(int_desc_6_axuser_4_axuser)
	,.int_desc_6_axuser_5_axuser(int_desc_6_axuser_5_axuser)
	,.int_desc_6_axuser_6_axuser(int_desc_6_axuser_6_axuser)
	,.int_desc_6_axuser_7_axuser(int_desc_6_axuser_7_axuser)
	,.int_desc_6_axuser_8_axuser(int_desc_6_axuser_8_axuser)
	,.int_desc_6_axuser_9_axuser(int_desc_6_axuser_9_axuser)
	,.int_desc_6_axuser_10_axuser(int_desc_6_axuser_10_axuser)
	,.int_desc_6_axuser_11_axuser(int_desc_6_axuser_11_axuser)
	,.int_desc_6_axuser_12_axuser(int_desc_6_axuser_12_axuser)
	,.int_desc_6_axuser_13_axuser(int_desc_6_axuser_13_axuser)
	,.int_desc_6_axuser_14_axuser(int_desc_6_axuser_14_axuser)
	,.int_desc_6_axuser_15_axuser(int_desc_6_axuser_15_axuser)
	,.int_desc_6_size_txn_size(int_desc_6_size_txn_size)
	,.int_desc_6_axsize_axsize(int_desc_6_axsize_axsize)
	,.int_desc_6_axaddr_0_addr(int_desc_6_axaddr_0_addr)
	,.int_desc_6_axaddr_1_addr(int_desc_6_axaddr_1_addr)
	,.int_desc_6_axaddr_2_addr(int_desc_6_axaddr_2_addr)
	,.int_desc_6_axaddr_3_addr(int_desc_6_axaddr_3_addr)
	,.int_desc_6_data_offset_addr(int_desc_6_data_offset_addr)
	,.int_desc_6_wuser_0_wuser(int_desc_6_wuser_0_wuser)
	,.int_desc_6_wuser_1_wuser(int_desc_6_wuser_1_wuser)
	,.int_desc_6_wuser_2_wuser(int_desc_6_wuser_2_wuser)
	,.int_desc_6_wuser_3_wuser(int_desc_6_wuser_3_wuser)
	,.int_desc_6_wuser_4_wuser(int_desc_6_wuser_4_wuser)
	,.int_desc_6_wuser_5_wuser(int_desc_6_wuser_5_wuser)
	,.int_desc_6_wuser_6_wuser(int_desc_6_wuser_6_wuser)
	,.int_desc_6_wuser_7_wuser(int_desc_6_wuser_7_wuser)
	,.int_desc_6_wuser_8_wuser(int_desc_6_wuser_8_wuser)
	,.int_desc_6_wuser_9_wuser(int_desc_6_wuser_9_wuser)
	,.int_desc_6_wuser_10_wuser(int_desc_6_wuser_10_wuser)
	,.int_desc_6_wuser_11_wuser(int_desc_6_wuser_11_wuser)
	,.int_desc_6_wuser_12_wuser(int_desc_6_wuser_12_wuser)
	,.int_desc_6_wuser_13_wuser(int_desc_6_wuser_13_wuser)
	,.int_desc_6_wuser_14_wuser(int_desc_6_wuser_14_wuser)
	,.int_desc_6_wuser_15_wuser(int_desc_6_wuser_15_wuser)
	,.int_desc_7_txn_type_wr_strb(int_desc_7_txn_type_wr_strb)
	,.int_desc_7_txn_type_wr_rd(int_desc_7_txn_type_wr_rd)
	,.int_desc_7_attr_axregion(int_desc_7_attr_axregion)
	,.int_desc_7_attr_axqos(int_desc_7_attr_axqos)
	,.int_desc_7_attr_axprot(int_desc_7_attr_axprot)
	,.int_desc_7_attr_axcache(int_desc_7_attr_axcache)
	,.int_desc_7_attr_axlock(int_desc_7_attr_axlock)
	,.int_desc_7_attr_axburst(int_desc_7_attr_axburst)
	,.int_desc_7_axid_0_axid(int_desc_7_axid_0_axid)
	,.int_desc_7_axid_1_axid(int_desc_7_axid_1_axid)
	,.int_desc_7_axid_2_axid(int_desc_7_axid_2_axid)
	,.int_desc_7_axid_3_axid(int_desc_7_axid_3_axid)
	,.int_desc_7_axuser_0_axuser(int_desc_7_axuser_0_axuser)
	,.int_desc_7_axuser_1_axuser(int_desc_7_axuser_1_axuser)
	,.int_desc_7_axuser_2_axuser(int_desc_7_axuser_2_axuser)
	,.int_desc_7_axuser_3_axuser(int_desc_7_axuser_3_axuser)
	,.int_desc_7_axuser_4_axuser(int_desc_7_axuser_4_axuser)
	,.int_desc_7_axuser_5_axuser(int_desc_7_axuser_5_axuser)
	,.int_desc_7_axuser_6_axuser(int_desc_7_axuser_6_axuser)
	,.int_desc_7_axuser_7_axuser(int_desc_7_axuser_7_axuser)
	,.int_desc_7_axuser_8_axuser(int_desc_7_axuser_8_axuser)
	,.int_desc_7_axuser_9_axuser(int_desc_7_axuser_9_axuser)
	,.int_desc_7_axuser_10_axuser(int_desc_7_axuser_10_axuser)
	,.int_desc_7_axuser_11_axuser(int_desc_7_axuser_11_axuser)
	,.int_desc_7_axuser_12_axuser(int_desc_7_axuser_12_axuser)
	,.int_desc_7_axuser_13_axuser(int_desc_7_axuser_13_axuser)
	,.int_desc_7_axuser_14_axuser(int_desc_7_axuser_14_axuser)
	,.int_desc_7_axuser_15_axuser(int_desc_7_axuser_15_axuser)
	,.int_desc_7_size_txn_size(int_desc_7_size_txn_size)
	,.int_desc_7_axsize_axsize(int_desc_7_axsize_axsize)
	,.int_desc_7_axaddr_0_addr(int_desc_7_axaddr_0_addr)
	,.int_desc_7_axaddr_1_addr(int_desc_7_axaddr_1_addr)
	,.int_desc_7_axaddr_2_addr(int_desc_7_axaddr_2_addr)
	,.int_desc_7_axaddr_3_addr(int_desc_7_axaddr_3_addr)
	,.int_desc_7_data_offset_addr(int_desc_7_data_offset_addr)
	,.int_desc_7_wuser_0_wuser(int_desc_7_wuser_0_wuser)
	,.int_desc_7_wuser_1_wuser(int_desc_7_wuser_1_wuser)
	,.int_desc_7_wuser_2_wuser(int_desc_7_wuser_2_wuser)
	,.int_desc_7_wuser_3_wuser(int_desc_7_wuser_3_wuser)
	,.int_desc_7_wuser_4_wuser(int_desc_7_wuser_4_wuser)
	,.int_desc_7_wuser_5_wuser(int_desc_7_wuser_5_wuser)
	,.int_desc_7_wuser_6_wuser(int_desc_7_wuser_6_wuser)
	,.int_desc_7_wuser_7_wuser(int_desc_7_wuser_7_wuser)
	,.int_desc_7_wuser_8_wuser(int_desc_7_wuser_8_wuser)
	,.int_desc_7_wuser_9_wuser(int_desc_7_wuser_9_wuser)
	,.int_desc_7_wuser_10_wuser(int_desc_7_wuser_10_wuser)
	,.int_desc_7_wuser_11_wuser(int_desc_7_wuser_11_wuser)
	,.int_desc_7_wuser_12_wuser(int_desc_7_wuser_12_wuser)
	,.int_desc_7_wuser_13_wuser(int_desc_7_wuser_13_wuser)
	,.int_desc_7_wuser_14_wuser(int_desc_7_wuser_14_wuser)
	,.int_desc_7_wuser_15_wuser(int_desc_7_wuser_15_wuser)
	,.int_desc_8_txn_type_wr_strb(int_desc_8_txn_type_wr_strb)
	,.int_desc_8_txn_type_wr_rd(int_desc_8_txn_type_wr_rd)
	,.int_desc_8_attr_axregion(int_desc_8_attr_axregion)
	,.int_desc_8_attr_axqos(int_desc_8_attr_axqos)
	,.int_desc_8_attr_axprot(int_desc_8_attr_axprot)
	,.int_desc_8_attr_axcache(int_desc_8_attr_axcache)
	,.int_desc_8_attr_axlock(int_desc_8_attr_axlock)
	,.int_desc_8_attr_axburst(int_desc_8_attr_axburst)
	,.int_desc_8_axid_0_axid(int_desc_8_axid_0_axid)
	,.int_desc_8_axid_1_axid(int_desc_8_axid_1_axid)
	,.int_desc_8_axid_2_axid(int_desc_8_axid_2_axid)
	,.int_desc_8_axid_3_axid(int_desc_8_axid_3_axid)
	,.int_desc_8_axuser_0_axuser(int_desc_8_axuser_0_axuser)
	,.int_desc_8_axuser_1_axuser(int_desc_8_axuser_1_axuser)
	,.int_desc_8_axuser_2_axuser(int_desc_8_axuser_2_axuser)
	,.int_desc_8_axuser_3_axuser(int_desc_8_axuser_3_axuser)
	,.int_desc_8_axuser_4_axuser(int_desc_8_axuser_4_axuser)
	,.int_desc_8_axuser_5_axuser(int_desc_8_axuser_5_axuser)
	,.int_desc_8_axuser_6_axuser(int_desc_8_axuser_6_axuser)
	,.int_desc_8_axuser_7_axuser(int_desc_8_axuser_7_axuser)
	,.int_desc_8_axuser_8_axuser(int_desc_8_axuser_8_axuser)
	,.int_desc_8_axuser_9_axuser(int_desc_8_axuser_9_axuser)
	,.int_desc_8_axuser_10_axuser(int_desc_8_axuser_10_axuser)
	,.int_desc_8_axuser_11_axuser(int_desc_8_axuser_11_axuser)
	,.int_desc_8_axuser_12_axuser(int_desc_8_axuser_12_axuser)
	,.int_desc_8_axuser_13_axuser(int_desc_8_axuser_13_axuser)
	,.int_desc_8_axuser_14_axuser(int_desc_8_axuser_14_axuser)
	,.int_desc_8_axuser_15_axuser(int_desc_8_axuser_15_axuser)
	,.int_desc_8_size_txn_size(int_desc_8_size_txn_size)
	,.int_desc_8_axsize_axsize(int_desc_8_axsize_axsize)
	,.int_desc_8_axaddr_0_addr(int_desc_8_axaddr_0_addr)
	,.int_desc_8_axaddr_1_addr(int_desc_8_axaddr_1_addr)
	,.int_desc_8_axaddr_2_addr(int_desc_8_axaddr_2_addr)
	,.int_desc_8_axaddr_3_addr(int_desc_8_axaddr_3_addr)
	,.int_desc_8_data_offset_addr(int_desc_8_data_offset_addr)
	,.int_desc_8_wuser_0_wuser(int_desc_8_wuser_0_wuser)
	,.int_desc_8_wuser_1_wuser(int_desc_8_wuser_1_wuser)
	,.int_desc_8_wuser_2_wuser(int_desc_8_wuser_2_wuser)
	,.int_desc_8_wuser_3_wuser(int_desc_8_wuser_3_wuser)
	,.int_desc_8_wuser_4_wuser(int_desc_8_wuser_4_wuser)
	,.int_desc_8_wuser_5_wuser(int_desc_8_wuser_5_wuser)
	,.int_desc_8_wuser_6_wuser(int_desc_8_wuser_6_wuser)
	,.int_desc_8_wuser_7_wuser(int_desc_8_wuser_7_wuser)
	,.int_desc_8_wuser_8_wuser(int_desc_8_wuser_8_wuser)
	,.int_desc_8_wuser_9_wuser(int_desc_8_wuser_9_wuser)
	,.int_desc_8_wuser_10_wuser(int_desc_8_wuser_10_wuser)
	,.int_desc_8_wuser_11_wuser(int_desc_8_wuser_11_wuser)
	,.int_desc_8_wuser_12_wuser(int_desc_8_wuser_12_wuser)
	,.int_desc_8_wuser_13_wuser(int_desc_8_wuser_13_wuser)
	,.int_desc_8_wuser_14_wuser(int_desc_8_wuser_14_wuser)
	,.int_desc_8_wuser_15_wuser(int_desc_8_wuser_15_wuser)
	,.int_desc_9_txn_type_wr_strb(int_desc_9_txn_type_wr_strb)
	,.int_desc_9_txn_type_wr_rd(int_desc_9_txn_type_wr_rd)
	,.int_desc_9_attr_axregion(int_desc_9_attr_axregion)
	,.int_desc_9_attr_axqos(int_desc_9_attr_axqos)
	,.int_desc_9_attr_axprot(int_desc_9_attr_axprot)
	,.int_desc_9_attr_axcache(int_desc_9_attr_axcache)
	,.int_desc_9_attr_axlock(int_desc_9_attr_axlock)
	,.int_desc_9_attr_axburst(int_desc_9_attr_axburst)
	,.int_desc_9_axid_0_axid(int_desc_9_axid_0_axid)
	,.int_desc_9_axid_1_axid(int_desc_9_axid_1_axid)
	,.int_desc_9_axid_2_axid(int_desc_9_axid_2_axid)
	,.int_desc_9_axid_3_axid(int_desc_9_axid_3_axid)
	,.int_desc_9_axuser_0_axuser(int_desc_9_axuser_0_axuser)
	,.int_desc_9_axuser_1_axuser(int_desc_9_axuser_1_axuser)
	,.int_desc_9_axuser_2_axuser(int_desc_9_axuser_2_axuser)
	,.int_desc_9_axuser_3_axuser(int_desc_9_axuser_3_axuser)
	,.int_desc_9_axuser_4_axuser(int_desc_9_axuser_4_axuser)
	,.int_desc_9_axuser_5_axuser(int_desc_9_axuser_5_axuser)
	,.int_desc_9_axuser_6_axuser(int_desc_9_axuser_6_axuser)
	,.int_desc_9_axuser_7_axuser(int_desc_9_axuser_7_axuser)
	,.int_desc_9_axuser_8_axuser(int_desc_9_axuser_8_axuser)
	,.int_desc_9_axuser_9_axuser(int_desc_9_axuser_9_axuser)
	,.int_desc_9_axuser_10_axuser(int_desc_9_axuser_10_axuser)
	,.int_desc_9_axuser_11_axuser(int_desc_9_axuser_11_axuser)
	,.int_desc_9_axuser_12_axuser(int_desc_9_axuser_12_axuser)
	,.int_desc_9_axuser_13_axuser(int_desc_9_axuser_13_axuser)
	,.int_desc_9_axuser_14_axuser(int_desc_9_axuser_14_axuser)
	,.int_desc_9_axuser_15_axuser(int_desc_9_axuser_15_axuser)
	,.int_desc_9_size_txn_size(int_desc_9_size_txn_size)
	,.int_desc_9_axsize_axsize(int_desc_9_axsize_axsize)
	,.int_desc_9_axaddr_0_addr(int_desc_9_axaddr_0_addr)
	,.int_desc_9_axaddr_1_addr(int_desc_9_axaddr_1_addr)
	,.int_desc_9_axaddr_2_addr(int_desc_9_axaddr_2_addr)
	,.int_desc_9_axaddr_3_addr(int_desc_9_axaddr_3_addr)
	,.int_desc_9_data_offset_addr(int_desc_9_data_offset_addr)
	,.int_desc_9_wuser_0_wuser(int_desc_9_wuser_0_wuser)
	,.int_desc_9_wuser_1_wuser(int_desc_9_wuser_1_wuser)
	,.int_desc_9_wuser_2_wuser(int_desc_9_wuser_2_wuser)
	,.int_desc_9_wuser_3_wuser(int_desc_9_wuser_3_wuser)
	,.int_desc_9_wuser_4_wuser(int_desc_9_wuser_4_wuser)
	,.int_desc_9_wuser_5_wuser(int_desc_9_wuser_5_wuser)
	,.int_desc_9_wuser_6_wuser(int_desc_9_wuser_6_wuser)
	,.int_desc_9_wuser_7_wuser(int_desc_9_wuser_7_wuser)
	,.int_desc_9_wuser_8_wuser(int_desc_9_wuser_8_wuser)
	,.int_desc_9_wuser_9_wuser(int_desc_9_wuser_9_wuser)
	,.int_desc_9_wuser_10_wuser(int_desc_9_wuser_10_wuser)
	,.int_desc_9_wuser_11_wuser(int_desc_9_wuser_11_wuser)
	,.int_desc_9_wuser_12_wuser(int_desc_9_wuser_12_wuser)
	,.int_desc_9_wuser_13_wuser(int_desc_9_wuser_13_wuser)
	,.int_desc_9_wuser_14_wuser(int_desc_9_wuser_14_wuser)
	,.int_desc_9_wuser_15_wuser(int_desc_9_wuser_15_wuser)
	,.int_desc_10_txn_type_wr_strb(int_desc_10_txn_type_wr_strb)
	,.int_desc_10_txn_type_wr_rd(int_desc_10_txn_type_wr_rd)
	,.int_desc_10_attr_axregion(int_desc_10_attr_axregion)
	,.int_desc_10_attr_axqos(int_desc_10_attr_axqos)
	,.int_desc_10_attr_axprot(int_desc_10_attr_axprot)
	,.int_desc_10_attr_axcache(int_desc_10_attr_axcache)
	,.int_desc_10_attr_axlock(int_desc_10_attr_axlock)
	,.int_desc_10_attr_axburst(int_desc_10_attr_axburst)
	,.int_desc_10_axid_0_axid(int_desc_10_axid_0_axid)
	,.int_desc_10_axid_1_axid(int_desc_10_axid_1_axid)
	,.int_desc_10_axid_2_axid(int_desc_10_axid_2_axid)
	,.int_desc_10_axid_3_axid(int_desc_10_axid_3_axid)
	,.int_desc_10_axuser_0_axuser(int_desc_10_axuser_0_axuser)
	,.int_desc_10_axuser_1_axuser(int_desc_10_axuser_1_axuser)
	,.int_desc_10_axuser_2_axuser(int_desc_10_axuser_2_axuser)
	,.int_desc_10_axuser_3_axuser(int_desc_10_axuser_3_axuser)
	,.int_desc_10_axuser_4_axuser(int_desc_10_axuser_4_axuser)
	,.int_desc_10_axuser_5_axuser(int_desc_10_axuser_5_axuser)
	,.int_desc_10_axuser_6_axuser(int_desc_10_axuser_6_axuser)
	,.int_desc_10_axuser_7_axuser(int_desc_10_axuser_7_axuser)
	,.int_desc_10_axuser_8_axuser(int_desc_10_axuser_8_axuser)
	,.int_desc_10_axuser_9_axuser(int_desc_10_axuser_9_axuser)
	,.int_desc_10_axuser_10_axuser(int_desc_10_axuser_10_axuser)
	,.int_desc_10_axuser_11_axuser(int_desc_10_axuser_11_axuser)
	,.int_desc_10_axuser_12_axuser(int_desc_10_axuser_12_axuser)
	,.int_desc_10_axuser_13_axuser(int_desc_10_axuser_13_axuser)
	,.int_desc_10_axuser_14_axuser(int_desc_10_axuser_14_axuser)
	,.int_desc_10_axuser_15_axuser(int_desc_10_axuser_15_axuser)
	,.int_desc_10_size_txn_size(int_desc_10_size_txn_size)
	,.int_desc_10_axsize_axsize(int_desc_10_axsize_axsize)
	,.int_desc_10_axaddr_0_addr(int_desc_10_axaddr_0_addr)
	,.int_desc_10_axaddr_1_addr(int_desc_10_axaddr_1_addr)
	,.int_desc_10_axaddr_2_addr(int_desc_10_axaddr_2_addr)
	,.int_desc_10_axaddr_3_addr(int_desc_10_axaddr_3_addr)
	,.int_desc_10_data_offset_addr(int_desc_10_data_offset_addr)
	,.int_desc_10_wuser_0_wuser(int_desc_10_wuser_0_wuser)
	,.int_desc_10_wuser_1_wuser(int_desc_10_wuser_1_wuser)
	,.int_desc_10_wuser_2_wuser(int_desc_10_wuser_2_wuser)
	,.int_desc_10_wuser_3_wuser(int_desc_10_wuser_3_wuser)
	,.int_desc_10_wuser_4_wuser(int_desc_10_wuser_4_wuser)
	,.int_desc_10_wuser_5_wuser(int_desc_10_wuser_5_wuser)
	,.int_desc_10_wuser_6_wuser(int_desc_10_wuser_6_wuser)
	,.int_desc_10_wuser_7_wuser(int_desc_10_wuser_7_wuser)
	,.int_desc_10_wuser_8_wuser(int_desc_10_wuser_8_wuser)
	,.int_desc_10_wuser_9_wuser(int_desc_10_wuser_9_wuser)
	,.int_desc_10_wuser_10_wuser(int_desc_10_wuser_10_wuser)
	,.int_desc_10_wuser_11_wuser(int_desc_10_wuser_11_wuser)
	,.int_desc_10_wuser_12_wuser(int_desc_10_wuser_12_wuser)
	,.int_desc_10_wuser_13_wuser(int_desc_10_wuser_13_wuser)
	,.int_desc_10_wuser_14_wuser(int_desc_10_wuser_14_wuser)
	,.int_desc_10_wuser_15_wuser(int_desc_10_wuser_15_wuser)
	,.int_desc_11_txn_type_wr_strb(int_desc_11_txn_type_wr_strb)
	,.int_desc_11_txn_type_wr_rd(int_desc_11_txn_type_wr_rd)
	,.int_desc_11_attr_axregion(int_desc_11_attr_axregion)
	,.int_desc_11_attr_axqos(int_desc_11_attr_axqos)
	,.int_desc_11_attr_axprot(int_desc_11_attr_axprot)
	,.int_desc_11_attr_axcache(int_desc_11_attr_axcache)
	,.int_desc_11_attr_axlock(int_desc_11_attr_axlock)
	,.int_desc_11_attr_axburst(int_desc_11_attr_axburst)
	,.int_desc_11_axid_0_axid(int_desc_11_axid_0_axid)
	,.int_desc_11_axid_1_axid(int_desc_11_axid_1_axid)
	,.int_desc_11_axid_2_axid(int_desc_11_axid_2_axid)
	,.int_desc_11_axid_3_axid(int_desc_11_axid_3_axid)
	,.int_desc_11_axuser_0_axuser(int_desc_11_axuser_0_axuser)
	,.int_desc_11_axuser_1_axuser(int_desc_11_axuser_1_axuser)
	,.int_desc_11_axuser_2_axuser(int_desc_11_axuser_2_axuser)
	,.int_desc_11_axuser_3_axuser(int_desc_11_axuser_3_axuser)
	,.int_desc_11_axuser_4_axuser(int_desc_11_axuser_4_axuser)
	,.int_desc_11_axuser_5_axuser(int_desc_11_axuser_5_axuser)
	,.int_desc_11_axuser_6_axuser(int_desc_11_axuser_6_axuser)
	,.int_desc_11_axuser_7_axuser(int_desc_11_axuser_7_axuser)
	,.int_desc_11_axuser_8_axuser(int_desc_11_axuser_8_axuser)
	,.int_desc_11_axuser_9_axuser(int_desc_11_axuser_9_axuser)
	,.int_desc_11_axuser_10_axuser(int_desc_11_axuser_10_axuser)
	,.int_desc_11_axuser_11_axuser(int_desc_11_axuser_11_axuser)
	,.int_desc_11_axuser_12_axuser(int_desc_11_axuser_12_axuser)
	,.int_desc_11_axuser_13_axuser(int_desc_11_axuser_13_axuser)
	,.int_desc_11_axuser_14_axuser(int_desc_11_axuser_14_axuser)
	,.int_desc_11_axuser_15_axuser(int_desc_11_axuser_15_axuser)
	,.int_desc_11_size_txn_size(int_desc_11_size_txn_size)
	,.int_desc_11_axsize_axsize(int_desc_11_axsize_axsize)
	,.int_desc_11_axaddr_0_addr(int_desc_11_axaddr_0_addr)
	,.int_desc_11_axaddr_1_addr(int_desc_11_axaddr_1_addr)
	,.int_desc_11_axaddr_2_addr(int_desc_11_axaddr_2_addr)
	,.int_desc_11_axaddr_3_addr(int_desc_11_axaddr_3_addr)
	,.int_desc_11_data_offset_addr(int_desc_11_data_offset_addr)
	,.int_desc_11_wuser_0_wuser(int_desc_11_wuser_0_wuser)
	,.int_desc_11_wuser_1_wuser(int_desc_11_wuser_1_wuser)
	,.int_desc_11_wuser_2_wuser(int_desc_11_wuser_2_wuser)
	,.int_desc_11_wuser_3_wuser(int_desc_11_wuser_3_wuser)
	,.int_desc_11_wuser_4_wuser(int_desc_11_wuser_4_wuser)
	,.int_desc_11_wuser_5_wuser(int_desc_11_wuser_5_wuser)
	,.int_desc_11_wuser_6_wuser(int_desc_11_wuser_6_wuser)
	,.int_desc_11_wuser_7_wuser(int_desc_11_wuser_7_wuser)
	,.int_desc_11_wuser_8_wuser(int_desc_11_wuser_8_wuser)
	,.int_desc_11_wuser_9_wuser(int_desc_11_wuser_9_wuser)
	,.int_desc_11_wuser_10_wuser(int_desc_11_wuser_10_wuser)
	,.int_desc_11_wuser_11_wuser(int_desc_11_wuser_11_wuser)
	,.int_desc_11_wuser_12_wuser(int_desc_11_wuser_12_wuser)
	,.int_desc_11_wuser_13_wuser(int_desc_11_wuser_13_wuser)
	,.int_desc_11_wuser_14_wuser(int_desc_11_wuser_14_wuser)
	,.int_desc_11_wuser_15_wuser(int_desc_11_wuser_15_wuser)
	,.int_desc_12_txn_type_wr_strb(int_desc_12_txn_type_wr_strb)
	,.int_desc_12_txn_type_wr_rd(int_desc_12_txn_type_wr_rd)
	,.int_desc_12_attr_axregion(int_desc_12_attr_axregion)
	,.int_desc_12_attr_axqos(int_desc_12_attr_axqos)
	,.int_desc_12_attr_axprot(int_desc_12_attr_axprot)
	,.int_desc_12_attr_axcache(int_desc_12_attr_axcache)
	,.int_desc_12_attr_axlock(int_desc_12_attr_axlock)
	,.int_desc_12_attr_axburst(int_desc_12_attr_axburst)
	,.int_desc_12_axid_0_axid(int_desc_12_axid_0_axid)
	,.int_desc_12_axid_1_axid(int_desc_12_axid_1_axid)
	,.int_desc_12_axid_2_axid(int_desc_12_axid_2_axid)
	,.int_desc_12_axid_3_axid(int_desc_12_axid_3_axid)
	,.int_desc_12_axuser_0_axuser(int_desc_12_axuser_0_axuser)
	,.int_desc_12_axuser_1_axuser(int_desc_12_axuser_1_axuser)
	,.int_desc_12_axuser_2_axuser(int_desc_12_axuser_2_axuser)
	,.int_desc_12_axuser_3_axuser(int_desc_12_axuser_3_axuser)
	,.int_desc_12_axuser_4_axuser(int_desc_12_axuser_4_axuser)
	,.int_desc_12_axuser_5_axuser(int_desc_12_axuser_5_axuser)
	,.int_desc_12_axuser_6_axuser(int_desc_12_axuser_6_axuser)
	,.int_desc_12_axuser_7_axuser(int_desc_12_axuser_7_axuser)
	,.int_desc_12_axuser_8_axuser(int_desc_12_axuser_8_axuser)
	,.int_desc_12_axuser_9_axuser(int_desc_12_axuser_9_axuser)
	,.int_desc_12_axuser_10_axuser(int_desc_12_axuser_10_axuser)
	,.int_desc_12_axuser_11_axuser(int_desc_12_axuser_11_axuser)
	,.int_desc_12_axuser_12_axuser(int_desc_12_axuser_12_axuser)
	,.int_desc_12_axuser_13_axuser(int_desc_12_axuser_13_axuser)
	,.int_desc_12_axuser_14_axuser(int_desc_12_axuser_14_axuser)
	,.int_desc_12_axuser_15_axuser(int_desc_12_axuser_15_axuser)
	,.int_desc_12_size_txn_size(int_desc_12_size_txn_size)
	,.int_desc_12_axsize_axsize(int_desc_12_axsize_axsize)
	,.int_desc_12_axaddr_0_addr(int_desc_12_axaddr_0_addr)
	,.int_desc_12_axaddr_1_addr(int_desc_12_axaddr_1_addr)
	,.int_desc_12_axaddr_2_addr(int_desc_12_axaddr_2_addr)
	,.int_desc_12_axaddr_3_addr(int_desc_12_axaddr_3_addr)
	,.int_desc_12_data_offset_addr(int_desc_12_data_offset_addr)
	,.int_desc_12_wuser_0_wuser(int_desc_12_wuser_0_wuser)
	,.int_desc_12_wuser_1_wuser(int_desc_12_wuser_1_wuser)
	,.int_desc_12_wuser_2_wuser(int_desc_12_wuser_2_wuser)
	,.int_desc_12_wuser_3_wuser(int_desc_12_wuser_3_wuser)
	,.int_desc_12_wuser_4_wuser(int_desc_12_wuser_4_wuser)
	,.int_desc_12_wuser_5_wuser(int_desc_12_wuser_5_wuser)
	,.int_desc_12_wuser_6_wuser(int_desc_12_wuser_6_wuser)
	,.int_desc_12_wuser_7_wuser(int_desc_12_wuser_7_wuser)
	,.int_desc_12_wuser_8_wuser(int_desc_12_wuser_8_wuser)
	,.int_desc_12_wuser_9_wuser(int_desc_12_wuser_9_wuser)
	,.int_desc_12_wuser_10_wuser(int_desc_12_wuser_10_wuser)
	,.int_desc_12_wuser_11_wuser(int_desc_12_wuser_11_wuser)
	,.int_desc_12_wuser_12_wuser(int_desc_12_wuser_12_wuser)
	,.int_desc_12_wuser_13_wuser(int_desc_12_wuser_13_wuser)
	,.int_desc_12_wuser_14_wuser(int_desc_12_wuser_14_wuser)
	,.int_desc_12_wuser_15_wuser(int_desc_12_wuser_15_wuser)
	,.int_desc_13_txn_type_wr_strb(int_desc_13_txn_type_wr_strb)
	,.int_desc_13_txn_type_wr_rd(int_desc_13_txn_type_wr_rd)
	,.int_desc_13_attr_axregion(int_desc_13_attr_axregion)
	,.int_desc_13_attr_axqos(int_desc_13_attr_axqos)
	,.int_desc_13_attr_axprot(int_desc_13_attr_axprot)
	,.int_desc_13_attr_axcache(int_desc_13_attr_axcache)
	,.int_desc_13_attr_axlock(int_desc_13_attr_axlock)
	,.int_desc_13_attr_axburst(int_desc_13_attr_axburst)
	,.int_desc_13_axid_0_axid(int_desc_13_axid_0_axid)
	,.int_desc_13_axid_1_axid(int_desc_13_axid_1_axid)
	,.int_desc_13_axid_2_axid(int_desc_13_axid_2_axid)
	,.int_desc_13_axid_3_axid(int_desc_13_axid_3_axid)
	,.int_desc_13_axuser_0_axuser(int_desc_13_axuser_0_axuser)
	,.int_desc_13_axuser_1_axuser(int_desc_13_axuser_1_axuser)
	,.int_desc_13_axuser_2_axuser(int_desc_13_axuser_2_axuser)
	,.int_desc_13_axuser_3_axuser(int_desc_13_axuser_3_axuser)
	,.int_desc_13_axuser_4_axuser(int_desc_13_axuser_4_axuser)
	,.int_desc_13_axuser_5_axuser(int_desc_13_axuser_5_axuser)
	,.int_desc_13_axuser_6_axuser(int_desc_13_axuser_6_axuser)
	,.int_desc_13_axuser_7_axuser(int_desc_13_axuser_7_axuser)
	,.int_desc_13_axuser_8_axuser(int_desc_13_axuser_8_axuser)
	,.int_desc_13_axuser_9_axuser(int_desc_13_axuser_9_axuser)
	,.int_desc_13_axuser_10_axuser(int_desc_13_axuser_10_axuser)
	,.int_desc_13_axuser_11_axuser(int_desc_13_axuser_11_axuser)
	,.int_desc_13_axuser_12_axuser(int_desc_13_axuser_12_axuser)
	,.int_desc_13_axuser_13_axuser(int_desc_13_axuser_13_axuser)
	,.int_desc_13_axuser_14_axuser(int_desc_13_axuser_14_axuser)
	,.int_desc_13_axuser_15_axuser(int_desc_13_axuser_15_axuser)
	,.int_desc_13_size_txn_size(int_desc_13_size_txn_size)
	,.int_desc_13_axsize_axsize(int_desc_13_axsize_axsize)
	,.int_desc_13_axaddr_0_addr(int_desc_13_axaddr_0_addr)
	,.int_desc_13_axaddr_1_addr(int_desc_13_axaddr_1_addr)
	,.int_desc_13_axaddr_2_addr(int_desc_13_axaddr_2_addr)
	,.int_desc_13_axaddr_3_addr(int_desc_13_axaddr_3_addr)
	,.int_desc_13_data_offset_addr(int_desc_13_data_offset_addr)
	,.int_desc_13_wuser_0_wuser(int_desc_13_wuser_0_wuser)
	,.int_desc_13_wuser_1_wuser(int_desc_13_wuser_1_wuser)
	,.int_desc_13_wuser_2_wuser(int_desc_13_wuser_2_wuser)
	,.int_desc_13_wuser_3_wuser(int_desc_13_wuser_3_wuser)
	,.int_desc_13_wuser_4_wuser(int_desc_13_wuser_4_wuser)
	,.int_desc_13_wuser_5_wuser(int_desc_13_wuser_5_wuser)
	,.int_desc_13_wuser_6_wuser(int_desc_13_wuser_6_wuser)
	,.int_desc_13_wuser_7_wuser(int_desc_13_wuser_7_wuser)
	,.int_desc_13_wuser_8_wuser(int_desc_13_wuser_8_wuser)
	,.int_desc_13_wuser_9_wuser(int_desc_13_wuser_9_wuser)
	,.int_desc_13_wuser_10_wuser(int_desc_13_wuser_10_wuser)
	,.int_desc_13_wuser_11_wuser(int_desc_13_wuser_11_wuser)
	,.int_desc_13_wuser_12_wuser(int_desc_13_wuser_12_wuser)
	,.int_desc_13_wuser_13_wuser(int_desc_13_wuser_13_wuser)
	,.int_desc_13_wuser_14_wuser(int_desc_13_wuser_14_wuser)
	,.int_desc_13_wuser_15_wuser(int_desc_13_wuser_15_wuser)
	,.int_desc_14_txn_type_wr_strb(int_desc_14_txn_type_wr_strb)
	,.int_desc_14_txn_type_wr_rd(int_desc_14_txn_type_wr_rd)
	,.int_desc_14_attr_axregion(int_desc_14_attr_axregion)
	,.int_desc_14_attr_axqos(int_desc_14_attr_axqos)
	,.int_desc_14_attr_axprot(int_desc_14_attr_axprot)
	,.int_desc_14_attr_axcache(int_desc_14_attr_axcache)
	,.int_desc_14_attr_axlock(int_desc_14_attr_axlock)
	,.int_desc_14_attr_axburst(int_desc_14_attr_axburst)
	,.int_desc_14_axid_0_axid(int_desc_14_axid_0_axid)
	,.int_desc_14_axid_1_axid(int_desc_14_axid_1_axid)
	,.int_desc_14_axid_2_axid(int_desc_14_axid_2_axid)
	,.int_desc_14_axid_3_axid(int_desc_14_axid_3_axid)
	,.int_desc_14_axuser_0_axuser(int_desc_14_axuser_0_axuser)
	,.int_desc_14_axuser_1_axuser(int_desc_14_axuser_1_axuser)
	,.int_desc_14_axuser_2_axuser(int_desc_14_axuser_2_axuser)
	,.int_desc_14_axuser_3_axuser(int_desc_14_axuser_3_axuser)
	,.int_desc_14_axuser_4_axuser(int_desc_14_axuser_4_axuser)
	,.int_desc_14_axuser_5_axuser(int_desc_14_axuser_5_axuser)
	,.int_desc_14_axuser_6_axuser(int_desc_14_axuser_6_axuser)
	,.int_desc_14_axuser_7_axuser(int_desc_14_axuser_7_axuser)
	,.int_desc_14_axuser_8_axuser(int_desc_14_axuser_8_axuser)
	,.int_desc_14_axuser_9_axuser(int_desc_14_axuser_9_axuser)
	,.int_desc_14_axuser_10_axuser(int_desc_14_axuser_10_axuser)
	,.int_desc_14_axuser_11_axuser(int_desc_14_axuser_11_axuser)
	,.int_desc_14_axuser_12_axuser(int_desc_14_axuser_12_axuser)
	,.int_desc_14_axuser_13_axuser(int_desc_14_axuser_13_axuser)
	,.int_desc_14_axuser_14_axuser(int_desc_14_axuser_14_axuser)
	,.int_desc_14_axuser_15_axuser(int_desc_14_axuser_15_axuser)
	,.int_desc_14_size_txn_size(int_desc_14_size_txn_size)
	,.int_desc_14_axsize_axsize(int_desc_14_axsize_axsize)
	,.int_desc_14_axaddr_0_addr(int_desc_14_axaddr_0_addr)
	,.int_desc_14_axaddr_1_addr(int_desc_14_axaddr_1_addr)
	,.int_desc_14_axaddr_2_addr(int_desc_14_axaddr_2_addr)
	,.int_desc_14_axaddr_3_addr(int_desc_14_axaddr_3_addr)
	,.int_desc_14_data_offset_addr(int_desc_14_data_offset_addr)
	,.int_desc_14_wuser_0_wuser(int_desc_14_wuser_0_wuser)
	,.int_desc_14_wuser_1_wuser(int_desc_14_wuser_1_wuser)
	,.int_desc_14_wuser_2_wuser(int_desc_14_wuser_2_wuser)
	,.int_desc_14_wuser_3_wuser(int_desc_14_wuser_3_wuser)
	,.int_desc_14_wuser_4_wuser(int_desc_14_wuser_4_wuser)
	,.int_desc_14_wuser_5_wuser(int_desc_14_wuser_5_wuser)
	,.int_desc_14_wuser_6_wuser(int_desc_14_wuser_6_wuser)
	,.int_desc_14_wuser_7_wuser(int_desc_14_wuser_7_wuser)
	,.int_desc_14_wuser_8_wuser(int_desc_14_wuser_8_wuser)
	,.int_desc_14_wuser_9_wuser(int_desc_14_wuser_9_wuser)
	,.int_desc_14_wuser_10_wuser(int_desc_14_wuser_10_wuser)
	,.int_desc_14_wuser_11_wuser(int_desc_14_wuser_11_wuser)
	,.int_desc_14_wuser_12_wuser(int_desc_14_wuser_12_wuser)
	,.int_desc_14_wuser_13_wuser(int_desc_14_wuser_13_wuser)
	,.int_desc_14_wuser_14_wuser(int_desc_14_wuser_14_wuser)
	,.int_desc_14_wuser_15_wuser(int_desc_14_wuser_15_wuser)
	,.int_desc_15_txn_type_wr_strb(int_desc_15_txn_type_wr_strb)
	,.int_desc_15_txn_type_wr_rd(int_desc_15_txn_type_wr_rd)
	,.int_desc_15_attr_axregion(int_desc_15_attr_axregion)
	,.int_desc_15_attr_axqos(int_desc_15_attr_axqos)
	,.int_desc_15_attr_axprot(int_desc_15_attr_axprot)
	,.int_desc_15_attr_axcache(int_desc_15_attr_axcache)
	,.int_desc_15_attr_axlock(int_desc_15_attr_axlock)
	,.int_desc_15_attr_axburst(int_desc_15_attr_axburst)
	,.int_desc_15_axid_0_axid(int_desc_15_axid_0_axid)
	,.int_desc_15_axid_1_axid(int_desc_15_axid_1_axid)
	,.int_desc_15_axid_2_axid(int_desc_15_axid_2_axid)
	,.int_desc_15_axid_3_axid(int_desc_15_axid_3_axid)
	,.int_desc_15_axuser_0_axuser(int_desc_15_axuser_0_axuser)
	,.int_desc_15_axuser_1_axuser(int_desc_15_axuser_1_axuser)
	,.int_desc_15_axuser_2_axuser(int_desc_15_axuser_2_axuser)
	,.int_desc_15_axuser_3_axuser(int_desc_15_axuser_3_axuser)
	,.int_desc_15_axuser_4_axuser(int_desc_15_axuser_4_axuser)
	,.int_desc_15_axuser_5_axuser(int_desc_15_axuser_5_axuser)
	,.int_desc_15_axuser_6_axuser(int_desc_15_axuser_6_axuser)
	,.int_desc_15_axuser_7_axuser(int_desc_15_axuser_7_axuser)
	,.int_desc_15_axuser_8_axuser(int_desc_15_axuser_8_axuser)
	,.int_desc_15_axuser_9_axuser(int_desc_15_axuser_9_axuser)
	,.int_desc_15_axuser_10_axuser(int_desc_15_axuser_10_axuser)
	,.int_desc_15_axuser_11_axuser(int_desc_15_axuser_11_axuser)
	,.int_desc_15_axuser_12_axuser(int_desc_15_axuser_12_axuser)
	,.int_desc_15_axuser_13_axuser(int_desc_15_axuser_13_axuser)
	,.int_desc_15_axuser_14_axuser(int_desc_15_axuser_14_axuser)
	,.int_desc_15_axuser_15_axuser(int_desc_15_axuser_15_axuser)
	,.int_desc_15_size_txn_size(int_desc_15_size_txn_size)
	,.int_desc_15_axsize_axsize(int_desc_15_axsize_axsize)
	,.int_desc_15_axaddr_0_addr(int_desc_15_axaddr_0_addr)
	,.int_desc_15_axaddr_1_addr(int_desc_15_axaddr_1_addr)
	,.int_desc_15_axaddr_2_addr(int_desc_15_axaddr_2_addr)
	,.int_desc_15_axaddr_3_addr(int_desc_15_axaddr_3_addr)
	,.int_desc_15_data_offset_addr(int_desc_15_data_offset_addr)
	,.int_desc_15_wuser_0_wuser(int_desc_15_wuser_0_wuser)
	,.int_desc_15_wuser_1_wuser(int_desc_15_wuser_1_wuser)
	,.int_desc_15_wuser_2_wuser(int_desc_15_wuser_2_wuser)
	,.int_desc_15_wuser_3_wuser(int_desc_15_wuser_3_wuser)
	,.int_desc_15_wuser_4_wuser(int_desc_15_wuser_4_wuser)
	,.int_desc_15_wuser_5_wuser(int_desc_15_wuser_5_wuser)
	,.int_desc_15_wuser_6_wuser(int_desc_15_wuser_6_wuser)
	,.int_desc_15_wuser_7_wuser(int_desc_15_wuser_7_wuser)
	,.int_desc_15_wuser_8_wuser(int_desc_15_wuser_8_wuser)
	,.int_desc_15_wuser_9_wuser(int_desc_15_wuser_9_wuser)
	,.int_desc_15_wuser_10_wuser(int_desc_15_wuser_10_wuser)
	,.int_desc_15_wuser_11_wuser(int_desc_15_wuser_11_wuser)
	,.int_desc_15_wuser_12_wuser(int_desc_15_wuser_12_wuser)
	,.int_desc_15_wuser_13_wuser(int_desc_15_wuser_13_wuser)
	,.int_desc_15_wuser_14_wuser(int_desc_15_wuser_14_wuser)
	,.int_desc_15_wuser_15_wuser(int_desc_15_wuser_15_wuser)
	,.uc2rb_rd_addr(uc2rb_rd_addr)
	,.uc2rb_wr_we(uc2rb_wr_we)
	,.uc2rb_wr_bwe(uc2rb_wr_bwe)
	,.uc2rb_wr_addr(uc2rb_wr_addr)
	,.uc2rb_wr_data(uc2rb_wr_data   )
	,.uc2rb_wr_wstrb(uc2rb_wr_wstrb   )
	,.uc2hm_trig(uc2hm_trig)
	,.int_version_major_ver(int_version_major_ver)
	,.int_version_minor_ver(int_version_minor_ver)
	,.int_bridge_type_type(int_bridge_type_type)
	,.int_axi_bridge_config_user_width(int_axi_bridge_config_user_width)
	,.int_axi_bridge_config_id_width(int_axi_bridge_config_id_width)
	,.int_axi_bridge_config_data_width(int_axi_bridge_config_data_width)
	,.int_reset_dut_srst_3(int_reset_dut_srst_3)
	,.int_reset_dut_srst_2(int_reset_dut_srst_2)
	,.int_reset_dut_srst_1(int_reset_dut_srst_1)
	,.int_reset_dut_srst_0(int_reset_dut_srst_0)
	,.int_reset_srst(int_reset_srst)
	,.int_mode_select_imm_bresp(int_mode_select_imm_bresp)
	,.int_mode_select_mode_2(int_mode_select_mode_2)
	,.int_mode_select_mode_0_1(int_mode_select_mode_0_1)
	,.int_ownership_flip_flip(int_ownership_flip_flip)
	,.int_status_resp_comp_resp_comp(int_status_resp_comp_resp_comp)
	,.int_status_resp_resp(int_status_resp_resp)
	,.int_intr_status_comp(int_intr_status_comp)
	,.int_intr_status_c2h(int_intr_status_c2h)
	,.int_intr_status_error(int_intr_status_error)
	,.int_intr_status_txn_avail(int_intr_status_txn_avail)
	,.int_intr_txn_avail_clear_clr_avail(int_intr_txn_avail_clear_clr_avail)
	,.int_intr_txn_avail_enable_en_avail(int_intr_txn_avail_enable_en_avail)
	,.int_intr_comp_clear_clr_comp(int_intr_comp_clear_clr_comp)
	,.int_intr_comp_enable_en_comp(int_intr_comp_enable_en_comp)
	,.int_intr_error_status_err_2(int_intr_error_status_err_2)
	,.int_intr_error_status_err_1(int_intr_error_status_err_1)
	,.int_intr_error_clear_clr_err_2(int_intr_error_clear_clr_err_2)
	,.int_intr_error_clear_clr_err_1(int_intr_error_clear_clr_err_1)
	,.int_intr_error_clear_clr_err_0(int_intr_error_clear_clr_err_0)
	,.int_intr_error_enable_en_err_2(int_intr_error_enable_en_err_2)
	,.int_intr_error_enable_en_err_1(int_intr_error_enable_en_err_1)
	,.int_intr_error_enable_en_err_0(int_intr_error_enable_en_err_0)
	,.int_intr_h2c_0_h2c(int_intr_h2c_0_h2c)
	,.int_intr_h2c_1_h2c(int_intr_h2c_1_h2c)
	,.int_intr_c2h_0_status_c2h(int_intr_c2h_0_status_c2h)
	,.int_intr_c2h_1_status_c2h(int_intr_c2h_1_status_c2h)
	,.int_c2h_gpio_0_status_gpio(int_c2h_gpio_0_status_gpio)
	,.int_c2h_gpio_1_status_gpio(int_c2h_gpio_1_status_gpio)
	,.int_c2h_gpio_2_status_gpio(int_c2h_gpio_2_status_gpio)
	,.int_c2h_gpio_3_status_gpio(int_c2h_gpio_3_status_gpio)
	,.int_c2h_gpio_4_status_gpio(int_c2h_gpio_4_status_gpio)
	,.int_c2h_gpio_5_status_gpio(int_c2h_gpio_5_status_gpio)
	,.int_c2h_gpio_6_status_gpio(int_c2h_gpio_6_status_gpio)
	,.int_c2h_gpio_7_status_gpio(int_c2h_gpio_7_status_gpio)
	,.int_c2h_gpio_8_status_gpio(int_c2h_gpio_8_status_gpio)
	,.int_c2h_gpio_9_status_gpio(int_c2h_gpio_9_status_gpio)
	,.int_c2h_gpio_10_status_gpio(int_c2h_gpio_10_status_gpio)
	,.int_c2h_gpio_11_status_gpio(int_c2h_gpio_11_status_gpio)
	,.int_c2h_gpio_12_status_gpio(int_c2h_gpio_12_status_gpio)
	,.int_c2h_gpio_13_status_gpio(int_c2h_gpio_13_status_gpio)
	,.int_c2h_gpio_14_status_gpio(int_c2h_gpio_14_status_gpio)
	,.int_c2h_gpio_15_status_gpio(int_c2h_gpio_15_status_gpio)
	,.int_addr_in_0_addr(int_addr_in_0_addr)
	,.int_addr_in_1_addr(int_addr_in_1_addr)
	,.int_addr_in_2_addr(int_addr_in_2_addr)
	,.int_addr_in_3_addr(int_addr_in_3_addr)
	,.int_trans_mask_0_addr(int_trans_mask_0_addr)
	,.int_trans_mask_1_addr(int_trans_mask_1_addr)
	,.int_trans_mask_2_addr(int_trans_mask_2_addr)
	,.int_trans_mask_3_addr(int_trans_mask_3_addr)
	,.int_trans_addr_0_addr(int_trans_addr_0_addr)
	,.int_trans_addr_1_addr(int_trans_addr_1_addr)
	,.int_trans_addr_2_addr(int_trans_addr_2_addr)
	,.int_trans_addr_3_addr(int_trans_addr_3_addr)
	,.int_desc_0_data_host_addr_0_addr(int_desc_0_data_host_addr_0_addr)
	,.int_desc_0_data_host_addr_1_addr(int_desc_0_data_host_addr_1_addr)
	,.int_desc_0_data_host_addr_2_addr(int_desc_0_data_host_addr_2_addr)
	,.int_desc_0_data_host_addr_3_addr(int_desc_0_data_host_addr_3_addr)
	,.int_desc_0_wstrb_host_addr_0_addr(int_desc_0_wstrb_host_addr_0_addr)
	,.int_desc_0_wstrb_host_addr_1_addr(int_desc_0_wstrb_host_addr_1_addr)
	,.int_desc_0_wstrb_host_addr_2_addr(int_desc_0_wstrb_host_addr_2_addr)
	,.int_desc_0_wstrb_host_addr_3_addr(int_desc_0_wstrb_host_addr_3_addr)
	,.int_desc_1_data_host_addr_0_addr(int_desc_1_data_host_addr_0_addr)
	,.int_desc_1_data_host_addr_1_addr(int_desc_1_data_host_addr_1_addr)
	,.int_desc_1_data_host_addr_2_addr(int_desc_1_data_host_addr_2_addr)
	,.int_desc_1_data_host_addr_3_addr(int_desc_1_data_host_addr_3_addr)
	,.int_desc_1_wstrb_host_addr_0_addr(int_desc_1_wstrb_host_addr_0_addr)
	,.int_desc_1_wstrb_host_addr_1_addr(int_desc_1_wstrb_host_addr_1_addr)
	,.int_desc_1_wstrb_host_addr_2_addr(int_desc_1_wstrb_host_addr_2_addr)
	,.int_desc_1_wstrb_host_addr_3_addr(int_desc_1_wstrb_host_addr_3_addr)
	,.int_desc_2_data_host_addr_0_addr(int_desc_2_data_host_addr_0_addr)
	,.int_desc_2_data_host_addr_1_addr(int_desc_2_data_host_addr_1_addr)
	,.int_desc_2_data_host_addr_2_addr(int_desc_2_data_host_addr_2_addr)
	,.int_desc_2_data_host_addr_3_addr(int_desc_2_data_host_addr_3_addr)
	,.int_desc_2_wstrb_host_addr_0_addr(int_desc_2_wstrb_host_addr_0_addr)
	,.int_desc_2_wstrb_host_addr_1_addr(int_desc_2_wstrb_host_addr_1_addr)
	,.int_desc_2_wstrb_host_addr_2_addr(int_desc_2_wstrb_host_addr_2_addr)
	,.int_desc_2_wstrb_host_addr_3_addr(int_desc_2_wstrb_host_addr_3_addr)
	,.int_desc_3_data_host_addr_0_addr(int_desc_3_data_host_addr_0_addr)
	,.int_desc_3_data_host_addr_1_addr(int_desc_3_data_host_addr_1_addr)
	,.int_desc_3_data_host_addr_2_addr(int_desc_3_data_host_addr_2_addr)
	,.int_desc_3_data_host_addr_3_addr(int_desc_3_data_host_addr_3_addr)
	,.int_desc_3_wstrb_host_addr_0_addr(int_desc_3_wstrb_host_addr_0_addr)
	,.int_desc_3_wstrb_host_addr_1_addr(int_desc_3_wstrb_host_addr_1_addr)
	,.int_desc_3_wstrb_host_addr_2_addr(int_desc_3_wstrb_host_addr_2_addr)
	,.int_desc_3_wstrb_host_addr_3_addr(int_desc_3_wstrb_host_addr_3_addr)
	,.int_desc_4_data_host_addr_0_addr(int_desc_4_data_host_addr_0_addr)
	,.int_desc_4_data_host_addr_1_addr(int_desc_4_data_host_addr_1_addr)
	,.int_desc_4_data_host_addr_2_addr(int_desc_4_data_host_addr_2_addr)
	,.int_desc_4_data_host_addr_3_addr(int_desc_4_data_host_addr_3_addr)
	,.int_desc_4_wstrb_host_addr_0_addr(int_desc_4_wstrb_host_addr_0_addr)
	,.int_desc_4_wstrb_host_addr_1_addr(int_desc_4_wstrb_host_addr_1_addr)
	,.int_desc_4_wstrb_host_addr_2_addr(int_desc_4_wstrb_host_addr_2_addr)
	,.int_desc_4_wstrb_host_addr_3_addr(int_desc_4_wstrb_host_addr_3_addr)
	,.int_desc_5_data_host_addr_0_addr(int_desc_5_data_host_addr_0_addr)
	,.int_desc_5_data_host_addr_1_addr(int_desc_5_data_host_addr_1_addr)
	,.int_desc_5_data_host_addr_2_addr(int_desc_5_data_host_addr_2_addr)
	,.int_desc_5_data_host_addr_3_addr(int_desc_5_data_host_addr_3_addr)
	,.int_desc_5_wstrb_host_addr_0_addr(int_desc_5_wstrb_host_addr_0_addr)
	,.int_desc_5_wstrb_host_addr_1_addr(int_desc_5_wstrb_host_addr_1_addr)
	,.int_desc_5_wstrb_host_addr_2_addr(int_desc_5_wstrb_host_addr_2_addr)
	,.int_desc_5_wstrb_host_addr_3_addr(int_desc_5_wstrb_host_addr_3_addr)
	,.int_desc_6_data_host_addr_0_addr(int_desc_6_data_host_addr_0_addr)
	,.int_desc_6_data_host_addr_1_addr(int_desc_6_data_host_addr_1_addr)
	,.int_desc_6_data_host_addr_2_addr(int_desc_6_data_host_addr_2_addr)
	,.int_desc_6_data_host_addr_3_addr(int_desc_6_data_host_addr_3_addr)
	,.int_desc_6_wstrb_host_addr_0_addr(int_desc_6_wstrb_host_addr_0_addr)
	,.int_desc_6_wstrb_host_addr_1_addr(int_desc_6_wstrb_host_addr_1_addr)
	,.int_desc_6_wstrb_host_addr_2_addr(int_desc_6_wstrb_host_addr_2_addr)
	,.int_desc_6_wstrb_host_addr_3_addr(int_desc_6_wstrb_host_addr_3_addr)
	,.int_desc_7_data_host_addr_0_addr(int_desc_7_data_host_addr_0_addr)
	,.int_desc_7_data_host_addr_1_addr(int_desc_7_data_host_addr_1_addr)
	,.int_desc_7_data_host_addr_2_addr(int_desc_7_data_host_addr_2_addr)
	,.int_desc_7_data_host_addr_3_addr(int_desc_7_data_host_addr_3_addr)
	,.int_desc_7_wstrb_host_addr_0_addr(int_desc_7_wstrb_host_addr_0_addr)
	,.int_desc_7_wstrb_host_addr_1_addr(int_desc_7_wstrb_host_addr_1_addr)
	,.int_desc_7_wstrb_host_addr_2_addr(int_desc_7_wstrb_host_addr_2_addr)
	,.int_desc_7_wstrb_host_addr_3_addr(int_desc_7_wstrb_host_addr_3_addr)
	,.int_desc_8_data_host_addr_0_addr(int_desc_8_data_host_addr_0_addr)
	,.int_desc_8_data_host_addr_1_addr(int_desc_8_data_host_addr_1_addr)
	,.int_desc_8_data_host_addr_2_addr(int_desc_8_data_host_addr_2_addr)
	,.int_desc_8_data_host_addr_3_addr(int_desc_8_data_host_addr_3_addr)
	,.int_desc_8_wstrb_host_addr_0_addr(int_desc_8_wstrb_host_addr_0_addr)
	,.int_desc_8_wstrb_host_addr_1_addr(int_desc_8_wstrb_host_addr_1_addr)
	,.int_desc_8_wstrb_host_addr_2_addr(int_desc_8_wstrb_host_addr_2_addr)
	,.int_desc_8_wstrb_host_addr_3_addr(int_desc_8_wstrb_host_addr_3_addr)
	,.int_desc_9_data_host_addr_0_addr(int_desc_9_data_host_addr_0_addr)
	,.int_desc_9_data_host_addr_1_addr(int_desc_9_data_host_addr_1_addr)
	,.int_desc_9_data_host_addr_2_addr(int_desc_9_data_host_addr_2_addr)
	,.int_desc_9_data_host_addr_3_addr(int_desc_9_data_host_addr_3_addr)
	,.int_desc_9_wstrb_host_addr_0_addr(int_desc_9_wstrb_host_addr_0_addr)
	,.int_desc_9_wstrb_host_addr_1_addr(int_desc_9_wstrb_host_addr_1_addr)
	,.int_desc_9_wstrb_host_addr_2_addr(int_desc_9_wstrb_host_addr_2_addr)
	,.int_desc_9_wstrb_host_addr_3_addr(int_desc_9_wstrb_host_addr_3_addr)
	,.int_desc_10_data_host_addr_0_addr(int_desc_10_data_host_addr_0_addr)
	,.int_desc_10_data_host_addr_1_addr(int_desc_10_data_host_addr_1_addr)
	,.int_desc_10_data_host_addr_2_addr(int_desc_10_data_host_addr_2_addr)
	,.int_desc_10_data_host_addr_3_addr(int_desc_10_data_host_addr_3_addr)
	,.int_desc_10_wstrb_host_addr_0_addr(int_desc_10_wstrb_host_addr_0_addr)
	,.int_desc_10_wstrb_host_addr_1_addr(int_desc_10_wstrb_host_addr_1_addr)
	,.int_desc_10_wstrb_host_addr_2_addr(int_desc_10_wstrb_host_addr_2_addr)
	,.int_desc_10_wstrb_host_addr_3_addr(int_desc_10_wstrb_host_addr_3_addr)
	,.int_desc_11_data_host_addr_0_addr(int_desc_11_data_host_addr_0_addr)
	,.int_desc_11_data_host_addr_1_addr(int_desc_11_data_host_addr_1_addr)
	,.int_desc_11_data_host_addr_2_addr(int_desc_11_data_host_addr_2_addr)
	,.int_desc_11_data_host_addr_3_addr(int_desc_11_data_host_addr_3_addr)
	,.int_desc_11_wstrb_host_addr_0_addr(int_desc_11_wstrb_host_addr_0_addr)
	,.int_desc_11_wstrb_host_addr_1_addr(int_desc_11_wstrb_host_addr_1_addr)
	,.int_desc_11_wstrb_host_addr_2_addr(int_desc_11_wstrb_host_addr_2_addr)
	,.int_desc_11_wstrb_host_addr_3_addr(int_desc_11_wstrb_host_addr_3_addr)
	,.int_desc_12_data_host_addr_0_addr(int_desc_12_data_host_addr_0_addr)
	,.int_desc_12_data_host_addr_1_addr(int_desc_12_data_host_addr_1_addr)
	,.int_desc_12_data_host_addr_2_addr(int_desc_12_data_host_addr_2_addr)
	,.int_desc_12_data_host_addr_3_addr(int_desc_12_data_host_addr_3_addr)
	,.int_desc_12_wstrb_host_addr_0_addr(int_desc_12_wstrb_host_addr_0_addr)
	,.int_desc_12_wstrb_host_addr_1_addr(int_desc_12_wstrb_host_addr_1_addr)
	,.int_desc_12_wstrb_host_addr_2_addr(int_desc_12_wstrb_host_addr_2_addr)
	,.int_desc_12_wstrb_host_addr_3_addr(int_desc_12_wstrb_host_addr_3_addr)
	,.int_desc_13_data_host_addr_0_addr(int_desc_13_data_host_addr_0_addr)
	,.int_desc_13_data_host_addr_1_addr(int_desc_13_data_host_addr_1_addr)
	,.int_desc_13_data_host_addr_2_addr(int_desc_13_data_host_addr_2_addr)
	,.int_desc_13_data_host_addr_3_addr(int_desc_13_data_host_addr_3_addr)
	,.int_desc_13_wstrb_host_addr_0_addr(int_desc_13_wstrb_host_addr_0_addr)
	,.int_desc_13_wstrb_host_addr_1_addr(int_desc_13_wstrb_host_addr_1_addr)
	,.int_desc_13_wstrb_host_addr_2_addr(int_desc_13_wstrb_host_addr_2_addr)
	,.int_desc_13_wstrb_host_addr_3_addr(int_desc_13_wstrb_host_addr_3_addr)
	,.int_desc_14_data_host_addr_0_addr(int_desc_14_data_host_addr_0_addr)
	,.int_desc_14_data_host_addr_1_addr(int_desc_14_data_host_addr_1_addr)
	,.int_desc_14_data_host_addr_2_addr(int_desc_14_data_host_addr_2_addr)
	,.int_desc_14_data_host_addr_3_addr(int_desc_14_data_host_addr_3_addr)
	,.int_desc_14_wstrb_host_addr_0_addr(int_desc_14_wstrb_host_addr_0_addr)
	,.int_desc_14_wstrb_host_addr_1_addr(int_desc_14_wstrb_host_addr_1_addr)
	,.int_desc_14_wstrb_host_addr_2_addr(int_desc_14_wstrb_host_addr_2_addr)
	,.int_desc_14_wstrb_host_addr_3_addr(int_desc_14_wstrb_host_addr_3_addr)
	,.int_desc_15_data_host_addr_0_addr(int_desc_15_data_host_addr_0_addr)
	,.int_desc_15_data_host_addr_1_addr(int_desc_15_data_host_addr_1_addr)
	,.int_desc_15_data_host_addr_2_addr(int_desc_15_data_host_addr_2_addr)
	,.int_desc_15_data_host_addr_3_addr(int_desc_15_data_host_addr_3_addr)
	,.int_desc_15_wstrb_host_addr_0_addr(int_desc_15_wstrb_host_addr_0_addr)
	,.int_desc_15_wstrb_host_addr_1_addr(int_desc_15_wstrb_host_addr_1_addr)
	,.int_desc_15_wstrb_host_addr_2_addr(int_desc_15_wstrb_host_addr_2_addr)
	,.int_desc_15_wstrb_host_addr_3_addr(int_desc_15_wstrb_host_addr_3_addr)
	,.int_desc_0_xuser_0_xuser(int_desc_0_xuser_0_xuser)
	,.int_desc_0_xuser_1_xuser(int_desc_0_xuser_1_xuser)
	,.int_desc_0_xuser_2_xuser(int_desc_0_xuser_2_xuser)
	,.int_desc_0_xuser_3_xuser(int_desc_0_xuser_3_xuser)
	,.int_desc_0_xuser_4_xuser(int_desc_0_xuser_4_xuser)
	,.int_desc_0_xuser_5_xuser(int_desc_0_xuser_5_xuser)
	,.int_desc_0_xuser_6_xuser(int_desc_0_xuser_6_xuser)
	,.int_desc_0_xuser_7_xuser(int_desc_0_xuser_7_xuser)
	,.int_desc_0_xuser_8_xuser(int_desc_0_xuser_8_xuser)
	,.int_desc_0_xuser_9_xuser(int_desc_0_xuser_9_xuser)
	,.int_desc_0_xuser_10_xuser(int_desc_0_xuser_10_xuser)
	,.int_desc_0_xuser_11_xuser(int_desc_0_xuser_11_xuser)
	,.int_desc_0_xuser_12_xuser(int_desc_0_xuser_12_xuser)
	,.int_desc_0_xuser_13_xuser(int_desc_0_xuser_13_xuser)
	,.int_desc_0_xuser_14_xuser(int_desc_0_xuser_14_xuser)
	,.int_desc_0_xuser_15_xuser(int_desc_0_xuser_15_xuser)
	,.int_desc_1_xuser_0_xuser(int_desc_1_xuser_0_xuser)
	,.int_desc_1_xuser_1_xuser(int_desc_1_xuser_1_xuser)
	,.int_desc_1_xuser_2_xuser(int_desc_1_xuser_2_xuser)
	,.int_desc_1_xuser_3_xuser(int_desc_1_xuser_3_xuser)
	,.int_desc_1_xuser_4_xuser(int_desc_1_xuser_4_xuser)
	,.int_desc_1_xuser_5_xuser(int_desc_1_xuser_5_xuser)
	,.int_desc_1_xuser_6_xuser(int_desc_1_xuser_6_xuser)
	,.int_desc_1_xuser_7_xuser(int_desc_1_xuser_7_xuser)
	,.int_desc_1_xuser_8_xuser(int_desc_1_xuser_8_xuser)
	,.int_desc_1_xuser_9_xuser(int_desc_1_xuser_9_xuser)
	,.int_desc_1_xuser_10_xuser(int_desc_1_xuser_10_xuser)
	,.int_desc_1_xuser_11_xuser(int_desc_1_xuser_11_xuser)
	,.int_desc_1_xuser_12_xuser(int_desc_1_xuser_12_xuser)
	,.int_desc_1_xuser_13_xuser(int_desc_1_xuser_13_xuser)
	,.int_desc_1_xuser_14_xuser(int_desc_1_xuser_14_xuser)
	,.int_desc_1_xuser_15_xuser(int_desc_1_xuser_15_xuser)
	,.int_desc_2_xuser_0_xuser(int_desc_2_xuser_0_xuser)
	,.int_desc_2_xuser_1_xuser(int_desc_2_xuser_1_xuser)
	,.int_desc_2_xuser_2_xuser(int_desc_2_xuser_2_xuser)
	,.int_desc_2_xuser_3_xuser(int_desc_2_xuser_3_xuser)
	,.int_desc_2_xuser_4_xuser(int_desc_2_xuser_4_xuser)
	,.int_desc_2_xuser_5_xuser(int_desc_2_xuser_5_xuser)
	,.int_desc_2_xuser_6_xuser(int_desc_2_xuser_6_xuser)
	,.int_desc_2_xuser_7_xuser(int_desc_2_xuser_7_xuser)
	,.int_desc_2_xuser_8_xuser(int_desc_2_xuser_8_xuser)
	,.int_desc_2_xuser_9_xuser(int_desc_2_xuser_9_xuser)
	,.int_desc_2_xuser_10_xuser(int_desc_2_xuser_10_xuser)
	,.int_desc_2_xuser_11_xuser(int_desc_2_xuser_11_xuser)
	,.int_desc_2_xuser_12_xuser(int_desc_2_xuser_12_xuser)
	,.int_desc_2_xuser_13_xuser(int_desc_2_xuser_13_xuser)
	,.int_desc_2_xuser_14_xuser(int_desc_2_xuser_14_xuser)
	,.int_desc_2_xuser_15_xuser(int_desc_2_xuser_15_xuser)
	,.int_desc_3_xuser_0_xuser(int_desc_3_xuser_0_xuser)
	,.int_desc_3_xuser_1_xuser(int_desc_3_xuser_1_xuser)
	,.int_desc_3_xuser_2_xuser(int_desc_3_xuser_2_xuser)
	,.int_desc_3_xuser_3_xuser(int_desc_3_xuser_3_xuser)
	,.int_desc_3_xuser_4_xuser(int_desc_3_xuser_4_xuser)
	,.int_desc_3_xuser_5_xuser(int_desc_3_xuser_5_xuser)
	,.int_desc_3_xuser_6_xuser(int_desc_3_xuser_6_xuser)
	,.int_desc_3_xuser_7_xuser(int_desc_3_xuser_7_xuser)
	,.int_desc_3_xuser_8_xuser(int_desc_3_xuser_8_xuser)
	,.int_desc_3_xuser_9_xuser(int_desc_3_xuser_9_xuser)
	,.int_desc_3_xuser_10_xuser(int_desc_3_xuser_10_xuser)
	,.int_desc_3_xuser_11_xuser(int_desc_3_xuser_11_xuser)
	,.int_desc_3_xuser_12_xuser(int_desc_3_xuser_12_xuser)
	,.int_desc_3_xuser_13_xuser(int_desc_3_xuser_13_xuser)
	,.int_desc_3_xuser_14_xuser(int_desc_3_xuser_14_xuser)
	,.int_desc_3_xuser_15_xuser(int_desc_3_xuser_15_xuser)
	,.int_desc_4_xuser_0_xuser(int_desc_4_xuser_0_xuser)
	,.int_desc_4_xuser_1_xuser(int_desc_4_xuser_1_xuser)
	,.int_desc_4_xuser_2_xuser(int_desc_4_xuser_2_xuser)
	,.int_desc_4_xuser_3_xuser(int_desc_4_xuser_3_xuser)
	,.int_desc_4_xuser_4_xuser(int_desc_4_xuser_4_xuser)
	,.int_desc_4_xuser_5_xuser(int_desc_4_xuser_5_xuser)
	,.int_desc_4_xuser_6_xuser(int_desc_4_xuser_6_xuser)
	,.int_desc_4_xuser_7_xuser(int_desc_4_xuser_7_xuser)
	,.int_desc_4_xuser_8_xuser(int_desc_4_xuser_8_xuser)
	,.int_desc_4_xuser_9_xuser(int_desc_4_xuser_9_xuser)
	,.int_desc_4_xuser_10_xuser(int_desc_4_xuser_10_xuser)
	,.int_desc_4_xuser_11_xuser(int_desc_4_xuser_11_xuser)
	,.int_desc_4_xuser_12_xuser(int_desc_4_xuser_12_xuser)
	,.int_desc_4_xuser_13_xuser(int_desc_4_xuser_13_xuser)
	,.int_desc_4_xuser_14_xuser(int_desc_4_xuser_14_xuser)
	,.int_desc_4_xuser_15_xuser(int_desc_4_xuser_15_xuser)
	,.int_desc_5_xuser_0_xuser(int_desc_5_xuser_0_xuser)
	,.int_desc_5_xuser_1_xuser(int_desc_5_xuser_1_xuser)
	,.int_desc_5_xuser_2_xuser(int_desc_5_xuser_2_xuser)
	,.int_desc_5_xuser_3_xuser(int_desc_5_xuser_3_xuser)
	,.int_desc_5_xuser_4_xuser(int_desc_5_xuser_4_xuser)
	,.int_desc_5_xuser_5_xuser(int_desc_5_xuser_5_xuser)
	,.int_desc_5_xuser_6_xuser(int_desc_5_xuser_6_xuser)
	,.int_desc_5_xuser_7_xuser(int_desc_5_xuser_7_xuser)
	,.int_desc_5_xuser_8_xuser(int_desc_5_xuser_8_xuser)
	,.int_desc_5_xuser_9_xuser(int_desc_5_xuser_9_xuser)
	,.int_desc_5_xuser_10_xuser(int_desc_5_xuser_10_xuser)
	,.int_desc_5_xuser_11_xuser(int_desc_5_xuser_11_xuser)
	,.int_desc_5_xuser_12_xuser(int_desc_5_xuser_12_xuser)
	,.int_desc_5_xuser_13_xuser(int_desc_5_xuser_13_xuser)
	,.int_desc_5_xuser_14_xuser(int_desc_5_xuser_14_xuser)
	,.int_desc_5_xuser_15_xuser(int_desc_5_xuser_15_xuser)
	,.int_desc_6_xuser_0_xuser(int_desc_6_xuser_0_xuser)
	,.int_desc_6_xuser_1_xuser(int_desc_6_xuser_1_xuser)
	,.int_desc_6_xuser_2_xuser(int_desc_6_xuser_2_xuser)
	,.int_desc_6_xuser_3_xuser(int_desc_6_xuser_3_xuser)
	,.int_desc_6_xuser_4_xuser(int_desc_6_xuser_4_xuser)
	,.int_desc_6_xuser_5_xuser(int_desc_6_xuser_5_xuser)
	,.int_desc_6_xuser_6_xuser(int_desc_6_xuser_6_xuser)
	,.int_desc_6_xuser_7_xuser(int_desc_6_xuser_7_xuser)
	,.int_desc_6_xuser_8_xuser(int_desc_6_xuser_8_xuser)
	,.int_desc_6_xuser_9_xuser(int_desc_6_xuser_9_xuser)
	,.int_desc_6_xuser_10_xuser(int_desc_6_xuser_10_xuser)
	,.int_desc_6_xuser_11_xuser(int_desc_6_xuser_11_xuser)
	,.int_desc_6_xuser_12_xuser(int_desc_6_xuser_12_xuser)
	,.int_desc_6_xuser_13_xuser(int_desc_6_xuser_13_xuser)
	,.int_desc_6_xuser_14_xuser(int_desc_6_xuser_14_xuser)
	,.int_desc_6_xuser_15_xuser(int_desc_6_xuser_15_xuser)
	,.int_desc_7_xuser_0_xuser(int_desc_7_xuser_0_xuser)
	,.int_desc_7_xuser_1_xuser(int_desc_7_xuser_1_xuser)
	,.int_desc_7_xuser_2_xuser(int_desc_7_xuser_2_xuser)
	,.int_desc_7_xuser_3_xuser(int_desc_7_xuser_3_xuser)
	,.int_desc_7_xuser_4_xuser(int_desc_7_xuser_4_xuser)
	,.int_desc_7_xuser_5_xuser(int_desc_7_xuser_5_xuser)
	,.int_desc_7_xuser_6_xuser(int_desc_7_xuser_6_xuser)
	,.int_desc_7_xuser_7_xuser(int_desc_7_xuser_7_xuser)
	,.int_desc_7_xuser_8_xuser(int_desc_7_xuser_8_xuser)
	,.int_desc_7_xuser_9_xuser(int_desc_7_xuser_9_xuser)
	,.int_desc_7_xuser_10_xuser(int_desc_7_xuser_10_xuser)
	,.int_desc_7_xuser_11_xuser(int_desc_7_xuser_11_xuser)
	,.int_desc_7_xuser_12_xuser(int_desc_7_xuser_12_xuser)
	,.int_desc_7_xuser_13_xuser(int_desc_7_xuser_13_xuser)
	,.int_desc_7_xuser_14_xuser(int_desc_7_xuser_14_xuser)
	,.int_desc_7_xuser_15_xuser(int_desc_7_xuser_15_xuser)
	,.int_desc_8_xuser_0_xuser(int_desc_8_xuser_0_xuser)
	,.int_desc_8_xuser_1_xuser(int_desc_8_xuser_1_xuser)
	,.int_desc_8_xuser_2_xuser(int_desc_8_xuser_2_xuser)
	,.int_desc_8_xuser_3_xuser(int_desc_8_xuser_3_xuser)
	,.int_desc_8_xuser_4_xuser(int_desc_8_xuser_4_xuser)
	,.int_desc_8_xuser_5_xuser(int_desc_8_xuser_5_xuser)
	,.int_desc_8_xuser_6_xuser(int_desc_8_xuser_6_xuser)
	,.int_desc_8_xuser_7_xuser(int_desc_8_xuser_7_xuser)
	,.int_desc_8_xuser_8_xuser(int_desc_8_xuser_8_xuser)
	,.int_desc_8_xuser_9_xuser(int_desc_8_xuser_9_xuser)
	,.int_desc_8_xuser_10_xuser(int_desc_8_xuser_10_xuser)
	,.int_desc_8_xuser_11_xuser(int_desc_8_xuser_11_xuser)
	,.int_desc_8_xuser_12_xuser(int_desc_8_xuser_12_xuser)
	,.int_desc_8_xuser_13_xuser(int_desc_8_xuser_13_xuser)
	,.int_desc_8_xuser_14_xuser(int_desc_8_xuser_14_xuser)
	,.int_desc_8_xuser_15_xuser(int_desc_8_xuser_15_xuser)
	,.int_desc_9_xuser_0_xuser(int_desc_9_xuser_0_xuser)
	,.int_desc_9_xuser_1_xuser(int_desc_9_xuser_1_xuser)
	,.int_desc_9_xuser_2_xuser(int_desc_9_xuser_2_xuser)
	,.int_desc_9_xuser_3_xuser(int_desc_9_xuser_3_xuser)
	,.int_desc_9_xuser_4_xuser(int_desc_9_xuser_4_xuser)
	,.int_desc_9_xuser_5_xuser(int_desc_9_xuser_5_xuser)
	,.int_desc_9_xuser_6_xuser(int_desc_9_xuser_6_xuser)
	,.int_desc_9_xuser_7_xuser(int_desc_9_xuser_7_xuser)
	,.int_desc_9_xuser_8_xuser(int_desc_9_xuser_8_xuser)
	,.int_desc_9_xuser_9_xuser(int_desc_9_xuser_9_xuser)
	,.int_desc_9_xuser_10_xuser(int_desc_9_xuser_10_xuser)
	,.int_desc_9_xuser_11_xuser(int_desc_9_xuser_11_xuser)
	,.int_desc_9_xuser_12_xuser(int_desc_9_xuser_12_xuser)
	,.int_desc_9_xuser_13_xuser(int_desc_9_xuser_13_xuser)
	,.int_desc_9_xuser_14_xuser(int_desc_9_xuser_14_xuser)
	,.int_desc_9_xuser_15_xuser(int_desc_9_xuser_15_xuser)
	,.int_desc_10_xuser_0_xuser(int_desc_10_xuser_0_xuser)
	,.int_desc_10_xuser_1_xuser(int_desc_10_xuser_1_xuser)
	,.int_desc_10_xuser_2_xuser(int_desc_10_xuser_2_xuser)
	,.int_desc_10_xuser_3_xuser(int_desc_10_xuser_3_xuser)
	,.int_desc_10_xuser_4_xuser(int_desc_10_xuser_4_xuser)
	,.int_desc_10_xuser_5_xuser(int_desc_10_xuser_5_xuser)
	,.int_desc_10_xuser_6_xuser(int_desc_10_xuser_6_xuser)
	,.int_desc_10_xuser_7_xuser(int_desc_10_xuser_7_xuser)
	,.int_desc_10_xuser_8_xuser(int_desc_10_xuser_8_xuser)
	,.int_desc_10_xuser_9_xuser(int_desc_10_xuser_9_xuser)
	,.int_desc_10_xuser_10_xuser(int_desc_10_xuser_10_xuser)
	,.int_desc_10_xuser_11_xuser(int_desc_10_xuser_11_xuser)
	,.int_desc_10_xuser_12_xuser(int_desc_10_xuser_12_xuser)
	,.int_desc_10_xuser_13_xuser(int_desc_10_xuser_13_xuser)
	,.int_desc_10_xuser_14_xuser(int_desc_10_xuser_14_xuser)
	,.int_desc_10_xuser_15_xuser(int_desc_10_xuser_15_xuser)
	,.int_desc_11_xuser_0_xuser(int_desc_11_xuser_0_xuser)
	,.int_desc_11_xuser_1_xuser(int_desc_11_xuser_1_xuser)
	,.int_desc_11_xuser_2_xuser(int_desc_11_xuser_2_xuser)
	,.int_desc_11_xuser_3_xuser(int_desc_11_xuser_3_xuser)
	,.int_desc_11_xuser_4_xuser(int_desc_11_xuser_4_xuser)
	,.int_desc_11_xuser_5_xuser(int_desc_11_xuser_5_xuser)
	,.int_desc_11_xuser_6_xuser(int_desc_11_xuser_6_xuser)
	,.int_desc_11_xuser_7_xuser(int_desc_11_xuser_7_xuser)
	,.int_desc_11_xuser_8_xuser(int_desc_11_xuser_8_xuser)
	,.int_desc_11_xuser_9_xuser(int_desc_11_xuser_9_xuser)
	,.int_desc_11_xuser_10_xuser(int_desc_11_xuser_10_xuser)
	,.int_desc_11_xuser_11_xuser(int_desc_11_xuser_11_xuser)
	,.int_desc_11_xuser_12_xuser(int_desc_11_xuser_12_xuser)
	,.int_desc_11_xuser_13_xuser(int_desc_11_xuser_13_xuser)
	,.int_desc_11_xuser_14_xuser(int_desc_11_xuser_14_xuser)
	,.int_desc_11_xuser_15_xuser(int_desc_11_xuser_15_xuser)
	,.int_desc_12_xuser_0_xuser(int_desc_12_xuser_0_xuser)
	,.int_desc_12_xuser_1_xuser(int_desc_12_xuser_1_xuser)
	,.int_desc_12_xuser_2_xuser(int_desc_12_xuser_2_xuser)
	,.int_desc_12_xuser_3_xuser(int_desc_12_xuser_3_xuser)
	,.int_desc_12_xuser_4_xuser(int_desc_12_xuser_4_xuser)
	,.int_desc_12_xuser_5_xuser(int_desc_12_xuser_5_xuser)
	,.int_desc_12_xuser_6_xuser(int_desc_12_xuser_6_xuser)
	,.int_desc_12_xuser_7_xuser(int_desc_12_xuser_7_xuser)
	,.int_desc_12_xuser_8_xuser(int_desc_12_xuser_8_xuser)
	,.int_desc_12_xuser_9_xuser(int_desc_12_xuser_9_xuser)
	,.int_desc_12_xuser_10_xuser(int_desc_12_xuser_10_xuser)
	,.int_desc_12_xuser_11_xuser(int_desc_12_xuser_11_xuser)
	,.int_desc_12_xuser_12_xuser(int_desc_12_xuser_12_xuser)
	,.int_desc_12_xuser_13_xuser(int_desc_12_xuser_13_xuser)
	,.int_desc_12_xuser_14_xuser(int_desc_12_xuser_14_xuser)
	,.int_desc_12_xuser_15_xuser(int_desc_12_xuser_15_xuser)
	,.int_desc_13_xuser_0_xuser(int_desc_13_xuser_0_xuser)
	,.int_desc_13_xuser_1_xuser(int_desc_13_xuser_1_xuser)
	,.int_desc_13_xuser_2_xuser(int_desc_13_xuser_2_xuser)
	,.int_desc_13_xuser_3_xuser(int_desc_13_xuser_3_xuser)
	,.int_desc_13_xuser_4_xuser(int_desc_13_xuser_4_xuser)
	,.int_desc_13_xuser_5_xuser(int_desc_13_xuser_5_xuser)
	,.int_desc_13_xuser_6_xuser(int_desc_13_xuser_6_xuser)
	,.int_desc_13_xuser_7_xuser(int_desc_13_xuser_7_xuser)
	,.int_desc_13_xuser_8_xuser(int_desc_13_xuser_8_xuser)
	,.int_desc_13_xuser_9_xuser(int_desc_13_xuser_9_xuser)
	,.int_desc_13_xuser_10_xuser(int_desc_13_xuser_10_xuser)
	,.int_desc_13_xuser_11_xuser(int_desc_13_xuser_11_xuser)
	,.int_desc_13_xuser_12_xuser(int_desc_13_xuser_12_xuser)
	,.int_desc_13_xuser_13_xuser(int_desc_13_xuser_13_xuser)
	,.int_desc_13_xuser_14_xuser(int_desc_13_xuser_14_xuser)
	,.int_desc_13_xuser_15_xuser(int_desc_13_xuser_15_xuser)
	,.int_desc_14_xuser_0_xuser(int_desc_14_xuser_0_xuser)
	,.int_desc_14_xuser_1_xuser(int_desc_14_xuser_1_xuser)
	,.int_desc_14_xuser_2_xuser(int_desc_14_xuser_2_xuser)
	,.int_desc_14_xuser_3_xuser(int_desc_14_xuser_3_xuser)
	,.int_desc_14_xuser_4_xuser(int_desc_14_xuser_4_xuser)
	,.int_desc_14_xuser_5_xuser(int_desc_14_xuser_5_xuser)
	,.int_desc_14_xuser_6_xuser(int_desc_14_xuser_6_xuser)
	,.int_desc_14_xuser_7_xuser(int_desc_14_xuser_7_xuser)
	,.int_desc_14_xuser_8_xuser(int_desc_14_xuser_8_xuser)
	,.int_desc_14_xuser_9_xuser(int_desc_14_xuser_9_xuser)
	,.int_desc_14_xuser_10_xuser(int_desc_14_xuser_10_xuser)
	,.int_desc_14_xuser_11_xuser(int_desc_14_xuser_11_xuser)
	,.int_desc_14_xuser_12_xuser(int_desc_14_xuser_12_xuser)
	,.int_desc_14_xuser_13_xuser(int_desc_14_xuser_13_xuser)
	,.int_desc_14_xuser_14_xuser(int_desc_14_xuser_14_xuser)
	,.int_desc_14_xuser_15_xuser(int_desc_14_xuser_15_xuser)
	,.int_desc_15_xuser_0_xuser(int_desc_15_xuser_0_xuser)
	,.int_desc_15_xuser_1_xuser(int_desc_15_xuser_1_xuser)
	,.int_desc_15_xuser_2_xuser(int_desc_15_xuser_2_xuser)
	,.int_desc_15_xuser_3_xuser(int_desc_15_xuser_3_xuser)
	,.int_desc_15_xuser_4_xuser(int_desc_15_xuser_4_xuser)
	,.int_desc_15_xuser_5_xuser(int_desc_15_xuser_5_xuser)
	,.int_desc_15_xuser_6_xuser(int_desc_15_xuser_6_xuser)
	,.int_desc_15_xuser_7_xuser(int_desc_15_xuser_7_xuser)
	,.int_desc_15_xuser_8_xuser(int_desc_15_xuser_8_xuser)
	,.int_desc_15_xuser_9_xuser(int_desc_15_xuser_9_xuser)
	,.int_desc_15_xuser_10_xuser(int_desc_15_xuser_10_xuser)
	,.int_desc_15_xuser_11_xuser(int_desc_15_xuser_11_xuser)
	,.int_desc_15_xuser_12_xuser(int_desc_15_xuser_12_xuser)
	,.int_desc_15_xuser_13_xuser(int_desc_15_xuser_13_xuser)
	,.int_desc_15_xuser_14_xuser(int_desc_15_xuser_14_xuser)
	,.int_desc_15_xuser_15_xuser(int_desc_15_xuser_15_xuser)
        ,.rb2uc_rd_data(rb2uc_rd_data)
        ,.hm2uc_done(hm2uc_done)

);

//////////////////////
//Tie all uc2rb_<reg>_reg_we to high because current implementation of uc2rb_<reg>_reg 
//such that it will always hold intended correct value.
//////////////////////
assign uc2rb_intr_error_status_reg_we = 32'hFFFFFFFF;
assign uc2rb_ownership_reg_we = 32'hFFFFFFFF;
assign uc2rb_intr_txn_avail_status_reg_we = 32'hFFFFFFFF;
assign uc2rb_intr_comp_status_reg_we = 32'hFFFFFFFF;
assign uc2rb_status_busy_reg_we = 32'hFFFFFFFF;
assign uc2rb_resp_fifo_free_level_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_0_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_1_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_2_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_3_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_4_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_5_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_6_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_7_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_8_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_9_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_10_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_11_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_12_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_13_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_14_wuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_txn_type_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_size_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_data_offset_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axsize_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_attr_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axaddr_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axaddr_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axaddr_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axaddr_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axid_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axid_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axid_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axid_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_axuser_15_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_0_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_1_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_2_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_3_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_4_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_5_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_6_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_7_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_8_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_9_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_10_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_11_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_12_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_13_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_14_reg_we = 32'hFFFFFFFF;
assign uc2rb_desc_15_wuser_15_reg_we = 32'hFFFFFFFF;

endmodule

